
module SNPS_CLOCK_GATE_HIGH_riscv_alu_div_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_alu_div_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_alu_div_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_30 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_29 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_28 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_27 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_26 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_25 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_24 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_23 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_22 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_21 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_20 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_19 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_18 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_17 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_16 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_15 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_14 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_13 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_12 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_11 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_10 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_9 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_8 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_7 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_6 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_5 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_4 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_3 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_2 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_1 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_0 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_L0_buffer_RDATA_IN_WIDTH128_2 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_L0_buffer_RDATA_IN_WIDTH128_1 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_L0_buffer_RDATA_IN_WIDTH128_0 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module riscv_alu_div ( Clk_CI, Rst_RBI, OpA_DI, OpB_DI, OpBShift_DI, 
        OpBIsZero_SI, OpBSign_SI, OpCode_SI, InVld_SI, OutRdy_SI, OutVld_SO, 
        Res_DO );
  input [31:0] OpA_DI;
  input [31:0] OpB_DI;
  input [5:0] OpBShift_DI;
  input [1:0] OpCode_SI;
  output [31:0] Res_DO;
  input Clk_CI, Rst_RBI, OpBIsZero_SI, OpBSign_SI, InVld_SI, OutRdy_SI;
  output OutVld_SO;
  wire   CompInv_SP, RemSel_SP, ResInv_SP, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n277, n278, n279, n280, n281, n282, n283, n284, n1,
         n2, n3, n5, n6, n7, n12, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n208, n213, n231, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n566, n570, n571, n574, n575,
         n576, n577, n578, n579, n580, n582, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n815, n817, n820, n821, n823, n824, n825,
         n826, n827, n828, n829, n830, n835, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1092, n1093, n1094, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159;
  wire   [31:0] BReg_DP;
  wire   [31:0] ResReg_DP_rev;
  wire   [31:0] AReg_DP;
  wire   [5:0] Cnt_DP;
  wire   [1:0] State_SP;

  INV_X1 U10 ( .A(n3), .ZN(n6) );
  NAND2_X1 U16 ( .A1(n594), .A2(AReg_DP[0]), .ZN(n21) );
  NAND2_X2 U17 ( .A1(n579), .A2(n830), .ZN(n577) );
  AOI21_X1 U21 ( .B1(n412), .B2(n410), .A(n369), .ZN(n407) );
  XNOR2_X1 U23 ( .A(n376), .B(n375), .ZN(n14) );
  XNOR2_X1 U24 ( .A(n613), .B(n603), .ZN(n602) );
  XNOR2_X1 U25 ( .A(n621), .B(n618), .ZN(n619) );
  AND2_X1 U27 ( .A1(n637), .A2(n636), .ZN(n641) );
  XNOR2_X1 U28 ( .A(n637), .B(n634), .ZN(n635) );
  XNOR2_X1 U29 ( .A(n661), .B(n658), .ZN(n659) );
  AND2_X1 U31 ( .A1(n653), .A2(n652), .ZN(n657) );
  AND2_X1 U32 ( .A1(n621), .A2(n620), .ZN(n625) );
  XNOR2_X1 U33 ( .A(n653), .B(n650), .ZN(n651) );
  AND2_X1 U34 ( .A1(n717), .A2(n716), .ZN(n721) );
  AND2_X1 U35 ( .A1(n709), .A2(n708), .ZN(n713) );
  XNOR2_X1 U36 ( .A(n709), .B(n706), .ZN(n707) );
  XNOR2_X1 U37 ( .A(n717), .B(n714), .ZN(n715) );
  NOR2_X1 U38 ( .A1(State_SP[1]), .A2(State_SP[0]), .ZN(n16) );
  OAI21_X1 U39 ( .B1(n407), .B2(n373), .A(n372), .ZN(n399) );
  INV_X1 U40 ( .A(n1086), .ZN(n570) );
  XOR2_X1 U41 ( .A(OpA_DI[31]), .B(OpBSign_SI), .Z(n15) );
  NAND2_X1 U42 ( .A1(n15), .A2(OpCode_SI[0]), .ZN(n588) );
  NAND2_X1 U44 ( .A1(n588), .A2(n586), .ZN(n19) );
  MUX2_X1 U45 ( .A(BReg_DP[1]), .B(OpA_DI[1]), .S(n586), .Z(n17) );
  XOR2_X1 U46 ( .A(n12), .B(n17), .Z(n24) );
  NOR2_X1 U47 ( .A1(n586), .A2(n754), .ZN(n23) );
  NOR2_X1 U48 ( .A1(n24), .A2(n23), .ZN(n529) );
  MUX2_X1 U49 ( .A(BReg_DP[2]), .B(OpA_DI[2]), .S(n586), .Z(n18) );
  XOR2_X1 U50 ( .A(n12), .B(n18), .Z(n26) );
  INV_X1 U51 ( .A(n586), .ZN(n594) );
  AND2_X1 U52 ( .A1(n594), .A2(AReg_DP[2]), .ZN(n25) );
  NOR2_X1 U54 ( .A1(n529), .A2(n523), .ZN(n28) );
  MUX2_X1 U55 ( .A(BReg_DP[0]), .B(OpA_DI[0]), .S(n586), .Z(n20) );
  XOR2_X1 U56 ( .A(n12), .B(n20), .Z(n536) );
  INV_X1 U57 ( .A(n536), .ZN(n22) );
  INV_X1 U58 ( .A(n12), .ZN(n535) );
  OAI21_X1 U59 ( .B1(n22), .B2(n535), .A(n21), .ZN(n522) );
  NAND2_X1 U60 ( .A1(n24), .A2(n23), .ZN(n530) );
  NAND2_X1 U61 ( .A1(n26), .A2(n25), .ZN(n524) );
  OAI21_X1 U62 ( .B1(n523), .B2(n530), .A(n524), .ZN(n27) );
  AOI21_X1 U63 ( .B1(n28), .B2(n522), .A(n27), .ZN(n494) );
  MUX2_X1 U64 ( .A(BReg_DP[3]), .B(OpA_DI[3]), .S(n586), .Z(n29) );
  XOR2_X1 U65 ( .A(n12), .B(n29), .Z(n34) );
  AND2_X1 U66 ( .A1(n829), .A2(AReg_DP[3]), .ZN(n33) );
  NOR2_X1 U67 ( .A1(n34), .A2(n33), .ZN(n509) );
  MUX2_X1 U68 ( .A(BReg_DP[4]), .B(OpA_DI[4]), .S(n586), .Z(n30) );
  XOR2_X1 U69 ( .A(n12), .B(n30), .Z(n36) );
  AND2_X1 U70 ( .A1(n830), .A2(AReg_DP[4]), .ZN(n35) );
  NOR2_X1 U71 ( .A1(n36), .A2(n35), .ZN(n511) );
  NOR2_X1 U72 ( .A1(n509), .A2(n511), .ZN(n496) );
  MUX2_X1 U73 ( .A(BReg_DP[5]), .B(OpA_DI[5]), .S(n586), .Z(n31) );
  XOR2_X1 U74 ( .A(n12), .B(n31), .Z(n38) );
  AND2_X1 U75 ( .A1(n830), .A2(AReg_DP[5]), .ZN(n37) );
  NOR2_X1 U76 ( .A1(n38), .A2(n37), .ZN(n503) );
  MUX2_X1 U77 ( .A(BReg_DP[6]), .B(OpA_DI[6]), .S(n586), .Z(n32) );
  XOR2_X1 U78 ( .A(n12), .B(n32), .Z(n40) );
  AND2_X1 U79 ( .A1(n830), .A2(AReg_DP[6]), .ZN(n39) );
  NOR2_X1 U80 ( .A1(n40), .A2(n39), .ZN(n497) );
  NOR2_X1 U81 ( .A1(n503), .A2(n497), .ZN(n42) );
  NAND2_X1 U82 ( .A1(n496), .A2(n42), .ZN(n44) );
  NAND2_X1 U83 ( .A1(n34), .A2(n33), .ZN(n517) );
  NAND2_X1 U84 ( .A1(n36), .A2(n35), .ZN(n512) );
  OAI21_X1 U85 ( .B1(n511), .B2(n517), .A(n512), .ZN(n495) );
  NAND2_X1 U86 ( .A1(n38), .A2(n37), .ZN(n504) );
  NAND2_X1 U87 ( .A1(n40), .A2(n39), .ZN(n498) );
  OAI21_X1 U88 ( .B1(n497), .B2(n504), .A(n498), .ZN(n41) );
  AOI21_X1 U89 ( .B1(n42), .B2(n495), .A(n41), .ZN(n43) );
  OAI21_X1 U90 ( .B1(n494), .B2(n44), .A(n43), .ZN(n481) );
  MUX2_X1 U91 ( .A(BReg_DP[7]), .B(OpA_DI[7]), .S(n586), .Z(n45) );
  XOR2_X1 U92 ( .A(n12), .B(n45), .Z(n48) );
  NOR2_X1 U93 ( .A1(n566), .A2(n732), .ZN(n47) );
  NOR2_X1 U94 ( .A1(n48), .A2(n47), .ZN(n488) );
  MUX2_X1 U95 ( .A(BReg_DP[8]), .B(OpA_DI[8]), .S(n586), .Z(n46) );
  XOR2_X1 U96 ( .A(n12), .B(n46), .Z(n50) );
  AND2_X1 U97 ( .A1(n830), .A2(AReg_DP[8]), .ZN(n49) );
  NOR2_X1 U98 ( .A1(n50), .A2(n49), .ZN(n482) );
  NOR2_X1 U99 ( .A1(n488), .A2(n482), .ZN(n52) );
  NAND2_X1 U100 ( .A1(n48), .A2(n47), .ZN(n489) );
  NAND2_X1 U101 ( .A1(n50), .A2(n49), .ZN(n483) );
  OAI21_X1 U102 ( .B1(n482), .B2(n489), .A(n483), .ZN(n51) );
  AOI21_X1 U103 ( .B1(n481), .B2(n52), .A(n51), .ZN(n479) );
  MUX2_X1 U104 ( .A(BReg_DP[9]), .B(OpA_DI[9]), .S(n586), .Z(n53) );
  XOR2_X1 U105 ( .A(n12), .B(n53), .Z(n55) );
  AND2_X1 U106 ( .A1(n829), .A2(AReg_DP[9]), .ZN(n54) );
  NOR2_X1 U107 ( .A1(n55), .A2(n54), .ZN(n475) );
  NAND2_X1 U108 ( .A1(n55), .A2(n54), .ZN(n476) );
  OAI21_X1 U109 ( .B1(n479), .B2(n475), .A(n476), .ZN(n473) );
  MUX2_X1 U110 ( .A(BReg_DP[10]), .B(OpA_DI[10]), .S(n586), .Z(n56) );
  XOR2_X1 U111 ( .A(n12), .B(n56), .Z(n58) );
  AND2_X1 U112 ( .A1(n594), .A2(AReg_DP[10]), .ZN(n57) );
  OR2_X1 U113 ( .A1(n58), .A2(n57), .ZN(n471) );
  NAND2_X1 U114 ( .A1(n58), .A2(n57), .ZN(n470) );
  INV_X1 U115 ( .A(n470), .ZN(n59) );
  AOI21_X1 U116 ( .B1(n473), .B2(n471), .A(n59), .ZN(n468) );
  MUX2_X1 U117 ( .A(BReg_DP[11]), .B(OpA_DI[11]), .S(n586), .Z(n60) );
  XOR2_X1 U118 ( .A(n12), .B(n60), .Z(n62) );
  AND2_X1 U119 ( .A1(n594), .A2(AReg_DP[11]), .ZN(n61) );
  NOR2_X1 U120 ( .A1(n62), .A2(n61), .ZN(n464) );
  NAND2_X1 U121 ( .A1(n62), .A2(n61), .ZN(n465) );
  OAI21_X1 U122 ( .B1(n468), .B2(n464), .A(n465), .ZN(n334) );
  MUX2_X1 U123 ( .A(BReg_DP[12]), .B(OpA_DI[12]), .S(n586), .Z(n63) );
  XOR2_X1 U124 ( .A(n12), .B(n63), .Z(n65) );
  AND2_X1 U125 ( .A1(n829), .A2(AReg_DP[12]), .ZN(n64) );
  OR2_X1 U126 ( .A1(n65), .A2(n64), .ZN(n333) );
  NAND2_X1 U127 ( .A1(n65), .A2(n64), .ZN(n331) );
  NAND2_X1 U128 ( .A1(n333), .A2(n331), .ZN(n66) );
  XNOR2_X1 U129 ( .A(n334), .B(n66), .ZN(n205) );
  NOR4_X1 U130 ( .A1(AReg_DP[31]), .A2(AReg_DP[2]), .A3(AReg_DP[30]), .A4(
        AReg_DP[1]), .ZN(n70) );
  NOR4_X1 U131 ( .A1(AReg_DP[3]), .A2(AReg_DP[4]), .A3(AReg_DP[5]), .A4(
        AReg_DP[6]), .ZN(n69) );
  NOR4_X1 U132 ( .A1(AReg_DP[8]), .A2(AReg_DP[9]), .A3(AReg_DP[10]), .A4(
        AReg_DP[11]), .ZN(n68) );
  NOR4_X1 U133 ( .A1(AReg_DP[7]), .A2(AReg_DP[0]), .A3(AReg_DP[16]), .A4(
        AReg_DP[21]), .ZN(n67) );
  NAND4_X1 U134 ( .A1(n70), .A2(n69), .A3(n68), .A4(n67), .ZN(n76) );
  NOR4_X1 U135 ( .A1(AReg_DP[12]), .A2(AReg_DP[13]), .A3(AReg_DP[14]), .A4(
        AReg_DP[15]), .ZN(n74) );
  NOR4_X1 U136 ( .A1(AReg_DP[17]), .A2(AReg_DP[18]), .A3(AReg_DP[19]), .A4(
        AReg_DP[20]), .ZN(n73) );
  NOR4_X1 U137 ( .A1(AReg_DP[22]), .A2(AReg_DP[23]), .A3(AReg_DP[24]), .A4(
        AReg_DP[25]), .ZN(n72) );
  NOR4_X1 U138 ( .A1(AReg_DP[26]), .A2(AReg_DP[27]), .A3(AReg_DP[28]), .A4(
        AReg_DP[29]), .ZN(n71) );
  NAND4_X1 U139 ( .A1(n74), .A2(n73), .A3(n72), .A4(n71), .ZN(n75) );
  OR3_X1 U140 ( .A1(OpBIsZero_SI), .A2(n76), .A3(n75), .ZN(n204) );
  NOR2_X2 U141 ( .A1(n802), .A2(State_SP[1]), .ZN(n580) );
  NOR2_X1 U142 ( .A1(n790), .A2(AReg_DP[31]), .ZN(n78) );
  AOI21_X1 U143 ( .B1(BReg_DP[30]), .B2(n772), .A(n78), .ZN(n174) );
  NOR2_X1 U144 ( .A1(n773), .A2(AReg_DP[29]), .ZN(n134) );
  NAND2_X1 U145 ( .A1(n809), .A2(AReg_DP[28]), .ZN(n154) );
  NAND2_X1 U146 ( .A1(n773), .A2(AReg_DP[29]), .ZN(n153) );
  OAI21_X1 U147 ( .B1(n134), .B2(n154), .A(n153), .ZN(n140) );
  NAND2_X1 U148 ( .A1(n810), .A2(AReg_DP[30]), .ZN(n151) );
  AND2_X1 U149 ( .A1(n790), .A2(AReg_DP[31]), .ZN(n170) );
  INV_X1 U150 ( .A(n170), .ZN(n77) );
  OAI21_X1 U151 ( .B1(n78), .B2(n151), .A(n77), .ZN(n139) );
  NOR2_X1 U152 ( .A1(n799), .A2(AReg_DP[20]), .ZN(n79) );
  NAND2_X1 U153 ( .A1(n804), .A2(BReg_DP[23]), .ZN(n122) );
  OAI21_X1 U154 ( .B1(AReg_DP[22]), .B2(n811), .A(n122), .ZN(n119) );
  AOI211_X1 U155 ( .C1(BReg_DP[21]), .C2(n748), .A(n79), .B(n119), .ZN(n191)
         );
  NOR2_X1 U156 ( .A1(n792), .A2(BReg_DP[11]), .ZN(n150) );
  NOR2_X1 U157 ( .A1(n751), .A2(AReg_DP[15]), .ZN(n104) );
  NOR2_X1 U158 ( .A1(n759), .A2(AReg_DP[12]), .ZN(n80) );
  NOR2_X1 U159 ( .A1(n104), .A2(n80), .ZN(n82) );
  NOR2_X1 U160 ( .A1(n753), .A2(AReg_DP[14]), .ZN(n103) );
  INV_X1 U161 ( .A(n103), .ZN(n81) );
  OR2_X1 U162 ( .A1(n755), .A2(AReg_DP[13]), .ZN(n102) );
  AND3_X1 U163 ( .A1(n82), .A2(n81), .A3(n102), .ZN(n194) );
  NOR2_X1 U164 ( .A1(n758), .A2(AReg_DP[11]), .ZN(n101) );
  AOI22_X1 U165 ( .A1(AReg_DP[8]), .A2(n761), .B1(n733), .B2(AReg_DP[9]), .ZN(
        n183) );
  NOR2_X1 U166 ( .A1(n733), .A2(AReg_DP[9]), .ZN(n95) );
  NOR2_X1 U167 ( .A1(n183), .A2(n95), .ZN(n83) );
  AND2_X1 U168 ( .A1(n769), .A2(AReg_DP[10]), .ZN(n168) );
  NAND2_X1 U169 ( .A1(n806), .A2(BReg_DP[10]), .ZN(n97) );
  OAI21_X1 U170 ( .B1(n83), .B2(n168), .A(n97), .ZN(n100) );
  NAND2_X1 U171 ( .A1(n750), .A2(AReg_DP[6]), .ZN(n162) );
  OAI21_X1 U172 ( .B1(n162), .B2(n732), .A(BReg_DP[7]), .ZN(n94) );
  NAND2_X1 U173 ( .A1(n162), .A2(n732), .ZN(n93) );
  NAND2_X1 U174 ( .A1(n762), .A2(BReg_DP[2]), .ZN(n187) );
  OAI21_X1 U175 ( .B1(AReg_DP[0]), .B2(n752), .A(n187), .ZN(n85) );
  AOI21_X1 U176 ( .B1(n752), .B2(AReg_DP[0]), .A(AReg_DP[1]), .ZN(n84) );
  NAND2_X1 U177 ( .A1(n766), .A2(AReg_DP[3]), .ZN(n186) );
  NAND2_X1 U178 ( .A1(n767), .A2(AReg_DP[2]), .ZN(n185) );
  OAI211_X1 U179 ( .C1(n85), .C2(n84), .A(n186), .B(n185), .ZN(n89) );
  NAND2_X1 U180 ( .A1(n763), .A2(BReg_DP[3]), .ZN(n180) );
  INV_X1 U181 ( .A(n180), .ZN(n86) );
  NOR2_X1 U182 ( .A1(n749), .A2(AReg_DP[4]), .ZN(n149) );
  NOR2_X1 U183 ( .A1(n86), .A2(n149), .ZN(n88) );
  NAND2_X1 U184 ( .A1(n749), .A2(AReg_DP[4]), .ZN(n184) );
  INV_X1 U185 ( .A(n184), .ZN(n87) );
  AND2_X1 U186 ( .A1(n768), .A2(AReg_DP[5]), .ZN(n179) );
  AOI211_X1 U187 ( .C1(n89), .C2(n88), .A(n87), .B(n179), .ZN(n91) );
  NOR2_X1 U188 ( .A1(n750), .A2(AReg_DP[6]), .ZN(n148) );
  AOI22_X1 U189 ( .A1(BReg_DP[5]), .A2(n760), .B1(n732), .B2(BReg_DP[7]), .ZN(
        n163) );
  INV_X1 U190 ( .A(n163), .ZN(n90) );
  NOR3_X1 U191 ( .A1(n91), .A2(n148), .A3(n90), .ZN(n92) );
  AOI21_X1 U192 ( .B1(n94), .B2(n93), .A(n92), .ZN(n99) );
  AOI21_X1 U193 ( .B1(BReg_DP[8]), .B2(n798), .A(n95), .ZN(n98) );
  INV_X1 U194 ( .A(n101), .ZN(n96) );
  NAND3_X1 U195 ( .A1(n98), .A2(n97), .A3(n96), .ZN(n198) );
  OAI22_X1 U196 ( .A1(n101), .A2(n100), .B1(n99), .B2(n198), .ZN(n108) );
  NOR2_X1 U197 ( .A1(n757), .A2(BReg_DP[12]), .ZN(n147) );
  AND2_X1 U198 ( .A1(n753), .A2(AReg_DP[14]), .ZN(n171) );
  AND2_X1 U199 ( .A1(n755), .A2(AReg_DP[13]), .ZN(n169) );
  AOI211_X1 U200 ( .C1(n147), .C2(n102), .A(n171), .B(n169), .ZN(n105) );
  OR3_X1 U201 ( .A1(n105), .A2(n104), .A3(n103), .ZN(n106) );
  NAND2_X1 U202 ( .A1(n751), .A2(AReg_DP[15]), .ZN(n173) );
  NAND2_X1 U203 ( .A1(n106), .A2(n173), .ZN(n107) );
  AOI221_X1 U204 ( .B1(n150), .B2(n194), .C1(n108), .C2(n194), .A(n107), .ZN(
        n118) );
  NAND2_X1 U205 ( .A1(n765), .A2(BReg_DP[19]), .ZN(n113) );
  INV_X1 U206 ( .A(n113), .ZN(n109) );
  AOI21_X1 U207 ( .B1(BReg_DP[18]), .B2(n770), .A(n109), .ZN(n115) );
  OR2_X1 U208 ( .A1(n756), .A2(AReg_DP[17]), .ZN(n110) );
  OAI211_X1 U209 ( .C1(AReg_DP[16]), .C2(n789), .A(n115), .B(n110), .ZN(n195)
         );
  INV_X1 U210 ( .A(n110), .ZN(n112) );
  NAND2_X1 U211 ( .A1(n789), .A2(AReg_DP[16]), .ZN(n172) );
  AND2_X1 U212 ( .A1(n756), .A2(AReg_DP[17]), .ZN(n178) );
  INV_X1 U213 ( .A(n178), .ZN(n111) );
  OAI21_X1 U214 ( .B1(n112), .B2(n172), .A(n111), .ZN(n114) );
  NOR2_X1 U215 ( .A1(n770), .A2(BReg_DP[18]), .ZN(n141) );
  AOI22_X1 U216 ( .A1(n115), .A2(n114), .B1(n141), .B2(n113), .ZN(n117) );
  AND2_X1 U217 ( .A1(n815), .A2(AReg_DP[19]), .ZN(n144) );
  INV_X1 U218 ( .A(n144), .ZN(n116) );
  OAI211_X1 U219 ( .C1(n118), .C2(n195), .A(n117), .B(n116), .ZN(n126) );
  NOR2_X1 U220 ( .A1(n793), .A2(BReg_DP[20]), .ZN(n145) );
  OAI21_X1 U221 ( .B1(n145), .B2(AReg_DP[21]), .A(n791), .ZN(n121) );
  NAND2_X1 U222 ( .A1(n145), .A2(AReg_DP[21]), .ZN(n120) );
  AOI21_X1 U223 ( .B1(n121), .B2(n120), .A(n119), .ZN(n125) );
  NOR2_X1 U224 ( .A1(n796), .A2(BReg_DP[22]), .ZN(n146) );
  NAND2_X1 U225 ( .A1(n146), .A2(n122), .ZN(n123) );
  NAND2_X1 U226 ( .A1(n807), .A2(AReg_DP[23]), .ZN(n152) );
  NAND2_X1 U227 ( .A1(n123), .A2(n152), .ZN(n124) );
  AOI211_X1 U228 ( .C1(n191), .C2(n126), .A(n125), .B(n124), .ZN(n137) );
  NOR2_X1 U229 ( .A1(n800), .A2(AReg_DP[27]), .ZN(n128) );
  AOI21_X1 U230 ( .B1(BReg_DP[26]), .B2(n771), .A(n128), .ZN(n133) );
  NOR2_X1 U231 ( .A1(n795), .A2(BReg_DP[24]), .ZN(n160) );
  NAND2_X1 U232 ( .A1(n803), .A2(BReg_DP[25]), .ZN(n132) );
  NAND2_X1 U233 ( .A1(n160), .A2(n132), .ZN(n127) );
  NAND2_X1 U234 ( .A1(n808), .A2(AReg_DP[25]), .ZN(n175) );
  NAND2_X1 U235 ( .A1(n127), .A2(n175), .ZN(n131) );
  NOR2_X1 U236 ( .A1(n794), .A2(BReg_DP[27]), .ZN(n143) );
  NOR2_X1 U237 ( .A1(n771), .A2(BReg_DP[26]), .ZN(n161) );
  INV_X1 U238 ( .A(n161), .ZN(n129) );
  NOR2_X1 U239 ( .A1(n129), .A2(n128), .ZN(n130) );
  AOI211_X1 U240 ( .C1(n133), .C2(n131), .A(n143), .B(n130), .ZN(n136) );
  OAI211_X1 U241 ( .C1(AReg_DP[24]), .C2(n812), .A(n133), .B(n132), .ZN(n196)
         );
  AOI21_X1 U242 ( .B1(BReg_DP[28]), .B2(n797), .A(n134), .ZN(n164) );
  NAND2_X1 U243 ( .A1(n164), .A2(n174), .ZN(n135) );
  AOI221_X1 U244 ( .B1(n137), .B2(n136), .C1(n196), .C2(n136), .A(n135), .ZN(
        n138) );
  AOI211_X1 U245 ( .C1(n174), .C2(n140), .A(n139), .B(n138), .ZN(n202) );
  INV_X1 U246 ( .A(n141), .ZN(n142) );
  OAI21_X1 U247 ( .B1(BReg_DP[21]), .B2(n748), .A(n142), .ZN(n159) );
  NOR4_X1 U248 ( .A1(n146), .A2(n145), .A3(n144), .A4(n143), .ZN(n157) );
  NOR4_X1 U249 ( .A1(n150), .A2(n149), .A3(n148), .A4(n147), .ZN(n156) );
  AND3_X1 U250 ( .A1(n153), .A2(n152), .A3(n151), .ZN(n155) );
  NAND4_X1 U251 ( .A1(n157), .A2(n156), .A3(n155), .A4(n154), .ZN(n158) );
  NOR4_X1 U252 ( .A1(n161), .A2(n160), .A3(n159), .A4(n158), .ZN(n193) );
  NAND3_X1 U253 ( .A1(n164), .A2(n163), .A3(n162), .ZN(n167) );
  XOR2_X1 U254 ( .A(BReg_DP[0]), .B(AReg_DP[0]), .Z(n166) );
  XOR2_X1 U255 ( .A(BReg_DP[1]), .B(AReg_DP[1]), .Z(n165) );
  NOR3_X1 U256 ( .A1(n167), .A2(n166), .A3(n165), .ZN(n192) );
  NOR4_X1 U257 ( .A1(n171), .A2(n170), .A3(n169), .A4(n168), .ZN(n182) );
  NAND3_X1 U258 ( .A1(n174), .A2(n173), .A3(n172), .ZN(n177) );
  OAI21_X1 U259 ( .B1(BReg_DP[7]), .B2(n732), .A(n175), .ZN(n176) );
  NOR4_X1 U260 ( .A1(n179), .A2(n178), .A3(n177), .A4(n176), .ZN(n181) );
  NAND4_X1 U261 ( .A1(n183), .A2(n182), .A3(n181), .A4(n180), .ZN(n189) );
  NAND4_X1 U262 ( .A1(n187), .A2(n186), .A3(n185), .A4(n184), .ZN(n188) );
  NOR2_X1 U263 ( .A1(n189), .A2(n188), .ZN(n190) );
  AND4_X1 U264 ( .A1(n193), .A2(n192), .A3(n191), .A4(n190), .ZN(n200) );
  INV_X1 U265 ( .A(n194), .ZN(n197) );
  NOR4_X1 U266 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(n199) );
  AOI22_X1 U267 ( .A1(n200), .A2(n199), .B1(n202), .B2(CompInv_SP), .ZN(n201)
         );
  OAI21_X1 U268 ( .B1(n202), .B2(CompInv_SP), .A(n201), .ZN(n203) );
  NAND3_X1 U269 ( .A1(n204), .A2(n570), .A3(n203), .ZN(n579) );
  MUX2_X1 U270 ( .A(AReg_DP[12]), .B(n205), .S(n577), .Z(n206) );
  INV_X1 U271 ( .A(n206), .ZN(n729) );
  INV_X1 U273 ( .A(n829), .ZN(n571) );
  NAND2_X1 U274 ( .A1(n830), .A2(n821), .ZN(n582) );
  INV_X1 U277 ( .A(OpBShift_DI[5]), .ZN(n213) );
  NOR3_X1 U278 ( .A1(Cnt_DP[2]), .A2(Cnt_DP[0]), .A3(Cnt_DP[1]), .ZN(n607) );
  NAND2_X1 U279 ( .A1(n607), .A2(n813), .ZN(n590) );
  OR2_X1 U280 ( .A1(Cnt_DP[4]), .A2(n590), .ZN(n317) );
  NAND3_X1 U281 ( .A1(n830), .A2(Cnt_DP[5]), .A3(n317), .ZN(n208) );
  OAI21_X1 U282 ( .B1(n213), .B2(n594), .A(n208), .ZN(n284) );
  INV_X1 U283 ( .A(OpBShift_DI[4]), .ZN(n319) );
  INV_X1 U284 ( .A(n317), .ZN(n231) );
  AOI21_X1 U285 ( .B1(Cnt_DP[4]), .B2(n590), .A(n231), .ZN(n318) );
  NOR2_X1 U286 ( .A1(n317), .A2(Cnt_DP[5]), .ZN(n322) );
  OR2_X1 U287 ( .A1(n571), .A2(n322), .ZN(n610) );
  OAI22_X1 U288 ( .A1(n319), .A2(n594), .B1(n318), .B2(n610), .ZN(n283) );
  INV_X1 U289 ( .A(InVld_SI), .ZN(n320) );
  NOR2_X1 U290 ( .A1(n320), .A2(State_SP[1]), .ZN(n321) );
  NOR2_X1 U291 ( .A1(n321), .A2(State_SP[0]), .ZN(OutVld_SO) );
  AOI21_X1 U292 ( .B1(n322), .B2(n570), .A(OutVld_SO), .ZN(n278) );
  OAI21_X1 U293 ( .B1(n322), .B2(State_SP[1]), .A(State_SP[0]), .ZN(n323) );
  OAI21_X1 U294 ( .B1(OutRdy_SI), .B2(n805), .A(n323), .ZN(n277) );
  INV_X2 U295 ( .A(n594), .ZN(n566) );
  MUX2_X1 U296 ( .A(BReg_DP[30]), .B(OpA_DI[30]), .S(n566), .Z(n324) );
  XOR2_X1 U297 ( .A(n12), .B(n324), .Z(n576) );
  NOR2_X1 U298 ( .A1(n566), .A2(n772), .ZN(n575) );
  MUX2_X1 U299 ( .A(BReg_DP[29]), .B(OpA_DI[29]), .S(n566), .Z(n325) );
  XOR2_X1 U300 ( .A(n12), .B(n325), .Z(n381) );
  AND2_X1 U301 ( .A1(n829), .A2(AReg_DP[29]), .ZN(n380) );
  MUX2_X1 U302 ( .A(BReg_DP[28]), .B(OpA_DI[28]), .S(n566), .Z(n326) );
  XOR2_X1 U303 ( .A(n12), .B(n326), .Z(n385) );
  AND2_X1 U304 ( .A1(n829), .A2(AReg_DP[28]), .ZN(n384) );
  MUX2_X1 U305 ( .A(BReg_DP[27]), .B(OpA_DI[27]), .S(n566), .Z(n327) );
  XOR2_X1 U306 ( .A(n12), .B(n327), .Z(n389) );
  AND2_X1 U307 ( .A1(n829), .A2(AReg_DP[27]), .ZN(n388) );
  MUX2_X1 U308 ( .A(BReg_DP[26]), .B(OpA_DI[26]), .S(n566), .Z(n328) );
  XOR2_X1 U309 ( .A(n12), .B(n328), .Z(n393) );
  AND2_X1 U310 ( .A1(n829), .A2(AReg_DP[26]), .ZN(n392) );
  MUX2_X1 U311 ( .A(BReg_DP[25]), .B(OpA_DI[25]), .S(n566), .Z(n329) );
  XOR2_X1 U312 ( .A(n12), .B(n329), .Z(n397) );
  AND2_X1 U313 ( .A1(n829), .A2(AReg_DP[25]), .ZN(n396) );
  MUX2_X1 U314 ( .A(BReg_DP[24]), .B(OpA_DI[24]), .S(n566), .Z(n330) );
  XOR2_X1 U315 ( .A(n12), .B(n330), .Z(n401) );
  AND2_X1 U316 ( .A1(n829), .A2(AReg_DP[24]), .ZN(n400) );
  INV_X1 U317 ( .A(n331), .ZN(n332) );
  AOI21_X1 U318 ( .B1(n334), .B2(n333), .A(n332), .ZN(n462) );
  MUX2_X1 U319 ( .A(BReg_DP[13]), .B(OpA_DI[13]), .S(n566), .Z(n335) );
  XOR2_X1 U320 ( .A(n12), .B(n335), .Z(n337) );
  AND2_X1 U321 ( .A1(n594), .A2(AReg_DP[13]), .ZN(n336) );
  NOR2_X1 U322 ( .A1(n337), .A2(n336), .ZN(n458) );
  NAND2_X1 U323 ( .A1(n337), .A2(n336), .ZN(n459) );
  OAI21_X1 U324 ( .B1(n462), .B2(n458), .A(n459), .ZN(n456) );
  MUX2_X1 U325 ( .A(BReg_DP[14]), .B(OpA_DI[14]), .S(n566), .Z(n338) );
  XOR2_X1 U326 ( .A(n12), .B(n338), .Z(n340) );
  AND2_X1 U327 ( .A1(n830), .A2(AReg_DP[14]), .ZN(n339) );
  OR2_X1 U328 ( .A1(n340), .A2(n339), .ZN(n454) );
  NAND2_X1 U329 ( .A1(n340), .A2(n339), .ZN(n453) );
  INV_X1 U330 ( .A(n453), .ZN(n341) );
  AOI21_X1 U331 ( .B1(n456), .B2(n454), .A(n341), .ZN(n451) );
  MUX2_X1 U332 ( .A(BReg_DP[15]), .B(OpA_DI[15]), .S(n566), .Z(n342) );
  XOR2_X1 U333 ( .A(n12), .B(n342), .Z(n344) );
  AND2_X1 U334 ( .A1(n594), .A2(AReg_DP[15]), .ZN(n343) );
  NOR2_X1 U335 ( .A1(n344), .A2(n343), .ZN(n447) );
  NAND2_X1 U336 ( .A1(n344), .A2(n343), .ZN(n448) );
  OAI21_X1 U337 ( .B1(n451), .B2(n447), .A(n448), .ZN(n445) );
  MUX2_X1 U338 ( .A(BReg_DP[16]), .B(OpA_DI[16]), .S(n566), .Z(n345) );
  XOR2_X1 U339 ( .A(n12), .B(n345), .Z(n347) );
  AND2_X1 U340 ( .A1(n829), .A2(AReg_DP[16]), .ZN(n346) );
  OR2_X1 U341 ( .A1(n347), .A2(n346), .ZN(n443) );
  NAND2_X1 U342 ( .A1(n347), .A2(n346), .ZN(n442) );
  INV_X1 U343 ( .A(n442), .ZN(n348) );
  AOI21_X1 U344 ( .B1(n445), .B2(n443), .A(n348), .ZN(n440) );
  MUX2_X1 U345 ( .A(BReg_DP[17]), .B(OpA_DI[17]), .S(n566), .Z(n349) );
  XOR2_X1 U346 ( .A(n12), .B(n349), .Z(n351) );
  AND2_X1 U347 ( .A1(n594), .A2(AReg_DP[17]), .ZN(n350) );
  NOR2_X1 U348 ( .A1(n351), .A2(n350), .ZN(n436) );
  NAND2_X1 U349 ( .A1(n351), .A2(n350), .ZN(n437) );
  OAI21_X1 U350 ( .B1(n440), .B2(n436), .A(n437), .ZN(n434) );
  MUX2_X1 U351 ( .A(BReg_DP[18]), .B(OpA_DI[18]), .S(n566), .Z(n352) );
  XOR2_X1 U352 ( .A(n12), .B(n352), .Z(n354) );
  AND2_X1 U353 ( .A1(n594), .A2(AReg_DP[18]), .ZN(n353) );
  OR2_X1 U354 ( .A1(n354), .A2(n353), .ZN(n432) );
  NAND2_X1 U355 ( .A1(n354), .A2(n353), .ZN(n431) );
  INV_X1 U356 ( .A(n431), .ZN(n355) );
  AOI21_X1 U357 ( .B1(n434), .B2(n432), .A(n355), .ZN(n429) );
  MUX2_X1 U358 ( .A(BReg_DP[19]), .B(OpA_DI[19]), .S(n566), .Z(n356) );
  XOR2_X1 U359 ( .A(n12), .B(n356), .Z(n358) );
  AND2_X1 U360 ( .A1(n594), .A2(AReg_DP[19]), .ZN(n357) );
  NOR2_X1 U361 ( .A1(n358), .A2(n357), .ZN(n425) );
  NAND2_X1 U362 ( .A1(n358), .A2(n357), .ZN(n426) );
  OAI21_X1 U363 ( .B1(n429), .B2(n425), .A(n426), .ZN(n423) );
  MUX2_X1 U364 ( .A(BReg_DP[20]), .B(OpA_DI[20]), .S(n566), .Z(n359) );
  XOR2_X1 U365 ( .A(n12), .B(n359), .Z(n361) );
  AND2_X1 U366 ( .A1(n829), .A2(AReg_DP[20]), .ZN(n360) );
  OR2_X1 U367 ( .A1(n361), .A2(n360), .ZN(n421) );
  NAND2_X1 U368 ( .A1(n361), .A2(n360), .ZN(n420) );
  INV_X1 U369 ( .A(n420), .ZN(n362) );
  AOI21_X1 U370 ( .B1(n423), .B2(n421), .A(n362), .ZN(n418) );
  MUX2_X1 U371 ( .A(BReg_DP[21]), .B(OpA_DI[21]), .S(n566), .Z(n363) );
  XOR2_X1 U372 ( .A(n12), .B(n363), .Z(n365) );
  NOR2_X1 U373 ( .A1(n566), .A2(n748), .ZN(n364) );
  NOR2_X1 U374 ( .A1(n365), .A2(n364), .ZN(n414) );
  NAND2_X1 U375 ( .A1(n365), .A2(n364), .ZN(n415) );
  OAI21_X1 U376 ( .B1(n418), .B2(n414), .A(n415), .ZN(n412) );
  MUX2_X1 U377 ( .A(BReg_DP[22]), .B(OpA_DI[22]), .S(n566), .Z(n366) );
  XOR2_X1 U378 ( .A(n12), .B(n366), .Z(n368) );
  AND2_X1 U379 ( .A1(n594), .A2(AReg_DP[22]), .ZN(n367) );
  OR2_X1 U380 ( .A1(n368), .A2(n367), .ZN(n410) );
  NAND2_X1 U381 ( .A1(n368), .A2(n367), .ZN(n409) );
  INV_X1 U382 ( .A(n409), .ZN(n369) );
  MUX2_X1 U383 ( .A(BReg_DP[23]), .B(OpA_DI[23]), .S(n566), .Z(n370) );
  XOR2_X1 U384 ( .A(n12), .B(n370), .Z(n405) );
  AND2_X1 U385 ( .A1(n830), .A2(AReg_DP[23]), .ZN(n403) );
  NOR2_X1 U386 ( .A1(n405), .A2(n403), .ZN(n373) );
  NAND2_X1 U387 ( .A1(n405), .A2(n403), .ZN(n372) );
  MUX2_X1 U388 ( .A(BReg_DP[31]), .B(OpA_DI[31]), .S(n566), .Z(n374) );
  XOR2_X1 U389 ( .A(n12), .B(n374), .Z(n376) );
  NOR2_X1 U390 ( .A1(n566), .A2(n801), .ZN(n375) );
  XNOR2_X1 U391 ( .A(n377), .B(n14), .ZN(n378) );
  MUX2_X1 U392 ( .A(AReg_DP[31]), .B(n378), .S(n577), .Z(n244) );
  FA_X1 U393 ( .A(n381), .B(n380), .CI(n379), .CO(n574), .S(n382) );
  MUX2_X1 U394 ( .A(AReg_DP[29]), .B(n382), .S(n577), .Z(n214) );
  FA_X1 U395 ( .A(n385), .B(n384), .CI(n383), .CO(n379), .S(n386) );
  MUX2_X1 U396 ( .A(AReg_DP[28]), .B(n386), .S(n577), .Z(n215) );
  FA_X1 U397 ( .A(n389), .B(n388), .CI(n387), .CO(n383), .S(n390) );
  MUX2_X1 U398 ( .A(AReg_DP[27]), .B(n390), .S(n577), .Z(n216) );
  FA_X1 U399 ( .A(n393), .B(n392), .CI(n391), .CO(n387), .S(n394) );
  MUX2_X1 U400 ( .A(AReg_DP[26]), .B(n394), .S(n577), .Z(n217) );
  FA_X1 U401 ( .A(n397), .B(n396), .CI(n395), .CO(n391), .S(n398) );
  MUX2_X1 U402 ( .A(AReg_DP[25]), .B(n398), .S(n577), .Z(n218) );
  FA_X1 U403 ( .A(n401), .B(n400), .CI(n399), .CO(n395), .S(n402) );
  MUX2_X1 U404 ( .A(AReg_DP[24]), .B(n402), .S(n577), .Z(n219) );
  INV_X1 U405 ( .A(n403), .ZN(n404) );
  XNOR2_X1 U406 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U407 ( .A(n827), .B(n406), .ZN(n408) );
  MUX2_X1 U408 ( .A(AReg_DP[23]), .B(n408), .S(n577), .Z(n220) );
  NAND2_X1 U409 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U410 ( .A(n412), .B(n411), .ZN(n413) );
  MUX2_X1 U411 ( .A(AReg_DP[22]), .B(n413), .S(n577), .Z(n221) );
  INV_X1 U412 ( .A(n414), .ZN(n416) );
  NAND2_X1 U413 ( .A1(n416), .A2(n415), .ZN(n417) );
  XOR2_X1 U414 ( .A(n418), .B(n417), .Z(n419) );
  MUX2_X1 U415 ( .A(AReg_DP[21]), .B(n419), .S(n577), .Z(n222) );
  NAND2_X1 U416 ( .A1(n421), .A2(n420), .ZN(n422) );
  XNOR2_X1 U417 ( .A(n423), .B(n422), .ZN(n424) );
  MUX2_X1 U418 ( .A(AReg_DP[20]), .B(n424), .S(n577), .Z(n223) );
  INV_X1 U419 ( .A(n425), .ZN(n427) );
  NAND2_X1 U420 ( .A1(n427), .A2(n426), .ZN(n428) );
  XOR2_X1 U421 ( .A(n826), .B(n428), .Z(n430) );
  MUX2_X1 U422 ( .A(AReg_DP[19]), .B(n430), .S(n577), .Z(n224) );
  NAND2_X1 U423 ( .A1(n432), .A2(n431), .ZN(n433) );
  XNOR2_X1 U424 ( .A(n434), .B(n433), .ZN(n435) );
  MUX2_X1 U425 ( .A(AReg_DP[18]), .B(n435), .S(n577), .Z(n225) );
  INV_X1 U426 ( .A(n436), .ZN(n438) );
  NAND2_X1 U427 ( .A1(n438), .A2(n437), .ZN(n439) );
  XOR2_X1 U428 ( .A(n440), .B(n439), .Z(n441) );
  MUX2_X1 U429 ( .A(AReg_DP[17]), .B(n441), .S(n577), .Z(n226) );
  NAND2_X1 U430 ( .A1(n443), .A2(n442), .ZN(n444) );
  XNOR2_X1 U431 ( .A(n445), .B(n444), .ZN(n446) );
  MUX2_X1 U432 ( .A(AReg_DP[16]), .B(n446), .S(n577), .Z(n227) );
  INV_X1 U433 ( .A(n447), .ZN(n449) );
  NAND2_X1 U434 ( .A1(n449), .A2(n448), .ZN(n450) );
  XOR2_X1 U435 ( .A(n451), .B(n450), .Z(n452) );
  MUX2_X1 U436 ( .A(AReg_DP[15]), .B(n452), .S(n577), .Z(n228) );
  NAND2_X1 U437 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U438 ( .A(n456), .B(n455), .ZN(n457) );
  MUX2_X1 U439 ( .A(AReg_DP[14]), .B(n457), .S(n577), .Z(n229) );
  INV_X1 U440 ( .A(n458), .ZN(n460) );
  NAND2_X1 U441 ( .A1(n460), .A2(n459), .ZN(n461) );
  XOR2_X1 U442 ( .A(n462), .B(n461), .Z(n463) );
  MUX2_X1 U443 ( .A(AReg_DP[13]), .B(n463), .S(n577), .Z(n230) );
  INV_X1 U444 ( .A(n464), .ZN(n466) );
  NAND2_X1 U445 ( .A1(n466), .A2(n465), .ZN(n467) );
  XOR2_X1 U446 ( .A(n468), .B(n467), .Z(n469) );
  MUX2_X1 U447 ( .A(AReg_DP[11]), .B(n469), .S(n577), .Z(n232) );
  NAND2_X1 U448 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U449 ( .A(n473), .B(n472), .ZN(n474) );
  MUX2_X1 U450 ( .A(AReg_DP[10]), .B(n474), .S(n577), .Z(n233) );
  INV_X1 U451 ( .A(n475), .ZN(n477) );
  NAND2_X1 U452 ( .A1(n477), .A2(n476), .ZN(n478) );
  XOR2_X1 U453 ( .A(n828), .B(n478), .Z(n480) );
  MUX2_X1 U454 ( .A(AReg_DP[9]), .B(n480), .S(n577), .Z(n234) );
  INV_X1 U455 ( .A(n481), .ZN(n492) );
  OAI21_X1 U456 ( .B1(n492), .B2(n488), .A(n489), .ZN(n486) );
  INV_X1 U457 ( .A(n482), .ZN(n484) );
  NAND2_X1 U458 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U459 ( .A(n486), .B(n485), .ZN(n487) );
  MUX2_X1 U460 ( .A(AReg_DP[8]), .B(n487), .S(n577), .Z(n235) );
  INV_X1 U461 ( .A(n488), .ZN(n490) );
  NAND2_X1 U462 ( .A1(n490), .A2(n489), .ZN(n491) );
  XOR2_X1 U463 ( .A(n492), .B(n491), .Z(n493) );
  MUX2_X1 U464 ( .A(AReg_DP[7]), .B(n493), .S(n577), .Z(n236) );
  INV_X1 U465 ( .A(n494), .ZN(n520) );
  AOI21_X1 U466 ( .B1(n520), .B2(n496), .A(n495), .ZN(n507) );
  OAI21_X1 U467 ( .B1(n507), .B2(n503), .A(n504), .ZN(n501) );
  INV_X1 U468 ( .A(n497), .ZN(n499) );
  NAND2_X1 U469 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U470 ( .A(n501), .B(n500), .ZN(n502) );
  MUX2_X1 U471 ( .A(AReg_DP[6]), .B(n502), .S(n577), .Z(n237) );
  INV_X1 U472 ( .A(n503), .ZN(n505) );
  NAND2_X1 U473 ( .A1(n505), .A2(n504), .ZN(n506) );
  XOR2_X1 U474 ( .A(n507), .B(n506), .Z(n508) );
  MUX2_X1 U475 ( .A(AReg_DP[5]), .B(n508), .S(n577), .Z(n238) );
  INV_X1 U476 ( .A(n509), .ZN(n518) );
  INV_X1 U477 ( .A(n517), .ZN(n510) );
  AOI21_X1 U478 ( .B1(n520), .B2(n518), .A(n510), .ZN(n515) );
  INV_X1 U479 ( .A(n511), .ZN(n513) );
  NAND2_X1 U480 ( .A1(n513), .A2(n512), .ZN(n514) );
  XOR2_X1 U481 ( .A(n515), .B(n514), .Z(n516) );
  MUX2_X1 U482 ( .A(AReg_DP[4]), .B(n516), .S(n577), .Z(n239) );
  NAND2_X1 U483 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U484 ( .A(n520), .B(n519), .ZN(n521) );
  MUX2_X1 U485 ( .A(AReg_DP[3]), .B(n521), .S(n577), .Z(n240) );
  INV_X1 U486 ( .A(n522), .ZN(n532) );
  OAI21_X1 U487 ( .B1(n529), .B2(n532), .A(n530), .ZN(n527) );
  INV_X1 U488 ( .A(n523), .ZN(n525) );
  NAND2_X1 U489 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U490 ( .A(n527), .B(n526), .ZN(n528) );
  MUX2_X1 U491 ( .A(AReg_DP[2]), .B(n528), .S(n577), .Z(n241) );
  INV_X1 U492 ( .A(n529), .ZN(n531) );
  NAND2_X1 U493 ( .A1(n531), .A2(n530), .ZN(n533) );
  XOR2_X1 U494 ( .A(n533), .B(n532), .Z(n534) );
  MUX2_X1 U495 ( .A(AReg_DP[1]), .B(n534), .S(n577), .Z(n242) );
  NAND2_X1 U496 ( .A1(n12), .A2(n21), .ZN(n537) );
  XNOR2_X1 U497 ( .A(n537), .B(n536), .ZN(n538) );
  MUX2_X1 U498 ( .A(AReg_DP[0]), .B(n538), .S(n577), .Z(n243) );
  FA_X1 U561 ( .A(n576), .B(n575), .CI(n574), .CO(n377), .S(n578) );
  MUX2_X1 U562 ( .A(AReg_DP[30]), .B(n578), .S(n577), .Z(n212) );
  INV_X1 U598 ( .A(OpBIsZero_SI), .ZN(n585) );
  OAI21_X1 U599 ( .B1(n585), .B2(OpCode_SI[1]), .A(n566), .ZN(n587) );
  NAND2_X1 U601 ( .A1(OpBShift_DI[0]), .A2(n566), .ZN(n589) );
  OAI21_X1 U602 ( .B1(Cnt_DP[0]), .B2(n610), .A(n589), .ZN(n279) );
  INV_X1 U603 ( .A(OpBShift_DI[3]), .ZN(n595) );
  INV_X1 U604 ( .A(n607), .ZN(n592) );
  INV_X1 U605 ( .A(n590), .ZN(n591) );
  AOI21_X1 U606 ( .B1(n592), .B2(Cnt_DP[3]), .A(n591), .ZN(n593) );
  OAI22_X1 U607 ( .A1(n595), .A2(n594), .B1(n593), .B2(n610), .ZN(n282) );
  NAND2_X1 U608 ( .A1(AReg_DP[1]), .A2(RemSel_SP), .ZN(n596) );
  OAI21_X1 U609 ( .B1(n731), .B2(n7), .A(n596), .ZN(n598) );
  INV_X1 U610 ( .A(Res_DO[0]), .ZN(n601) );
  INV_X1 U611 ( .A(n598), .ZN(n600) );
  MUX2_X1 U612 ( .A(n598), .B(n597), .S(ResInv_SP), .Z(Res_DO[1]) );
  NAND2_X1 U613 ( .A1(AReg_DP[2]), .A2(n6), .ZN(n599) );
  OAI21_X1 U614 ( .B1(n730), .B2(n6), .A(n599), .ZN(n603) );
  INV_X1 U616 ( .A(n603), .ZN(n612) );
  MUX2_X1 U617 ( .A(n603), .B(n602), .S(ResInv_SP), .Z(Res_DO[2]) );
  NOR2_X1 U618 ( .A1(Cnt_DP[0]), .A2(Cnt_DP[1]), .ZN(n606) );
  AOI21_X1 U619 ( .B1(Cnt_DP[1]), .B2(Cnt_DP[0]), .A(n606), .ZN(n605) );
  NAND2_X1 U620 ( .A1(OpBShift_DI[1]), .A2(n566), .ZN(n604) );
  OAI21_X1 U621 ( .B1(n605), .B2(n610), .A(n604), .ZN(n280) );
  INV_X1 U622 ( .A(n606), .ZN(n608) );
  AOI21_X1 U623 ( .B1(Cnt_DP[2]), .B2(n608), .A(n607), .ZN(n611) );
  NAND2_X1 U624 ( .A1(OpBShift_DI[2]), .A2(n566), .ZN(n609) );
  OAI21_X1 U625 ( .B1(n611), .B2(n610), .A(n609), .ZN(n281) );
  MUX2_X1 U626 ( .A(ResReg_DP_rev[3]), .B(AReg_DP[3]), .S(n1), .Z(n614) );
  INV_X1 U627 ( .A(n614), .ZN(n616) );
  MUX2_X1 U628 ( .A(n615), .B(n614), .S(n764), .Z(Res_DO[3]) );
  HA_X1 U629 ( .A(n617), .B(n616), .CO(n621), .S(n615) );
  MUX2_X1 U630 ( .A(ResReg_DP_rev[4]), .B(AReg_DP[4]), .S(n2), .Z(n618) );
  INV_X1 U631 ( .A(n618), .ZN(n620) );
  MUX2_X1 U632 ( .A(n619), .B(n618), .S(n764), .Z(Res_DO[4]) );
  MUX2_X1 U633 ( .A(ResReg_DP_rev[5]), .B(AReg_DP[5]), .S(n1), .Z(n622) );
  INV_X1 U634 ( .A(n622), .ZN(n624) );
  MUX2_X1 U635 ( .A(n623), .B(n622), .S(n764), .Z(Res_DO[5]) );
  MUX2_X1 U637 ( .A(ResReg_DP_rev[6]), .B(AReg_DP[6]), .S(n1), .Z(n626) );
  INV_X1 U638 ( .A(n626), .ZN(n628) );
  XNOR2_X1 U639 ( .A(n629), .B(n626), .ZN(n627) );
  MUX2_X1 U640 ( .A(n627), .B(n626), .S(n764), .Z(Res_DO[6]) );
  MUX2_X1 U641 ( .A(ResReg_DP_rev[7]), .B(AReg_DP[7]), .S(n2), .Z(n630) );
  INV_X1 U642 ( .A(n630), .ZN(n632) );
  MUX2_X1 U643 ( .A(n631), .B(n630), .S(n764), .Z(Res_DO[7]) );
  HA_X1 U644 ( .A(n633), .B(n632), .CO(n637), .S(n631) );
  MUX2_X1 U645 ( .A(ResReg_DP_rev[8]), .B(AReg_DP[8]), .S(n5), .Z(n634) );
  INV_X1 U646 ( .A(n634), .ZN(n636) );
  MUX2_X1 U647 ( .A(n635), .B(n634), .S(n764), .Z(Res_DO[8]) );
  MUX2_X1 U648 ( .A(ResReg_DP_rev[9]), .B(AReg_DP[9]), .S(n2), .Z(n638) );
  INV_X1 U649 ( .A(n638), .ZN(n640) );
  MUX2_X1 U650 ( .A(n639), .B(n638), .S(n764), .Z(Res_DO[9]) );
  MUX2_X1 U652 ( .A(ResReg_DP_rev[10]), .B(AReg_DP[10]), .S(n5), .Z(n642) );
  INV_X1 U653 ( .A(n642), .ZN(n644) );
  XNOR2_X1 U654 ( .A(n645), .B(n642), .ZN(n643) );
  MUX2_X1 U655 ( .A(n643), .B(n642), .S(n764), .Z(Res_DO[10]) );
  MUX2_X1 U656 ( .A(ResReg_DP_rev[11]), .B(AReg_DP[11]), .S(n5), .Z(n646) );
  INV_X1 U657 ( .A(n646), .ZN(n648) );
  MUX2_X1 U658 ( .A(n647), .B(n646), .S(n764), .Z(Res_DO[11]) );
  HA_X1 U659 ( .A(n649), .B(n648), .CO(n653), .S(n647) );
  MUX2_X1 U660 ( .A(ResReg_DP_rev[12]), .B(AReg_DP[12]), .S(n6), .Z(n650) );
  INV_X1 U661 ( .A(n650), .ZN(n652) );
  MUX2_X1 U662 ( .A(n651), .B(n650), .S(n764), .Z(Res_DO[12]) );
  MUX2_X1 U663 ( .A(ResReg_DP_rev[13]), .B(AReg_DP[13]), .S(n7), .Z(n654) );
  INV_X1 U664 ( .A(n654), .ZN(n656) );
  MUX2_X1 U665 ( .A(n655), .B(n654), .S(n764), .Z(Res_DO[13]) );
  MUX2_X1 U667 ( .A(ResReg_DP_rev[14]), .B(AReg_DP[14]), .S(n2), .Z(n658) );
  INV_X1 U668 ( .A(n658), .ZN(n660) );
  MUX2_X1 U669 ( .A(n659), .B(n658), .S(n764), .Z(Res_DO[14]) );
  MUX2_X1 U670 ( .A(ResReg_DP_rev[15]), .B(AReg_DP[15]), .S(n2), .Z(n662) );
  INV_X1 U671 ( .A(n662), .ZN(n664) );
  MUX2_X1 U672 ( .A(n663), .B(n662), .S(n764), .Z(Res_DO[15]) );
  HA_X1 U673 ( .A(n665), .B(n664), .CO(n669), .S(n663) );
  MUX2_X1 U674 ( .A(ResReg_DP_rev[16]), .B(AReg_DP[16]), .S(n2), .Z(n666) );
  INV_X1 U675 ( .A(n666), .ZN(n668) );
  MUX2_X1 U676 ( .A(n667), .B(n666), .S(n764), .Z(Res_DO[16]) );
  MUX2_X1 U678 ( .A(ResReg_DP_rev[17]), .B(AReg_DP[17]), .S(n1), .Z(n670) );
  INV_X1 U679 ( .A(n670), .ZN(n672) );
  MUX2_X1 U680 ( .A(n671), .B(n670), .S(n764), .Z(Res_DO[17]) );
  HA_X1 U681 ( .A(n673), .B(n672), .CO(n677), .S(n671) );
  MUX2_X1 U682 ( .A(ResReg_DP_rev[18]), .B(AReg_DP[18]), .S(n1), .Z(n674) );
  INV_X1 U683 ( .A(n674), .ZN(n676) );
  MUX2_X1 U684 ( .A(n675), .B(n674), .S(n764), .Z(Res_DO[18]) );
  MUX2_X1 U686 ( .A(ResReg_DP_rev[19]), .B(AReg_DP[19]), .S(n2), .Z(n678) );
  INV_X1 U687 ( .A(n678), .ZN(n680) );
  MUX2_X1 U688 ( .A(n679), .B(n678), .S(n764), .Z(Res_DO[19]) );
  HA_X1 U689 ( .A(n681), .B(n680), .CO(n685), .S(n679) );
  MUX2_X1 U690 ( .A(ResReg_DP_rev[20]), .B(AReg_DP[20]), .S(n2), .Z(n682) );
  INV_X1 U691 ( .A(n682), .ZN(n684) );
  MUX2_X1 U692 ( .A(n683), .B(n682), .S(n764), .Z(Res_DO[20]) );
  MUX2_X1 U694 ( .A(ResReg_DP_rev[21]), .B(AReg_DP[21]), .S(n2), .Z(n686) );
  INV_X1 U695 ( .A(n686), .ZN(n688) );
  MUX2_X1 U696 ( .A(n687), .B(n686), .S(n764), .Z(Res_DO[21]) );
  HA_X1 U697 ( .A(n689), .B(n688), .CO(n693), .S(n687) );
  MUX2_X1 U698 ( .A(ResReg_DP_rev[22]), .B(AReg_DP[22]), .S(n5), .Z(n690) );
  INV_X1 U699 ( .A(n690), .ZN(n692) );
  MUX2_X1 U700 ( .A(n691), .B(n690), .S(n764), .Z(Res_DO[22]) );
  MUX2_X1 U702 ( .A(ResReg_DP_rev[23]), .B(AReg_DP[23]), .S(n5), .Z(n694) );
  INV_X1 U703 ( .A(n694), .ZN(n696) );
  MUX2_X1 U704 ( .A(n695), .B(n694), .S(n764), .Z(Res_DO[23]) );
  HA_X1 U705 ( .A(n697), .B(n696), .CO(n701), .S(n695) );
  MUX2_X1 U706 ( .A(ResReg_DP_rev[24]), .B(AReg_DP[24]), .S(n6), .Z(n698) );
  INV_X1 U707 ( .A(n698), .ZN(n700) );
  MUX2_X1 U708 ( .A(n699), .B(n698), .S(n764), .Z(Res_DO[24]) );
  HA_X1 U709 ( .A(n701), .B(n700), .CO(n705), .S(n699) );
  MUX2_X1 U710 ( .A(ResReg_DP_rev[25]), .B(AReg_DP[25]), .S(n7), .Z(n702) );
  INV_X1 U711 ( .A(n702), .ZN(n704) );
  MUX2_X1 U712 ( .A(n703), .B(n702), .S(n764), .Z(Res_DO[25]) );
  HA_X1 U713 ( .A(n705), .B(n704), .CO(n709), .S(n703) );
  MUX2_X1 U714 ( .A(ResReg_DP_rev[26]), .B(AReg_DP[26]), .S(n2), .Z(n706) );
  INV_X1 U715 ( .A(n706), .ZN(n708) );
  MUX2_X1 U716 ( .A(n707), .B(n706), .S(n764), .Z(Res_DO[26]) );
  MUX2_X1 U717 ( .A(ResReg_DP_rev[27]), .B(AReg_DP[27]), .S(n2), .Z(n710) );
  INV_X1 U718 ( .A(n710), .ZN(n712) );
  MUX2_X1 U719 ( .A(n711), .B(n710), .S(n764), .Z(Res_DO[27]) );
  HA_X1 U720 ( .A(n713), .B(n712), .CO(n717), .S(n711) );
  MUX2_X1 U721 ( .A(ResReg_DP_rev[28]), .B(AReg_DP[28]), .S(n2), .Z(n714) );
  INV_X1 U722 ( .A(n714), .ZN(n716) );
  MUX2_X1 U723 ( .A(n715), .B(n714), .S(n764), .Z(Res_DO[28]) );
  MUX2_X1 U724 ( .A(ResReg_DP_rev[29]), .B(AReg_DP[29]), .S(n1), .Z(n718) );
  INV_X1 U725 ( .A(n718), .ZN(n720) );
  MUX2_X1 U726 ( .A(n719), .B(n718), .S(n764), .Z(Res_DO[29]) );
  HA_X1 U727 ( .A(n721), .B(n720), .CO(n724), .S(n719) );
  MUX2_X1 U728 ( .A(ResReg_DP_rev[30]), .B(AReg_DP[30]), .S(n1), .Z(n722) );
  INV_X1 U729 ( .A(n722), .ZN(n725) );
  XNOR2_X1 U730 ( .A(n724), .B(n722), .ZN(n723) );
  MUX2_X1 U731 ( .A(n723), .B(n722), .S(n764), .Z(Res_DO[30]) );
  AND2_X1 U732 ( .A1(n725), .A2(n724), .ZN(n726) );
  MUX2_X1 U733 ( .A(ResReg_DP_rev[31]), .B(AReg_DP[31]), .S(n2), .Z(n727) );
  XNOR2_X1 U734 ( .A(n726), .B(n727), .ZN(n728) );
  MUX2_X1 U735 ( .A(n728), .B(n727), .S(n764), .Z(Res_DO[31]) );
  SDFFR_X1 Cnt_DP_reg_0_ ( .D(n279), .SI(1'b0), .SE(1'b0), .CK(Clk_CI), .RN(
        Rst_RBI), .Q(Cnt_DP[0]) );
  SDFFR_X1 State_SP_reg_1_ ( .D(n277), .SI(1'b0), .SE(1'b0), .CK(n1090), .RN(
        Rst_RBI), .Q(State_SP[1]), .QN(n805) );
  SDFFR_X1 State_SP_reg_0_ ( .D(n278), .SI(1'b0), .SE(1'b0), .CK(Clk_CI), .RN(
        Rst_RBI), .Q(State_SP[0]), .QN(n802) );
  SDFFR_X1 Cnt_DP_reg_5_ ( .D(n284), .SI(1'b0), .SE(1'b0), .CK(n1090), .RN(
        Rst_RBI), .Q(Cnt_DP[5]) );
  SDFFR_X1 Cnt_DP_reg_4_ ( .D(n283), .SI(1'b0), .SE(1'b0), .CK(n1090), .RN(
        Rst_RBI), .Q(Cnt_DP[4]) );
  SDFFR_X1 Cnt_DP_reg_3_ ( .D(n282), .SI(1'b0), .SE(1'b0), .CK(n1090), .RN(
        Rst_RBI), .Q(Cnt_DP[3]), .QN(n813) );
  SDFFR_X1 Cnt_DP_reg_2_ ( .D(n281), .SI(1'b0), .SE(1'b0), .CK(n1090), .RN(
        Rst_RBI), .Q(Cnt_DP[2]) );
  SDFFR_X1 Cnt_DP_reg_1_ ( .D(n280), .SI(1'b0), .SE(1'b0), .CK(n1090), .RN(
        Rst_RBI), .Q(Cnt_DP[1]) );
  SDFFR_X1 BReg_DP_reg_31_ ( .D(n1096), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[31]), .QN(n790) );
  SDFFR_X1 BReg_DP_reg_30_ ( .D(n1097), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[30]), .QN(n810) );
  SDFFR_X1 BReg_DP_reg_29_ ( .D(n1098), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[29]), .QN(n773) );
  SDFFR_X1 BReg_DP_reg_28_ ( .D(n1099), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[28]), .QN(n809) );
  SDFFR_X1 BReg_DP_reg_27_ ( .D(n1100), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[27]), .QN(n800) );
  SDFFR_X1 BReg_DP_reg_26_ ( .D(n1101), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[26]), .QN(n825) );
  SDFFR_X1 BReg_DP_reg_25_ ( .D(n1102), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[25]), .QN(n808) );
  SDFFR_X1 BReg_DP_reg_23_ ( .D(n1103), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[23]), .QN(n807) );
  SDFFR_X1 BReg_DP_reg_22_ ( .D(n1104), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[22]), .QN(n811) );
  SDFFR_X1 BReg_DP_reg_21_ ( .D(n1105), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[21]), .QN(n791) );
  SDFFR_X1 BReg_DP_reg_20_ ( .D(n1106), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[20]), .QN(n799) );
  SDFFR_X1 BReg_DP_reg_19_ ( .D(n1107), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[19]), .QN(n815) );
  SDFFR_X1 BReg_DP_reg_18_ ( .D(n1108), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[18]) );
  SDFFR_X1 BReg_DP_reg_17_ ( .D(n1109), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[17]), .QN(n756) );
  SDFFR_X1 BReg_DP_reg_16_ ( .D(n1110), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[16]), .QN(n789) );
  SDFFR_X1 BReg_DP_reg_15_ ( .D(n1111), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[15]), .QN(n751) );
  SDFFR_X1 BReg_DP_reg_14_ ( .D(n1112), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[14]), .QN(n753) );
  SDFFR_X1 BReg_DP_reg_13_ ( .D(n1113), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[13]), .QN(n755) );
  SDFFR_X1 BReg_DP_reg_12_ ( .D(n1114), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[12]), .QN(n759) );
  SDFFR_X1 BReg_DP_reg_11_ ( .D(n1115), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[11]), .QN(n758) );
  SDFFR_X1 BReg_DP_reg_10_ ( .D(n1116), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[10]), .QN(n769) );
  SDFFR_X1 BReg_DP_reg_9_ ( .D(n1117), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[9]), .QN(n733) );
  SDFFR_X1 BReg_DP_reg_8_ ( .D(n1118), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[8]), .QN(n761) );
  SDFFR_X1 BReg_DP_reg_7_ ( .D(n1119), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[7]), .QN(n824) );
  SDFFR_X1 BReg_DP_reg_6_ ( .D(n1120), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[6]), .QN(n750) );
  SDFFR_X1 BReg_DP_reg_5_ ( .D(n1121), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[5]), .QN(n768) );
  SDFFR_X1 BReg_DP_reg_4_ ( .D(n1122), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[4]), .QN(n749) );
  SDFFR_X1 BReg_DP_reg_3_ ( .D(n1123), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[3]), .QN(n766) );
  SDFFR_X1 BReg_DP_reg_2_ ( .D(n1124), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[2]), .QN(n767) );
  SDFFR_X1 BReg_DP_reg_1_ ( .D(n1125), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[1]), .QN(n752) );
  SDFFR_X1 BReg_DP_reg_0_ ( .D(n1126), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[0]) );
  SDFFR_X1 ResReg_DP_reg_31_ ( .D(n1127), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[0]), .QN(n788) );
  SDFFR_X1 ResReg_DP_reg_30_ ( .D(n1128), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .QN(n731) );
  SDFFR_X1 ResReg_DP_reg_29_ ( .D(n1129), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .QN(n730) );
  SDFFR_X1 ResReg_DP_reg_28_ ( .D(n1130), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[3]), .QN(n774) );
  SDFFR_X1 ResReg_DP_reg_27_ ( .D(n1131), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[4]), .QN(n734) );
  SDFFR_X1 ResReg_DP_reg_26_ ( .D(n1132), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[5]), .QN(n775) );
  SDFFR_X1 ResReg_DP_reg_25_ ( .D(n1133), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[6]), .QN(n735) );
  SDFFR_X1 ResReg_DP_reg_24_ ( .D(n1134), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[7]), .QN(n776) );
  SDFFR_X1 ResReg_DP_reg_23_ ( .D(n1135), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[8]), .QN(n736) );
  SDFFR_X1 ResReg_DP_reg_22_ ( .D(n1136), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[9]), .QN(n777) );
  SDFFR_X1 ResReg_DP_reg_21_ ( .D(n1137), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[10]), .QN(n737) );
  SDFFR_X1 ResReg_DP_reg_20_ ( .D(n1138), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[11]), .QN(n778) );
  SDFFR_X1 ResReg_DP_reg_19_ ( .D(n1139), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[12]), .QN(n738) );
  SDFFR_X1 ResReg_DP_reg_18_ ( .D(n1140), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[13]), .QN(n779) );
  SDFFR_X1 ResReg_DP_reg_17_ ( .D(n1141), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[14]), .QN(n739) );
  SDFFR_X1 ResReg_DP_reg_16_ ( .D(n1142), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[15]), .QN(n780) );
  SDFFR_X1 ResReg_DP_reg_15_ ( .D(n1143), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[16]), .QN(n740) );
  SDFFR_X1 ResReg_DP_reg_14_ ( .D(n1144), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[17]), .QN(n781) );
  SDFFR_X1 ResReg_DP_reg_13_ ( .D(n1145), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[18]), .QN(n741) );
  SDFFR_X1 ResReg_DP_reg_12_ ( .D(n1146), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[19]), .QN(n782) );
  SDFFR_X1 ResReg_DP_reg_11_ ( .D(n1147), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[20]), .QN(n742) );
  SDFFR_X1 ResReg_DP_reg_10_ ( .D(n1148), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[21]), .QN(n783) );
  SDFFR_X1 ResReg_DP_reg_9_ ( .D(n1149), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[22]), .QN(n743) );
  SDFFR_X1 ResReg_DP_reg_8_ ( .D(n1150), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[23]), .QN(n784) );
  SDFFR_X1 ResReg_DP_reg_7_ ( .D(n1151), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[24]), .QN(n744) );
  SDFFR_X1 ResReg_DP_reg_6_ ( .D(n1152), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[25]), .QN(n785) );
  SDFFR_X1 ResReg_DP_reg_5_ ( .D(n1153), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[26]), .QN(n745) );
  SDFFR_X1 ResReg_DP_reg_4_ ( .D(n1154), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[27]), .QN(n786) );
  SDFFR_X1 ResReg_DP_reg_3_ ( .D(n1155), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[28]), .QN(n746) );
  SDFFR_X1 ResReg_DP_reg_2_ ( .D(n1156), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[29]), .QN(n787) );
  SDFFR_X1 ResReg_DP_reg_1_ ( .D(n1157), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[30]), .QN(n747) );
  SDFFR_X1 ResReg_DP_reg_0_ ( .D(n1158), .SI(1'b0), .SE(1'b0), .CK(n1159), 
        .RN(Rst_RBI), .Q(ResReg_DP_rev[31]) );
  SDFFR_X1 AReg_DP_reg_31_ ( .D(n244), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[31]), .QN(n801) );
  SDFFR_X1 AReg_DP_reg_0_ ( .D(n243), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[0]) );
  SDFFR_X1 AReg_DP_reg_1_ ( .D(n242), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[1]), .QN(n754) );
  SDFFR_X1 AReg_DP_reg_2_ ( .D(n241), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[2]), .QN(n762) );
  SDFFR_X1 AReg_DP_reg_3_ ( .D(n240), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[3]), .QN(n763) );
  SDFFR_X1 AReg_DP_reg_4_ ( .D(n239), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[4]) );
  SDFFR_X1 AReg_DP_reg_5_ ( .D(n238), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[5]), .QN(n760) );
  SDFFR_X1 AReg_DP_reg_6_ ( .D(n237), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[6]) );
  SDFFR_X1 AReg_DP_reg_7_ ( .D(n236), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[7]), .QN(n732) );
  SDFFR_X1 AReg_DP_reg_8_ ( .D(n235), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[8]), .QN(n798) );
  SDFFR_X1 AReg_DP_reg_9_ ( .D(n234), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[9]) );
  SDFFR_X1 AReg_DP_reg_10_ ( .D(n233), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[10]), .QN(n806) );
  SDFFR_X1 AReg_DP_reg_11_ ( .D(n232), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[11]), .QN(n792) );
  SDFFR_X1 AReg_DP_reg_13_ ( .D(n230), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[13]) );
  SDFFR_X1 AReg_DP_reg_14_ ( .D(n229), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[14]) );
  SDFFR_X1 AReg_DP_reg_15_ ( .D(n228), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[15]) );
  SDFFR_X1 AReg_DP_reg_16_ ( .D(n227), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[16]) );
  SDFFR_X1 AReg_DP_reg_17_ ( .D(n226), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[17]) );
  SDFFR_X1 AReg_DP_reg_18_ ( .D(n225), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[18]), .QN(n770) );
  SDFFR_X1 AReg_DP_reg_19_ ( .D(n224), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[19]), .QN(n765) );
  SDFFR_X1 AReg_DP_reg_20_ ( .D(n223), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[20]), .QN(n793) );
  SDFFR_X1 AReg_DP_reg_21_ ( .D(n222), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[21]), .QN(n748) );
  SDFFR_X1 AReg_DP_reg_22_ ( .D(n221), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[22]), .QN(n796) );
  SDFFR_X1 AReg_DP_reg_23_ ( .D(n220), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[23]), .QN(n804) );
  SDFFR_X1 AReg_DP_reg_24_ ( .D(n219), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[24]), .QN(n795) );
  SDFFR_X1 AReg_DP_reg_28_ ( .D(n215), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[28]), .QN(n797) );
  SDFFR_X1 AReg_DP_reg_29_ ( .D(n214), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[29]) );
  SDFFR_X1 AReg_DP_reg_30_ ( .D(n212), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[30]), .QN(n772) );
  SDFFR_X1 RemSel_SP_reg ( .D(OpCode_SI[1]), .SI(1'b0), .SE(1'b0), .CK(n1094), 
        .RN(Rst_RBI), .Q(RemSel_SP), .QN(n3) );
  SDFFR_X1 CompInv_SP_reg ( .D(OpBSign_SI), .SI(1'b0), .SE(1'b0), .CK(n1094), 
        .RN(Rst_RBI), .Q(CompInv_SP), .QN(n823) );
  SDFFS_X1 AReg_DP_reg_12_ ( .D(n729), .SI(1'b0), .SE(1'b0), .CK(n1159), .SN(
        Rst_RBI), .Q(n757), .QN(AReg_DP[12]) );
  SNPS_CLOCK_GATE_HIGH_riscv_alu_div_0 clk_gate_ResReg_DP_reg_0_ ( .CLK(Clk_CI), .EN(n582), .ENCLK(n1159), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_alu_div_1 clk_gate_ResInv_SP_reg ( .CLK(Clk_CI), 
        .EN(n566), .ENCLK(n1094), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_alu_div_2 clk_gate_State_SP_reg_1_ ( .CLK(Clk_CI), 
        .EN(n1092), .ENCLK(n1090), .TE(1'b0) );
  SDFFR_X1 AReg_DP_reg_25_ ( .D(n218), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[25]), .QN(n803) );
  SDFFR_X1 AReg_DP_reg_26_ ( .D(n217), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[26]), .QN(n771) );
  SDFFR_X1 AReg_DP_reg_27_ ( .D(n216), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(AReg_DP[27]), .QN(n794) );
  SDFFR_X2 ResInv_SP_reg ( .D(n1093), .SI(1'b0), .SE(1'b0), .CK(n1094), .RN(
        Rst_RBI), .Q(ResInv_SP), .QN(n764) );
  BUF_X2 U6 ( .A(RemSel_SP), .Z(n1) );
  CLKBUF_X1 U11 ( .A(RemSel_SP), .Z(n7) );
  AND2_X2 U3 ( .A1(InVld_SI), .A2(n16), .ZN(n586) );
  BUF_X2 U4 ( .A(n19), .Z(n12) );
  BUF_X2 U7 ( .A(RemSel_SP), .Z(n2) );
  SDFFR_X1 BReg_DP_reg_24_ ( .D(n835), .SI(1'b0), .SE(1'b0), .CK(n1159), .RN(
        Rst_RBI), .Q(BReg_DP[24]), .QN(n812) );
  INV_X1 U5 ( .A(n580), .ZN(n817) );
  INV_X1 U8 ( .A(n580), .ZN(n821) );
  AND2_X1 U9 ( .A1(n661), .A2(n660), .ZN(n665) );
  AND2_X1 U12 ( .A1(n657), .A2(n656), .ZN(n661) );
  AND2_X1 U13 ( .A1(n645), .A2(n644), .ZN(n649) );
  AND2_X1 U14 ( .A1(n641), .A2(n640), .ZN(n645) );
  AND2_X1 U15 ( .A1(n629), .A2(n628), .ZN(n633) );
  NOR2_X1 U18 ( .A1(n26), .A2(n25), .ZN(n523) );
  AND2_X1 U19 ( .A1(n625), .A2(n624), .ZN(n629) );
  AND2_X1 U20 ( .A1(n613), .A2(n612), .ZN(n617) );
  AND2_X1 U22 ( .A1(n601), .A2(n600), .ZN(n613) );
  INV_X1 U26 ( .A(n570), .ZN(n820) );
  AND2_X1 U30 ( .A1(n677), .A2(n676), .ZN(n681) );
  AND2_X1 U43 ( .A1(n669), .A2(n668), .ZN(n673) );
  AND2_X1 U53 ( .A1(n693), .A2(n692), .ZN(n697) );
  AND2_X1 U272 ( .A1(n685), .A2(n684), .ZN(n689) );
  AOI21_X1 U275 ( .B1(n434), .B2(n432), .A(n355), .ZN(n826) );
  AOI21_X1 U276 ( .B1(n412), .B2(n410), .A(n369), .ZN(n827) );
  AOI21_X1 U499 ( .B1(n481), .B2(n52), .A(n51), .ZN(n828) );
  INV_X1 U500 ( .A(n586), .ZN(n829) );
  INV_X1 U501 ( .A(n586), .ZN(n830) );
  INV_X1 U506 ( .A(n3), .ZN(n5) );
  MUX2_X1 U507 ( .A(AReg_DP[0]), .B(ResReg_DP_rev[0]), .S(n3), .Z(Res_DO[0])
         );
  XOR2_X1 U508 ( .A(n641), .B(n640), .Z(n639) );
  XOR2_X1 U509 ( .A(n657), .B(n656), .Z(n655) );
  XOR2_X1 U510 ( .A(n625), .B(n624), .Z(n623) );
  XOR2_X1 U511 ( .A(n601), .B(n600), .Z(n597) );
  XOR2_X1 U512 ( .A(n693), .B(n692), .Z(n691) );
  XOR2_X1 U513 ( .A(n685), .B(n684), .Z(n683) );
  XOR2_X1 U514 ( .A(n677), .B(n676), .Z(n675) );
  XOR2_X1 U515 ( .A(n669), .B(n668), .Z(n667) );
  NAND2_X1 U853 ( .A1(Cnt_DP[0]), .A2(State_SP[0]), .ZN(n1092) );
  NOR2_X1 U854 ( .A1(n587), .A2(n588), .ZN(n1093) );
  OAI21_X1 U855 ( .B1(n823), .B2(n821), .A(n1042), .ZN(n1096) );
  NAND2_X1 U856 ( .A1(OpB_DI[31]), .A2(n566), .ZN(n1042) );
  OAI21_X1 U857 ( .B1(n790), .B2(n821), .A(n1043), .ZN(n1097) );
  NAND2_X1 U858 ( .A1(OpB_DI[30]), .A2(n566), .ZN(n1043) );
  OAI21_X1 U859 ( .B1(n810), .B2(n817), .A(n1044), .ZN(n1098) );
  NAND2_X1 U860 ( .A1(OpB_DI[29]), .A2(n566), .ZN(n1044) );
  OAI22_X1 U861 ( .A1(n1089), .A2(n773), .B1(n829), .B2(n1045), .ZN(n1099) );
  INV_X1 U862 ( .A(OpB_DI[28]), .ZN(n1045) );
  OAI22_X1 U863 ( .A1(n821), .A2(n809), .B1(n829), .B2(n1046), .ZN(n1100) );
  INV_X1 U864 ( .A(OpB_DI[27]), .ZN(n1046) );
  OAI22_X1 U865 ( .A1(n1087), .A2(n800), .B1(n830), .B2(n1047), .ZN(n1101) );
  INV_X1 U866 ( .A(OpB_DI[26]), .ZN(n1047) );
  OAI22_X1 U867 ( .A1(n821), .A2(n825), .B1(n829), .B2(n1048), .ZN(n1102) );
  INV_X1 U868 ( .A(OpB_DI[25]), .ZN(n1048) );
  OAI21_X1 U869 ( .B1(n808), .B2(n1089), .A(n1049), .ZN(n835) );
  NAND2_X1 U870 ( .A1(OpB_DI[24]), .A2(n566), .ZN(n1049) );
  OAI21_X1 U871 ( .B1(n1050), .B2(n829), .A(n1051), .ZN(n1103) );
  NAND2_X1 U872 ( .A1(n580), .A2(BReg_DP[24]), .ZN(n1051) );
  INV_X1 U873 ( .A(OpB_DI[23]), .ZN(n1050) );
  OAI21_X1 U874 ( .B1(n1052), .B2(n829), .A(n1053), .ZN(n1104) );
  NAND2_X1 U875 ( .A1(n580), .A2(BReg_DP[23]), .ZN(n1053) );
  INV_X1 U876 ( .A(OpB_DI[22]), .ZN(n1052) );
  OAI21_X1 U877 ( .B1(n1054), .B2(n830), .A(n1055), .ZN(n1105) );
  NAND2_X1 U878 ( .A1(n580), .A2(BReg_DP[22]), .ZN(n1055) );
  INV_X1 U879 ( .A(OpB_DI[21]), .ZN(n1054) );
  OAI21_X1 U880 ( .B1(n1056), .B2(n829), .A(n1057), .ZN(n1106) );
  NAND2_X1 U881 ( .A1(n580), .A2(BReg_DP[21]), .ZN(n1057) );
  INV_X1 U882 ( .A(OpB_DI[20]), .ZN(n1056) );
  OAI21_X1 U883 ( .B1(n1058), .B2(n829), .A(n1059), .ZN(n1107) );
  NAND2_X1 U884 ( .A1(n580), .A2(BReg_DP[20]), .ZN(n1059) );
  INV_X1 U885 ( .A(OpB_DI[19]), .ZN(n1058) );
  OAI22_X1 U886 ( .A1(n1087), .A2(n815), .B1(n829), .B2(n1060), .ZN(n1108) );
  INV_X1 U887 ( .A(OpB_DI[18]), .ZN(n1060) );
  OAI21_X1 U888 ( .B1(n1061), .B2(n830), .A(n1062), .ZN(n1109) );
  NAND2_X1 U889 ( .A1(n580), .A2(BReg_DP[18]), .ZN(n1062) );
  INV_X1 U890 ( .A(OpB_DI[17]), .ZN(n1061) );
  OAI21_X1 U891 ( .B1(n1063), .B2(n829), .A(n1064), .ZN(n1110) );
  NAND2_X1 U892 ( .A1(n580), .A2(BReg_DP[17]), .ZN(n1064) );
  INV_X1 U893 ( .A(OpB_DI[16]), .ZN(n1063) );
  OAI21_X1 U894 ( .B1(n1065), .B2(n829), .A(n1066), .ZN(n1111) );
  NAND2_X1 U895 ( .A1(n580), .A2(BReg_DP[16]), .ZN(n1066) );
  INV_X1 U896 ( .A(OpB_DI[15]), .ZN(n1065) );
  OAI21_X1 U897 ( .B1(n1067), .B2(n830), .A(n1068), .ZN(n1112) );
  NAND2_X1 U898 ( .A1(n580), .A2(BReg_DP[15]), .ZN(n1068) );
  INV_X1 U899 ( .A(OpB_DI[14]), .ZN(n1067) );
  OAI21_X1 U900 ( .B1(n1069), .B2(n829), .A(n1070), .ZN(n1113) );
  NAND2_X1 U901 ( .A1(n580), .A2(BReg_DP[14]), .ZN(n1070) );
  INV_X1 U902 ( .A(OpB_DI[13]), .ZN(n1069) );
  AOI221_X1 U903 ( .B1(State_SP[0]), .B2(n1071), .C1(n1072), .C2(n1071), .A(
        State_SP[1]), .ZN(n1114) );
  NAND2_X1 U904 ( .A1(InVld_SI), .A2(OpB_DI[12]), .ZN(n1072) );
  NAND2_X1 U905 ( .A1(BReg_DP[13]), .A2(State_SP[0]), .ZN(n1071) );
  OAI21_X1 U906 ( .B1(n759), .B2(n1088), .A(n1073), .ZN(n1115) );
  NAND2_X1 U907 ( .A1(OpB_DI[11]), .A2(n586), .ZN(n1073) );
  OAI22_X1 U908 ( .A1(n1088), .A2(n758), .B1(n830), .B2(n1074), .ZN(n1116) );
  INV_X1 U909 ( .A(OpB_DI[10]), .ZN(n1074) );
  OAI22_X1 U910 ( .A1(n817), .A2(n769), .B1(n829), .B2(n1075), .ZN(n1117) );
  INV_X1 U911 ( .A(OpB_DI[9]), .ZN(n1075) );
  OAI22_X1 U912 ( .A1(n1088), .A2(n733), .B1(n829), .B2(n1076), .ZN(n1118) );
  INV_X1 U913 ( .A(OpB_DI[8]), .ZN(n1076) );
  OAI22_X1 U914 ( .A1(n1089), .A2(n761), .B1(n830), .B2(n1077), .ZN(n1119) );
  INV_X1 U915 ( .A(OpB_DI[7]), .ZN(n1077) );
  OAI21_X1 U916 ( .B1(n824), .B2(n817), .A(n1078), .ZN(n1120) );
  NAND2_X1 U917 ( .A1(OpB_DI[6]), .A2(n566), .ZN(n1078) );
  OAI22_X1 U918 ( .A1(n817), .A2(n750), .B1(n829), .B2(n1079), .ZN(n1121) );
  INV_X1 U919 ( .A(OpB_DI[5]), .ZN(n1079) );
  OAI21_X1 U920 ( .B1(n768), .B2(n1087), .A(n1080), .ZN(n1122) );
  NAND2_X1 U921 ( .A1(OpB_DI[4]), .A2(n566), .ZN(n1080) );
  OAI22_X1 U922 ( .A1(n1089), .A2(n749), .B1(n829), .B2(n1081), .ZN(n1123) );
  INV_X1 U923 ( .A(OpB_DI[3]), .ZN(n1081) );
  OAI22_X1 U924 ( .A1(n1087), .A2(n766), .B1(n830), .B2(n1082), .ZN(n1124) );
  INV_X1 U925 ( .A(OpB_DI[2]), .ZN(n1082) );
  OAI22_X1 U926 ( .A1(n1088), .A2(n767), .B1(n830), .B2(n1083), .ZN(n1125) );
  INV_X1 U927 ( .A(OpB_DI[1]), .ZN(n1083) );
  INV_X1 U928 ( .A(n1084), .ZN(n1126) );
  AOI22_X1 U929 ( .A1(n580), .A2(BReg_DP[1]), .B1(OpB_DI[0]), .B2(n566), .ZN(
        n1084) );
  NOR2_X1 U930 ( .A1(n817), .A2(n1085), .ZN(n1127) );
  NAND2_X1 U931 ( .A1(n203), .A2(n204), .ZN(n1085) );
  NOR2_X1 U932 ( .A1(n788), .A2(n817), .ZN(n1128) );
  NOR2_X1 U933 ( .A1(n731), .A2(n1089), .ZN(n1129) );
  NOR2_X1 U934 ( .A1(n730), .A2(n821), .ZN(n1130) );
  NOR2_X1 U935 ( .A1(n774), .A2(n1088), .ZN(n1131) );
  NOR2_X1 U936 ( .A1(n734), .A2(n820), .ZN(n1132) );
  NOR2_X1 U937 ( .A1(n775), .A2(n1087), .ZN(n1133) );
  NOR2_X1 U938 ( .A1(n735), .A2(n817), .ZN(n1134) );
  NOR2_X1 U939 ( .A1(n776), .A2(n817), .ZN(n1135) );
  NOR2_X1 U940 ( .A1(n736), .A2(n821), .ZN(n1136) );
  NOR2_X1 U941 ( .A1(n777), .A2(n821), .ZN(n1137) );
  NOR2_X1 U942 ( .A1(n737), .A2(n820), .ZN(n1138) );
  NOR2_X1 U943 ( .A1(n778), .A2(n821), .ZN(n1139) );
  NOR2_X1 U944 ( .A1(n738), .A2(n821), .ZN(n1140) );
  NOR2_X1 U945 ( .A1(n779), .A2(n817), .ZN(n1141) );
  NOR2_X1 U946 ( .A1(n739), .A2(n817), .ZN(n1142) );
  NOR2_X1 U947 ( .A1(n780), .A2(n1089), .ZN(n1143) );
  NOR2_X1 U948 ( .A1(n740), .A2(n817), .ZN(n1144) );
  NOR2_X1 U949 ( .A1(n781), .A2(n817), .ZN(n1145) );
  NOR2_X1 U950 ( .A1(n741), .A2(n821), .ZN(n1146) );
  NOR2_X1 U951 ( .A1(n782), .A2(n1088), .ZN(n1147) );
  NOR2_X1 U952 ( .A1(n742), .A2(n1086), .ZN(n1148) );
  INV_X1 U953 ( .A(n580), .ZN(n1086) );
  NOR2_X1 U954 ( .A1(n783), .A2(n1087), .ZN(n1149) );
  NOR2_X1 U955 ( .A1(n743), .A2(n1087), .ZN(n1150) );
  INV_X1 U956 ( .A(n580), .ZN(n1087) );
  NOR2_X1 U957 ( .A1(n784), .A2(n817), .ZN(n1151) );
  NOR2_X1 U958 ( .A1(n744), .A2(n1088), .ZN(n1152) );
  INV_X1 U959 ( .A(n580), .ZN(n1088) );
  NOR2_X1 U960 ( .A1(n785), .A2(n821), .ZN(n1153) );
  NOR2_X1 U961 ( .A1(n745), .A2(n1089), .ZN(n1154) );
  INV_X1 U962 ( .A(n580), .ZN(n1089) );
  NOR2_X1 U963 ( .A1(n786), .A2(n821), .ZN(n1155) );
  NOR2_X1 U964 ( .A1(n746), .A2(n820), .ZN(n1156) );
  NOR2_X1 U965 ( .A1(n787), .A2(n817), .ZN(n1157) );
  NOR2_X1 U966 ( .A1(n747), .A2(n821), .ZN(n1158) );
endmodule


module alu_ff ( in_i, first_one_o, no_ones_o );
  input [31:0] in_i;
  output [4:0] first_one_o;
  output no_ones_o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n55, n56, n57, n58, n59,
         n60, n61, n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;

  OR2_X1 U1 ( .A1(in_i[16]), .A2(in_i[17]), .ZN(n35) );
  MUX2_X1 U3 ( .A(n43), .B(n42), .S(n74), .Z(first_one_o[1]) );
  CLKBUF_X1 U4 ( .A(n74), .Z(first_one_o[4]) );
  NOR2_X1 U7 ( .A1(n32), .A2(in_i[24]), .ZN(n23) );
  NAND3_X1 U8 ( .A1(n30), .A2(n29), .A3(n1), .ZN(n43) );
  OR2_X1 U9 ( .A1(n25), .A2(n31), .ZN(n1) );
  AND2_X1 U10 ( .A1(n37), .A2(n5), .ZN(n3) );
  INV_X1 U11 ( .A(n20), .ZN(n5) );
  NOR2_X1 U12 ( .A1(n33), .A2(in_i[24]), .ZN(n6) );
  AND3_X1 U13 ( .A1(n23), .A2(n44), .A3(n9), .ZN(n73) );
  INV_X1 U14 ( .A(in_i[28]), .ZN(n9) );
  NOR2_X1 U15 ( .A1(n44), .A2(n8), .ZN(n7) );
  AND2_X1 U16 ( .A1(n23), .A2(n44), .ZN(n4) );
  INV_X1 U17 ( .A(n34), .ZN(n8) );
  NOR2_X1 U18 ( .A1(n3), .A2(n36), .ZN(n38) );
  NOR2_X1 U19 ( .A1(n15), .A2(n11), .ZN(n10) );
  NOR2_X1 U20 ( .A1(n46), .A2(n74), .ZN(n83) );
  NOR2_X1 U21 ( .A1(in_i[14]), .A2(in_i[15]), .ZN(n2) );
  AND3_X1 U22 ( .A1(n74), .A2(n73), .A3(n24), .ZN(no_ones_o) );
  NAND2_X1 U23 ( .A1(n40), .A2(n41), .ZN(n42) );
  NOR2_X1 U25 ( .A1(n7), .A2(n4), .ZN(n47) );
  NAND2_X1 U26 ( .A1(n25), .A2(n14), .ZN(n27) );
  NAND2_X1 U28 ( .A1(n44), .A2(n6), .ZN(n70) );
  INV_X1 U29 ( .A(n27), .ZN(n12) );
  NAND3_X1 U30 ( .A1(n12), .A2(n10), .A3(n79), .ZN(n29) );
  AND4_X2 U31 ( .A1(n12), .A2(n10), .A3(n79), .A4(n2), .ZN(n74) );
  NAND2_X1 U32 ( .A1(n17), .A2(n78), .ZN(n11) );
  OR2_X1 U33 ( .A1(in_i[1]), .A2(in_i[0]), .ZN(n31) );
  OR2_X1 U34 ( .A1(in_i[2]), .A2(in_i[3]), .ZN(n13) );
  NOR2_X1 U35 ( .A1(in_i[5]), .A2(in_i[4]), .ZN(n14) );
  OR2_X1 U36 ( .A1(in_i[6]), .A2(in_i[7]), .ZN(n15) );
  OR2_X1 U37 ( .A1(in_i[9]), .A2(in_i[8]), .ZN(n26) );
  OR2_X1 U38 ( .A1(in_i[10]), .A2(in_i[11]), .ZN(n16) );
  NOR2_X2 U39 ( .A1(n26), .A2(n16), .ZN(n79) );
  INV_X1 U40 ( .A(in_i[13]), .ZN(n78) );
  INV_X1 U41 ( .A(in_i[12]), .ZN(n17) );
  OR2_X1 U42 ( .A1(in_i[18]), .A2(in_i[19]), .ZN(n18) );
  NOR2_X1 U44 ( .A1(in_i[20]), .A2(in_i[21]), .ZN(n19) );
  AND2_X1 U45 ( .A1(n34), .A2(n19), .ZN(n37) );
  NOR2_X1 U46 ( .A1(in_i[22]), .A2(in_i[23]), .ZN(n20) );
  NOR2_X1 U47 ( .A1(in_i[26]), .A2(in_i[27]), .ZN(n22) );
  INV_X1 U48 ( .A(in_i[25]), .ZN(n21) );
  NAND2_X1 U49 ( .A1(n22), .A2(n21), .ZN(n32) );
  NOR3_X1 U50 ( .A1(in_i[29]), .A2(in_i[30]), .A3(in_i[31]), .ZN(n24) );
  OAI21_X1 U51 ( .B1(n79), .B2(n26), .A(n56), .ZN(n28) );
  NAND2_X1 U52 ( .A1(n28), .A2(n12), .ZN(n30) );
  INV_X1 U53 ( .A(in_i[29]), .ZN(n60) );
  NAND2_X1 U54 ( .A1(n73), .A2(n60), .ZN(n41) );
  INV_X1 U55 ( .A(n32), .ZN(n33) );
  NOR2_X1 U56 ( .A1(n34), .A2(n35), .ZN(n36) );
  OAI21_X1 U57 ( .B1(n70), .B2(in_i[25]), .A(n38), .ZN(n39) );
  INV_X1 U58 ( .A(n39), .ZN(n40) );
  INV_X1 U59 ( .A(n56), .ZN(n46) );
  AND2_X1 U60 ( .A1(n44), .A2(first_one_o[4]), .ZN(n45) );
  OR2_X1 U61 ( .A1(n83), .A2(n45), .ZN(first_one_o[3]) );
  INV_X1 U62 ( .A(n83), .ZN(n51) );
  INV_X1 U63 ( .A(n79), .ZN(n50) );
  NAND2_X1 U64 ( .A1(n46), .A2(n25), .ZN(n48) );
  MUX2_X1 U65 ( .A(n48), .B(n47), .S(n74), .Z(n49) );
  OAI21_X1 U66 ( .B1(n51), .B2(n50), .A(n49), .ZN(first_one_o[2]) );
  INV_X1 U67 ( .A(in_i[6]), .ZN(n53) );
  INV_X1 U68 ( .A(in_i[4]), .ZN(n52) );
  OAI21_X1 U69 ( .B1(n53), .B2(in_i[5]), .A(n52), .ZN(n55) );
  OAI21_X1 U70 ( .B1(n56), .B2(n55), .A(n25), .ZN(n59) );
  INV_X1 U71 ( .A(in_i[1]), .ZN(n57) );
  AOI21_X1 U72 ( .B1(n57), .B2(in_i[2]), .A(in_i[0]), .ZN(n58) );
  NAND2_X1 U73 ( .A1(n59), .A2(n58), .ZN(n76) );
  NAND2_X1 U74 ( .A1(n60), .A2(in_i[30]), .ZN(n72) );
  INV_X1 U75 ( .A(in_i[26]), .ZN(n61) );
  NOR2_X1 U76 ( .A1(n61), .A2(in_i[25]), .ZN(n69) );
  INV_X1 U77 ( .A(in_i[22]), .ZN(n62) );
  AOI21_X1 U78 ( .B1(n62), .B2(in_i[23]), .A(in_i[21]), .ZN(n64) );
  OAI21_X1 U79 ( .B1(in_i[20]), .B2(n64), .A(n34), .ZN(n67) );
  INV_X1 U80 ( .A(in_i[17]), .ZN(n65) );
  AOI21_X1 U81 ( .B1(n65), .B2(in_i[18]), .A(in_i[16]), .ZN(n66) );
  NAND2_X1 U82 ( .A1(n67), .A2(n66), .ZN(n68) );
  OAI21_X1 U83 ( .B1(n70), .B2(n69), .A(n68), .ZN(n71) );
  AOI21_X1 U84 ( .B1(n73), .B2(n72), .A(n71), .ZN(n75) );
  MUX2_X1 U85 ( .A(n76), .B(n75), .S(n74), .Z(n85) );
  INV_X1 U86 ( .A(in_i[9]), .ZN(n77) );
  AOI21_X1 U87 ( .B1(n77), .B2(in_i[10]), .A(in_i[8]), .ZN(n81) );
  AOI21_X1 U88 ( .B1(n78), .B2(in_i[14]), .A(in_i[12]), .ZN(n80) );
  MUX2_X1 U89 ( .A(n81), .B(n80), .S(n79), .Z(n82) );
  NAND2_X1 U90 ( .A1(n83), .A2(n82), .ZN(n84) );
  NAND2_X1 U91 ( .A1(n85), .A2(n84), .ZN(first_one_o[0]) );
  AND2_X1 U27 ( .A1(n37), .A2(n20), .ZN(n44) );
  NOR2_X1 U2 ( .A1(n27), .A2(n15), .ZN(n56) );
  NOR2_X2 U43 ( .A1(n35), .A2(n18), .ZN(n34) );
  NOR2_X2 U5 ( .A1(n13), .A2(n31), .ZN(n25) );
endmodule


module alu_popcnt ( in_i, result_o );
  input [31:0] in_i;
  output [5:0] result_o;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;

  FA_X1 U1 ( .A(in_i[6]), .B(in_i[2]), .CI(in_i[4]), .CO(n10), .S(n32) );
  FA_X1 U2 ( .A(in_i[22]), .B(in_i[20]), .CI(in_i[18]), .CO(n8), .S(n31) );
  FA_X1 U3 ( .A(in_i[16]), .B(in_i[14]), .CI(in_i[12]), .CO(n9), .S(n21) );
  FA_X1 U4 ( .A(in_i[10]), .B(in_i[0]), .CI(in_i[8]), .CO(n12), .S(n23) );
  HA_X1 U5 ( .A(in_i[5]), .B(in_i[3]), .CO(n11), .S(n22) );
  FA_X1 U6 ( .A(in_i[28]), .B(in_i[26]), .CI(in_i[24]), .CO(n5), .S(n30) );
  FA_X1 U7 ( .A(n4), .B(n3), .CI(n2), .CO(n15), .S(n36) );
  FA_X1 U8 ( .A(n7), .B(n6), .CI(n5), .CO(n14), .S(n24) );
  FA_X1 U9 ( .A(n10), .B(n9), .CI(n8), .CO(n17), .S(n37) );
  HA_X1 U10 ( .A(n12), .B(n11), .CO(n16), .S(n25) );
  FA_X1 U11 ( .A(n15), .B(n14), .CI(n13), .CO(n43), .S(n18) );
  HA_X1 U12 ( .A(n17), .B(n16), .CO(n42), .S(n13) );
  FA_X1 U13 ( .A(n20), .B(n19), .CI(n18), .CO(n48), .S(n51) );
  FA_X1 U14 ( .A(in_i[11]), .B(in_i[13]), .CI(in_i[15]), .CO(n3), .S(n35) );
  FA_X1 U15 ( .A(in_i[1]), .B(in_i[7]), .CI(in_i[9]), .CO(n7), .S(n34) );
  FA_X1 U16 ( .A(n23), .B(n22), .CI(n21), .CO(n26), .S(n33) );
  FA_X1 U17 ( .A(in_i[29]), .B(in_i[31]), .CI(in_i[30]), .CO(n4), .S(n29) );
  FA_X1 U18 ( .A(in_i[23]), .B(in_i[25]), .CI(in_i[27]), .CO(n6), .S(n28) );
  FA_X1 U19 ( .A(in_i[17]), .B(in_i[21]), .CI(in_i[19]), .CO(n2), .S(n27) );
  FA_X1 U20 ( .A(n26), .B(n25), .CI(n24), .CO(n19), .S(n39) );
  FA_X1 U21 ( .A(n29), .B(n28), .CI(n27), .CO(n40), .S(n57) );
  FA_X1 U22 ( .A(n32), .B(n31), .CI(n30), .CO(n38), .S(n56) );
  FA_X1 U23 ( .A(n35), .B(n34), .CI(n33), .CO(n41), .S(n55) );
  FA_X1 U24 ( .A(n38), .B(n37), .CI(n36), .CO(n20), .S(n53) );
  FA_X1 U25 ( .A(n41), .B(n40), .CI(n39), .CO(n50), .S(n52) );
  HA_X1 U26 ( .A(n43), .B(n42), .CO(n44), .S(n47) );
  HA_X1 U27 ( .A(n45), .B(n44), .CO(result_o[5]), .S(result_o[4]) );
  FA_X1 U28 ( .A(n48), .B(n47), .CI(n46), .CO(n45), .S(result_o[3]) );
  FA_X1 U29 ( .A(n51), .B(n50), .CI(n49), .CO(n46), .S(result_o[2]) );
  FA_X1 U30 ( .A(n54), .B(n53), .CI(n52), .CO(n49), .S(result_o[1]) );
  FA_X1 U31 ( .A(n57), .B(n56), .CI(n55), .CO(n54), .S(result_o[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_hwloop_regs_N_REGS2_4 ( CLK, EN, ENCLK, TE
 );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_hwloop_regs_N_REGS2_3 ( CLK, EN, ENCLK, TE
 );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_hwloop_regs_N_REGS2_2 ( CLK, EN, ENCLK, TE
 );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_hwloop_regs_N_REGS2_1 ( CLK, EN, ENCLK, TE
 );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_hwloop_regs_N_REGS2_0 ( CLK, EN, ENCLK, TE
 );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_int_controller_PULP_SECURE1_0 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net8, net11;
  assign net8 = EN;
  assign net11 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net8), .SE(net11), .GCK(ENCLK) );
endmodule


module riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0 ( clk, rst_n, 
        test_en_i, raddr_a_i, rdata_a_o, raddr_b_i, rdata_b_o, raddr_c_i, 
        rdata_c_o, waddr_a_i, wdata_a_i, we_a_i, waddr_b_i, wdata_b_i, we_b_i
 );
  input [5:0] raddr_a_i;
  output [31:0] rdata_a_o;
  input [5:0] raddr_b_i;
  output [31:0] rdata_b_o;
  input [5:0] raddr_c_i;
  output [31:0] rdata_c_o;
  input [5:0] waddr_a_i;
  input [31:0] wdata_a_i;
  input [5:0] waddr_b_i;
  input [31:0] wdata_b_i;
  input clk, rst_n, test_en_i, we_a_i, we_b_i;
  wire   n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1031, n1033, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1539, n1541, n1543,
         n1545, n1546, n1548, n1550, n1551, n1554, n1555, n1556, n1559, n1560,
         n1561, n1563, n1565, n1566, n1568, n1570, n1571, n1575, n1576, n1577,
         n1579, n1581, n1582, n1585, n1586, n1587, n1591, n1592, n1593, n1596,
         n1597, n1598, n1601, n1602, n1603, n1604, n1606, n1608, n1609, n1610,
         n1611, n1614, n1615, n1616, n1617, n1618, n1620, n1621, n1622, n1623,
         n1624, n1625, n1627, n1629, n1631, n1632, n1634, n1636, n1637, n1638,
         n1639, n1640, n1641, n1643, n1644, n1645, n1646, n1647, n1648, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1688, n1689, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2259, n2260,
         n2261, n2262, n2263, n2264, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2468, n2469, n2473, n2474, n2478,
         n2479, n2480, n2481, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2530, n2532, n2533,
         n2534, n2535, n2539, n2540, n2541, n2542, n2546, n2547, n2548, n2549,
         n2550, n2551, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3768, n3769, n3770, n3771, n3772, n3774, n3845, n3846, n3847, n3848,
         n3849, n3851, n4002, n4004, n4011, n4017, n4037, n4040, n4043, n4047,
         n4374, n4380, n4382, n4385, n4386, n4394, n4408, n4410, n4412, n4414,
         n4416, n4418, n4420, n4422, n4424, n4426, n4430, n4432, n4434, n4436,
         n4439, n4441, n4444, n4447, n4449, n4452, n4458, n4459, n4461, n4467,
         n4468, n4470, n4472, n4474, n4477, n4486, n4614, n4618, n4623, n4729,
         n4730, n4731, n4732, n4734, n4736, n4737, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9198;
  wire   [991:0] mem;

  OR2_X1 U11 ( .A1(n1344), .A2(raddr_c_i[1]), .ZN(n1362) );
  OR2_X1 U12 ( .A1(raddr_c_i[1]), .A2(raddr_c_i[0]), .ZN(n1358) );
  BUF_X1 U15 ( .A(n3092), .Z(n3066) );
  BUF_X1 U47 ( .A(raddr_a_i[2]), .Z(n997) );
  OR2_X2 U49 ( .A1(n1720), .A2(n1719), .ZN(n1723) );
  NOR2_X1 U50 ( .A1(n3415), .A2(n993), .ZN(n3416) );
  NAND4_X1 U51 ( .A1(n3410), .A2(n3411), .A3(n3412), .A4(n3413), .ZN(n993) );
  BUF_X2 U54 ( .A(n3131), .Z(n3351) );
  BUF_X2 U57 ( .A(n3207), .Z(n994) );
  BUF_X2 U58 ( .A(n3207), .Z(n995) );
  BUF_X2 U61 ( .A(n2162), .Z(n3350) );
  NAND4_X1 U70 ( .A1(n998), .A2(n999), .A3(n1000), .A4(n1001), .ZN(
        rdata_a_o[5]) );
  AND4_X1 U71 ( .A1(n2152), .A2(n2151), .A3(n2150), .A4(n2149), .ZN(n998) );
  AND4_X1 U72 ( .A1(n2160), .A2(n2159), .A3(n2158), .A4(n2157), .ZN(n999) );
  AND4_X1 U73 ( .A1(n2168), .A2(n2167), .A3(n2166), .A4(n2165), .ZN(n1000) );
  AND4_X1 U74 ( .A1(n2174), .A2(n2173), .A3(n2172), .A4(n2171), .ZN(n1001) );
  BUF_X2 U75 ( .A(n3040), .Z(n3592) );
  BUF_X1 U81 ( .A(n2170), .Z(n3269) );
  BUF_X2 U83 ( .A(n3176), .Z(n1083) );
  AND2_X1 U87 ( .A1(n3206), .A2(n3205), .ZN(n1002) );
  AND2_X1 U88 ( .A1(n2892), .A2(n2894), .ZN(n1003) );
  AND4_X1 U89 ( .A1(n2902), .A2(n2901), .A3(n2900), .A4(n2899), .ZN(n1004) );
  BUF_X2 U96 ( .A(n2147), .Z(n1011) );
  BUF_X2 U97 ( .A(n2147), .Z(n1012) );
  BUF_X2 U98 ( .A(n2147), .Z(n1013) );
  BUF_X2 U103 ( .A(n2156), .Z(n1017) );
  BUF_X2 U106 ( .A(n3102), .Z(n1020) );
  BUF_X2 U107 ( .A(n3102), .Z(n1021) );
  BUF_X2 U108 ( .A(n3102), .Z(n1022) );
  BUF_X2 U109 ( .A(n2161), .Z(n1023) );
  BUF_X2 U110 ( .A(n2161), .Z(n1024) );
  AND2_X1 U111 ( .A1(n1704), .A2(n1710), .ZN(n2161) );
  BUF_X1 U116 ( .A(n2155), .Z(n1028) );
  BUF_X2 U117 ( .A(n2155), .Z(n1029) );
  BUF_X1 U119 ( .A(n1028), .Z(n1031) );
  AND2_X1 U121 ( .A1(n1698), .A2(n1710), .ZN(n2155) );
  BUF_X1 U147 ( .A(n1414), .Z(n3001) );
  BUF_X1 U152 ( .A(n2164), .Z(n1067) );
  BUF_X1 U153 ( .A(n2164), .Z(n1092) );
  BUF_X1 U154 ( .A(n2164), .Z(n1093) );
  AND2_X1 U155 ( .A1(n1718), .A2(n1710), .ZN(n2164) );
  INV_X1 U158 ( .A(wdata_b_i[12]), .ZN(n4432) );
  CLKBUF_X1 U163 ( .A(wdata_a_i[27]), .Z(n4394) );
  CLKBUF_X1 U165 ( .A(wdata_a_i[29]), .Z(n4468) );
  CLKBUF_X1 U166 ( .A(wdata_a_i[30]), .Z(n4472) );
  CLKBUF_X1 U167 ( .A(wdata_a_i[30]), .Z(n4623) );
  CLKBUF_X1 U169 ( .A(wdata_a_i[28]), .Z(n4618) );
  CLKBUF_X1 U170 ( .A(wdata_a_i[31]), .Z(n4477) );
  CLKBUF_X1 U171 ( .A(wdata_a_i[25]), .Z(n4614) );
  CLKBUF_X1 U172 ( .A(wdata_a_i[24]), .Z(n4386) );
  CLKBUF_X1 U174 ( .A(wdata_a_i[26]), .Z(n4459) );
  NAND4_X1 U177 ( .A1(n1076), .A2(n1003), .A3(n1074), .A4(n1004), .ZN(
        rdata_a_o[3]) );
  NOR2_X1 U178 ( .A1(n3215), .A2(n3216), .ZN(n1079) );
  AND4_X1 U179 ( .A1(n2898), .A2(n2897), .A3(n2896), .A4(n2895), .ZN(n1076) );
  CLKBUF_X2 U201 ( .A(n3061), .Z(n3358) );
  BUF_X1 U206 ( .A(n3222), .Z(n1089) );
  BUF_X1 U208 ( .A(n3222), .Z(n1091) );
  BUF_X2 U210 ( .A(n3196), .Z(n1069) );
  BUF_X1 U211 ( .A(n3222), .Z(n1090) );
  BUF_X2 U214 ( .A(n3114), .Z(n1072) );
  BUF_X2 U218 ( .A(n2169), .Z(n1073) );
  AND2_X2 U219 ( .A1(n1691), .A2(n1717), .ZN(n3131) );
  NOR2_X1 U220 ( .A1(n2907), .A2(n1075), .ZN(n1074) );
  NAND2_X1 U221 ( .A1(n2891), .A2(n2893), .ZN(n1075) );
  NOR3_X1 U222 ( .A1(n3450), .A2(n1078), .A3(n1077), .ZN(n3463) );
  NAND2_X1 U223 ( .A1(n3443), .A2(n3442), .ZN(n1077) );
  NAND2_X1 U224 ( .A1(n3445), .A2(n3444), .ZN(n1078) );
  NAND3_X1 U226 ( .A1(n3229), .A2(n1079), .A3(n1002), .ZN(rdata_a_o[11]) );
  NAND2_X1 U227 ( .A1(n3076), .A2(n3077), .ZN(n3087) );
  NOR2_X1 U228 ( .A1(n1696), .A2(n1719), .ZN(n1706) );
  NOR2_X1 U232 ( .A1(n4773), .A2(raddr_a_i[0]), .ZN(n1708) );
  INV_X1 U233 ( .A(waddr_b_i[4]), .ZN(n3768) );
  INV_X1 U234 ( .A(waddr_a_i[1]), .ZN(n2527) );
  OR2_X1 U235 ( .A1(waddr_a_i[3]), .A2(waddr_a_i[4]), .ZN(n2525) );
  OR2_X1 U236 ( .A1(n1535), .A2(waddr_a_i[0]), .ZN(n2532) );
  INV_X1 U237 ( .A(waddr_a_i[2]), .ZN(n2533) );
  AND4_X1 U300 ( .A1(n3158), .A2(n3157), .A3(n3156), .A4(n3155), .ZN(n1094) );
  OR2_X1 U301 ( .A1(n4773), .A2(raddr_a_i[0]), .ZN(n1095) );
  NAND2_X1 U302 ( .A1(n1096), .A2(n3099), .ZN(rdata_a_o[6]) );
  NOR2_X1 U303 ( .A1(n3098), .A2(n3097), .ZN(n1096) );
  BUF_X2 U304 ( .A(n3061), .Z(n3587) );
  NAND3_X1 U305 ( .A1(n3175), .A2(n1097), .A3(n1094), .ZN(rdata_a_o[9]) );
  NOR2_X1 U306 ( .A1(n3160), .A2(n3159), .ZN(n1097) );
  INV_X1 U315 ( .A(we_a_i), .ZN(n1535) );
  NAND2_X1 U316 ( .A1(waddr_a_i[0]), .A2(we_a_i), .ZN(n1586) );
  NOR2_X1 U317 ( .A1(n1622), .A2(n2533), .ZN(n1637) );
  OR2_X1 U318 ( .A1(waddr_a_i[1]), .A2(n1586), .ZN(n2480) );
  AND2_X1 U319 ( .A1(waddr_b_i[1]), .A2(waddr_b_i[3]), .ZN(n3770) );
  NAND3_X1 U320 ( .A1(n2468), .A2(waddr_b_i[1]), .A3(waddr_b_i[4]), .ZN(n1608)
         );
  NAND2_X1 U321 ( .A1(n2478), .A2(waddr_b_i[4]), .ZN(n1591) );
  NAND2_X1 U322 ( .A1(n3845), .A2(n3768), .ZN(n1601) );
  OR2_X1 U323 ( .A1(n1614), .A2(n1559), .ZN(n2540) );
  OR2_X1 U324 ( .A1(n1560), .A2(waddr_b_i[2]), .ZN(n3769) );
  INV_X1 U325 ( .A(wdata_b_i[13]), .ZN(n4434) );
  INV_X1 U327 ( .A(wdata_b_i[29]), .ZN(n4467) );
  INV_X1 U329 ( .A(raddr_b_i[0]), .ZN(n1098) );
  NAND2_X1 U330 ( .A1(raddr_b_i[1]), .A2(n1098), .ZN(n1121) );
  NAND3_X1 U331 ( .A1(raddr_b_i[4]), .A2(raddr_b_i[2]), .A3(raddr_b_i[3]), 
        .ZN(n1104) );
  NOR2_X1 U332 ( .A1(n1121), .A2(n1104), .ZN(n2797) );
  CLKBUF_X1 U333 ( .A(n2797), .Z(n2963) );
  INV_X1 U334 ( .A(raddr_b_i[1]), .ZN(n1103) );
  NAND2_X1 U335 ( .A1(n1103), .A2(n1098), .ZN(n1120) );
  INV_X1 U336 ( .A(raddr_b_i[2]), .ZN(n1107) );
  NAND3_X1 U337 ( .A1(raddr_b_i[4]), .A2(raddr_b_i[3]), .A3(n1107), .ZN(n1114)
         );
  NOR2_X1 U338 ( .A1(n1120), .A2(n1114), .ZN(n2980) );
  CLKBUF_X1 U339 ( .A(n2980), .Z(n2764) );
  AOI22_X1 U340 ( .A1(mem[928]), .A2(n2963), .B1(mem[736]), .B2(n2764), .ZN(
        n1102) );
  INV_X1 U341 ( .A(raddr_b_i[4]), .ZN(n1108) );
  NAND3_X1 U342 ( .A1(raddr_b_i[2]), .A2(raddr_b_i[3]), .A3(n1108), .ZN(n1125)
         );
  NAND2_X1 U343 ( .A1(raddr_b_i[1]), .A2(raddr_b_i[0]), .ZN(n1126) );
  NOR2_X1 U344 ( .A1(n1125), .A2(n1126), .ZN(n2952) );
  CLKBUF_X1 U345 ( .A(n2952), .Z(n2833) );
  NOR2_X1 U346 ( .A1(n1104), .A2(n1120), .ZN(n2992) );
  CLKBUF_X1 U347 ( .A(n2992), .Z(n2853) );
  AOI22_X1 U348 ( .A1(mem[448]), .A2(n2833), .B1(mem[864]), .B2(n2853), .ZN(
        n1101) );
  INV_X1 U349 ( .A(raddr_b_i[3]), .ZN(n1105) );
  NAND3_X1 U350 ( .A1(raddr_b_i[2]), .A2(raddr_b_i[4]), .A3(n1105), .ZN(n1127)
         );
  NOR2_X1 U351 ( .A1(n1127), .A2(n1120), .ZN(n2956) );
  CLKBUF_X1 U352 ( .A(n2956), .Z(n2770) );
  NOR2_X1 U353 ( .A1(raddr_b_i[2]), .A2(raddr_b_i[3]), .ZN(n1106) );
  NAND2_X1 U354 ( .A1(n1106), .A2(n1108), .ZN(n1122) );
  NOR2_X1 U355 ( .A1(n1121), .A2(n1122), .ZN(n2990) );
  CLKBUF_X1 U356 ( .A(n2990), .Z(n2775) );
  AOI22_X1 U357 ( .A1(mem[608]), .A2(n2770), .B1(mem[32]), .B2(n2775), .ZN(
        n1100) );
  NOR2_X1 U358 ( .A1(n1121), .A2(n1127), .ZN(n2969) );
  CLKBUF_X1 U359 ( .A(n2969), .Z(n2850) );
  NAND2_X1 U360 ( .A1(mem[672]), .A2(n2850), .ZN(n1099) );
  NAND4_X1 U361 ( .A1(n1102), .A2(n1101), .A3(n1100), .A4(n1099), .ZN(n1135)
         );
  NOR2_X1 U362 ( .A1(n1114), .A2(n1126), .ZN(n2639) );
  CLKBUF_X1 U363 ( .A(n2639), .Z(n2962) );
  NAND2_X1 U364 ( .A1(raddr_b_i[0]), .A2(n1103), .ZN(n1124) );
  NOR2_X1 U365 ( .A1(n1127), .A2(n1124), .ZN(n2967) );
  CLKBUF_X1 U366 ( .A(n2967), .Z(n2796) );
  AOI22_X1 U367 ( .A1(mem[832]), .A2(n2962), .B1(mem[640]), .B2(n2796), .ZN(
        n1112) );
  NOR2_X1 U368 ( .A1(n1104), .A2(n1126), .ZN(n2791) );
  CLKBUF_X1 U369 ( .A(n2791), .Z(n2989) );
  NOR2_X1 U370 ( .A1(n1114), .A2(n1124), .ZN(n2975) );
  CLKBUF_X1 U371 ( .A(n2975), .Z(n2852) );
  AOI22_X1 U372 ( .A1(mem[960]), .A2(n2989), .B1(mem[768]), .B2(n2852), .ZN(
        n1111) );
  NOR2_X1 U373 ( .A1(n1104), .A2(n1124), .ZN(n2785) );
  CLKBUF_X1 U374 ( .A(n2785), .Z(n2968) );
  NAND3_X1 U375 ( .A1(raddr_b_i[2]), .A2(n1108), .A3(n1105), .ZN(n1113) );
  NOR2_X1 U376 ( .A1(n1120), .A2(n1113), .ZN(n2843) );
  CLKBUF_X1 U377 ( .A(n2843), .Z(n2974) );
  AOI22_X1 U378 ( .A1(mem[896]), .A2(n2968), .B1(mem[96]), .B2(n2974), .ZN(
        n1110) );
  NAND2_X1 U379 ( .A1(raddr_b_i[4]), .A2(n1106), .ZN(n1123) );
  NOR2_X1 U380 ( .A1(n1126), .A2(n1123), .ZN(n2986) );
  CLKBUF_X1 U381 ( .A(n2986), .Z(n2765) );
  NAND3_X1 U382 ( .A1(raddr_b_i[3]), .A2(n1108), .A3(n1107), .ZN(n1119) );
  NOR2_X1 U383 ( .A1(n1126), .A2(n1119), .ZN(n2759) );
  CLKBUF_X1 U384 ( .A(n2759), .Z(n2985) );
  AOI22_X1 U385 ( .A1(mem[576]), .A2(n2765), .B1(mem[320]), .B2(n2985), .ZN(
        n1109) );
  NAND4_X1 U386 ( .A1(n1112), .A2(n1111), .A3(n1110), .A4(n1109), .ZN(n1134)
         );
  NOR2_X1 U387 ( .A1(n1120), .A2(n1119), .ZN(n2803) );
  CLKBUF_X1 U388 ( .A(n2803), .Z(n2957) );
  NOR2_X1 U389 ( .A1(n1126), .A2(n1122), .ZN(n2798) );
  AOI22_X1 U390 ( .A1(mem[224]), .A2(n2957), .B1(mem[64]), .B2(n2798), .ZN(
        n1118) );
  NOR2_X1 U391 ( .A1(n1126), .A2(n1113), .ZN(n2776) );
  CLKBUF_X1 U392 ( .A(n2776), .Z(n2977) );
  NOR2_X1 U393 ( .A1(n1124), .A2(n1119), .ZN(n2978) );
  CLKBUF_X1 U394 ( .A(n2978), .Z(n2848) );
  AOI22_X1 U395 ( .A1(mem[192]), .A2(n2977), .B1(mem[256]), .B2(n2848), .ZN(
        n1117) );
  NOR2_X1 U396 ( .A1(n1120), .A2(n1123), .ZN(n2849) );
  NOR2_X1 U397 ( .A1(n1124), .A2(n1113), .ZN(n2859) );
  AOI22_X1 U398 ( .A1(mem[480]), .A2(n2849), .B1(mem[128]), .B2(n2859), .ZN(
        n1116) );
  NOR2_X1 U399 ( .A1(n1121), .A2(n1113), .ZN(n1228) );
  CLKBUF_X1 U400 ( .A(n1228), .Z(n2860) );
  NOR2_X1 U401 ( .A1(n1121), .A2(n1114), .ZN(n2840) );
  AOI22_X1 U402 ( .A1(mem[160]), .A2(n2860), .B1(mem[800]), .B2(n2840), .ZN(
        n1115) );
  NAND4_X1 U403 ( .A1(n1118), .A2(n1117), .A3(n1116), .A4(n1115), .ZN(n1133)
         );
  NOR2_X1 U404 ( .A1(n1121), .A2(n1119), .ZN(n2858) );
  NOR2_X1 U405 ( .A1(n1121), .A2(n1123), .ZN(n2991) );
  AOI22_X1 U406 ( .A1(mem[288]), .A2(n2858), .B1(mem[544]), .B2(n2991), .ZN(
        n1131) );
  NOR2_X1 U407 ( .A1(n1120), .A2(n1125), .ZN(n2842) );
  NOR2_X1 U408 ( .A1(n1121), .A2(n1125), .ZN(n2964) );
  CLKBUF_X1 U409 ( .A(n2964), .Z(n2832) );
  AOI22_X1 U410 ( .A1(mem[352]), .A2(n2842), .B1(mem[416]), .B2(n2832), .ZN(
        n1130) );
  NOR2_X1 U411 ( .A1(n1122), .A2(n1124), .ZN(n2834) );
  NOR2_X1 U412 ( .A1(n1124), .A2(n1123), .ZN(n2988) );
  CLKBUF_X1 U413 ( .A(n2988), .Z(n2835) );
  AOI22_X1 U414 ( .A1(mem[0]), .A2(n2834), .B1(mem[512]), .B2(n2835), .ZN(
        n1129) );
  NOR2_X1 U415 ( .A1(n1125), .A2(n1124), .ZN(n2987) );
  CLKBUF_X1 U416 ( .A(n2987), .Z(n2851) );
  NOR2_X1 U417 ( .A1(n1127), .A2(n1126), .ZN(n2953) );
  CLKBUF_X1 U418 ( .A(n2953), .Z(n2841) );
  AOI22_X1 U419 ( .A1(mem[384]), .A2(n2851), .B1(mem[704]), .B2(n2841), .ZN(
        n1128) );
  NAND4_X1 U420 ( .A1(n1131), .A2(n1130), .A3(n1129), .A4(n1128), .ZN(n1132)
         );
  OR4_X1 U421 ( .A1(n1135), .A2(n1134), .A3(n1133), .A4(n1132), .ZN(
        rdata_b_o[0]) );
  AOI22_X1 U422 ( .A1(n2977), .A2(mem[193]), .B1(n2848), .B2(mem[257]), .ZN(
        n1139) );
  CLKBUF_X1 U423 ( .A(n2991), .Z(n2786) );
  AOI22_X1 U424 ( .A1(n2764), .A2(mem[737]), .B1(n2786), .B2(mem[545]), .ZN(
        n1138) );
  AOI22_X1 U425 ( .A1(n2850), .A2(mem[673]), .B1(n2765), .B2(mem[577]), .ZN(
        n1137) );
  NAND2_X1 U426 ( .A1(n2962), .A2(mem[833]), .ZN(n1136) );
  NAND4_X1 U427 ( .A1(n1139), .A2(n1138), .A3(n1137), .A4(n1136), .ZN(n1155)
         );
  AOI22_X1 U428 ( .A1(n2852), .A2(mem[769]), .B1(n2840), .B2(mem[801]), .ZN(
        n1143) );
  AOI22_X1 U429 ( .A1(n2796), .A2(mem[641]), .B1(n2957), .B2(mem[225]), .ZN(
        n1142) );
  AOI22_X1 U430 ( .A1(n2992), .A2(mem[865]), .B1(n2833), .B2(mem[449]), .ZN(
        n1141) );
  AOI22_X1 U431 ( .A1(n2860), .A2(mem[161]), .B1(n2988), .B2(mem[513]), .ZN(
        n1140) );
  NAND4_X1 U432 ( .A1(n1143), .A2(n1142), .A3(n1141), .A4(n1140), .ZN(n1154)
         );
  AOI22_X1 U433 ( .A1(n2963), .A2(mem[929]), .B1(n2985), .B2(mem[321]), .ZN(
        n1147) );
  AOI22_X1 U434 ( .A1(n2770), .A2(mem[609]), .B1(n2832), .B2(mem[417]), .ZN(
        n1146) );
  AOI22_X1 U435 ( .A1(n2849), .A2(mem[481]), .B1(n2842), .B2(mem[353]), .ZN(
        n1145) );
  AOI22_X1 U436 ( .A1(n2791), .A2(mem[961]), .B1(n2859), .B2(mem[129]), .ZN(
        n1144) );
  NAND4_X1 U437 ( .A1(n1147), .A2(n1146), .A3(n1145), .A4(n1144), .ZN(n1153)
         );
  CLKBUF_X1 U438 ( .A(n2798), .Z(n2966) );
  AOI22_X1 U439 ( .A1(n2974), .A2(mem[97]), .B1(n2966), .B2(mem[65]), .ZN(
        n1151) );
  AOI22_X1 U440 ( .A1(n2968), .A2(mem[897]), .B1(n2858), .B2(mem[289]), .ZN(
        n1150) );
  AOI22_X1 U441 ( .A1(n2834), .A2(mem[1]), .B1(n2841), .B2(mem[705]), .ZN(
        n1149) );
  AOI22_X1 U442 ( .A1(n2775), .A2(mem[33]), .B1(n2851), .B2(mem[385]), .ZN(
        n1148) );
  NAND4_X1 U443 ( .A1(n1151), .A2(n1150), .A3(n1149), .A4(n1148), .ZN(n1152)
         );
  OR4_X1 U444 ( .A1(n1155), .A2(n1154), .A3(n1153), .A4(n1152), .ZN(
        rdata_b_o[1]) );
  AOI22_X1 U445 ( .A1(n2764), .A2(mem[741]), .B1(n2786), .B2(mem[549]), .ZN(
        n1159) );
  AOI22_X1 U446 ( .A1(n2796), .A2(mem[645]), .B1(n2985), .B2(mem[325]), .ZN(
        n1158) );
  AOI22_X1 U447 ( .A1(n2989), .A2(mem[965]), .B1(n2851), .B2(mem[389]), .ZN(
        n1157) );
  NAND2_X1 U448 ( .A1(n2957), .A2(mem[229]), .ZN(n1156) );
  NAND4_X1 U449 ( .A1(n1159), .A2(n1158), .A3(n1157), .A4(n1156), .ZN(n1175)
         );
  AOI22_X1 U450 ( .A1(n2833), .A2(mem[453]), .B1(n2962), .B2(mem[837]), .ZN(
        n1163) );
  AOI22_X1 U451 ( .A1(n2798), .A2(mem[69]), .B1(n2841), .B2(mem[709]), .ZN(
        n1162) );
  AOI22_X1 U452 ( .A1(n2850), .A2(mem[677]), .B1(n2785), .B2(mem[901]), .ZN(
        n1161) );
  AOI22_X1 U453 ( .A1(n2770), .A2(mem[613]), .B1(n2860), .B2(mem[165]), .ZN(
        n1160) );
  NAND4_X1 U454 ( .A1(n1163), .A2(n1162), .A3(n1161), .A4(n1160), .ZN(n1174)
         );
  CLKBUF_X1 U455 ( .A(n2840), .Z(n2955) );
  AOI22_X1 U456 ( .A1(n2849), .A2(mem[485]), .B1(n2955), .B2(mem[805]), .ZN(
        n1167) );
  AOI22_X1 U457 ( .A1(n2775), .A2(mem[37]), .B1(n2835), .B2(mem[517]), .ZN(
        n1166) );
  AOI22_X1 U458 ( .A1(n2974), .A2(mem[101]), .B1(n2978), .B2(mem[261]), .ZN(
        n1165) );
  AOI22_X1 U459 ( .A1(n2797), .A2(mem[933]), .B1(n2977), .B2(mem[197]), .ZN(
        n1164) );
  NAND4_X1 U460 ( .A1(n1167), .A2(n1166), .A3(n1165), .A4(n1164), .ZN(n1173)
         );
  CLKBUF_X1 U461 ( .A(n2842), .Z(n2954) );
  AOI22_X1 U462 ( .A1(n2858), .A2(mem[293]), .B1(n2954), .B2(mem[357]), .ZN(
        n1171) );
  AOI22_X1 U463 ( .A1(n2852), .A2(mem[773]), .B1(n2832), .B2(mem[421]), .ZN(
        n1170) );
  CLKBUF_X1 U464 ( .A(n2834), .Z(n2979) );
  AOI22_X1 U465 ( .A1(n2859), .A2(mem[133]), .B1(n2979), .B2(mem[5]), .ZN(
        n1169) );
  AOI22_X1 U466 ( .A1(n2853), .A2(mem[869]), .B1(n2765), .B2(mem[581]), .ZN(
        n1168) );
  NAND4_X1 U467 ( .A1(n1171), .A2(n1170), .A3(n1169), .A4(n1168), .ZN(n1172)
         );
  OR4_X1 U468 ( .A1(n1175), .A2(n1174), .A3(n1173), .A4(n1172), .ZN(
        rdata_b_o[5]) );
  CLKBUF_X1 U469 ( .A(n2858), .Z(n2976) );
  AOI22_X1 U470 ( .A1(n2775), .A2(mem[36]), .B1(n2976), .B2(mem[292]), .ZN(
        n1179) );
  AOI22_X1 U471 ( .A1(n2850), .A2(mem[676]), .B1(n2954), .B2(mem[356]), .ZN(
        n1178) );
  AOI22_X1 U472 ( .A1(n2966), .A2(mem[68]), .B1(n2860), .B2(mem[164]), .ZN(
        n1177) );
  NAND2_X1 U473 ( .A1(n2963), .A2(mem[932]), .ZN(n1176) );
  NAND4_X1 U474 ( .A1(n1179), .A2(n1178), .A3(n1177), .A4(n1176), .ZN(n1195)
         );
  AOI22_X1 U475 ( .A1(n2852), .A2(mem[772]), .B1(n2968), .B2(mem[900]), .ZN(
        n1183) );
  AOI22_X1 U476 ( .A1(n2803), .A2(mem[228]), .B1(n2786), .B2(mem[548]), .ZN(
        n1182) );
  AOI22_X1 U477 ( .A1(n2978), .A2(mem[260]), .B1(n2979), .B2(mem[4]), .ZN(
        n1181) );
  AOI22_X1 U478 ( .A1(n2985), .A2(mem[324]), .B1(n2955), .B2(mem[804]), .ZN(
        n1180) );
  NAND4_X1 U479 ( .A1(n1183), .A2(n1182), .A3(n1181), .A4(n1180), .ZN(n1194)
         );
  AOI22_X1 U480 ( .A1(n2796), .A2(mem[644]), .B1(n2849), .B2(mem[484]), .ZN(
        n1187) );
  AOI22_X1 U481 ( .A1(n2962), .A2(mem[836]), .B1(n2776), .B2(mem[196]), .ZN(
        n1186) );
  CLKBUF_X1 U482 ( .A(n2859), .Z(n2951) );
  AOI22_X1 U483 ( .A1(n2952), .A2(mem[452]), .B1(n2951), .B2(mem[132]), .ZN(
        n1185) );
  AOI22_X1 U484 ( .A1(n2988), .A2(mem[516]), .B1(n2841), .B2(mem[708]), .ZN(
        n1184) );
  NAND4_X1 U485 ( .A1(n1187), .A2(n1186), .A3(n1185), .A4(n1184), .ZN(n1193)
         );
  AOI22_X1 U486 ( .A1(n2764), .A2(mem[740]), .B1(n2992), .B2(mem[868]), .ZN(
        n1191) );
  AOI22_X1 U487 ( .A1(n2791), .A2(mem[964]), .B1(n2851), .B2(mem[388]), .ZN(
        n1190) );
  AOI22_X1 U488 ( .A1(n2956), .A2(mem[612]), .B1(n2964), .B2(mem[420]), .ZN(
        n1189) );
  AOI22_X1 U489 ( .A1(n2974), .A2(mem[100]), .B1(n2765), .B2(mem[580]), .ZN(
        n1188) );
  NAND4_X1 U490 ( .A1(n1191), .A2(n1190), .A3(n1189), .A4(n1188), .ZN(n1192)
         );
  OR4_X1 U491 ( .A1(n1195), .A2(n1194), .A3(n1193), .A4(n1192), .ZN(
        rdata_b_o[4]) );
  AOI22_X1 U492 ( .A1(n2974), .A2(mem[99]), .B1(n2765), .B2(mem[579]), .ZN(
        n1199) );
  AOI22_X1 U493 ( .A1(n2796), .A2(mem[643]), .B1(n2786), .B2(mem[547]), .ZN(
        n1198) );
  AOI22_X1 U494 ( .A1(n2955), .A2(mem[803]), .B1(n2832), .B2(mem[419]), .ZN(
        n1197) );
  NAND2_X1 U495 ( .A1(n2963), .A2(mem[931]), .ZN(n1196) );
  NAND4_X1 U496 ( .A1(n1199), .A2(n1198), .A3(n1197), .A4(n1196), .ZN(n1215)
         );
  AOI22_X1 U497 ( .A1(n2849), .A2(mem[483]), .B1(n1228), .B2(mem[163]), .ZN(
        n1203) );
  AOI22_X1 U498 ( .A1(n2770), .A2(mem[611]), .B1(n2962), .B2(mem[835]), .ZN(
        n1202) );
  AOI22_X1 U499 ( .A1(n2852), .A2(mem[771]), .B1(n2978), .B2(mem[259]), .ZN(
        n1201) );
  AOI22_X1 U500 ( .A1(n2969), .A2(mem[675]), .B1(n2835), .B2(mem[515]), .ZN(
        n1200) );
  NAND4_X1 U501 ( .A1(n1203), .A2(n1202), .A3(n1201), .A4(n1200), .ZN(n1214)
         );
  AOI22_X1 U502 ( .A1(n2980), .A2(mem[739]), .B1(n2977), .B2(mem[195]), .ZN(
        n1207) );
  AOI22_X1 U503 ( .A1(n2992), .A2(mem[867]), .B1(n2954), .B2(mem[355]), .ZN(
        n1206) );
  AOI22_X1 U504 ( .A1(n2858), .A2(mem[291]), .B1(n2851), .B2(mem[387]), .ZN(
        n1205) );
  AOI22_X1 U505 ( .A1(n2833), .A2(mem[451]), .B1(n2990), .B2(mem[35]), .ZN(
        n1204) );
  NAND4_X1 U506 ( .A1(n1207), .A2(n1206), .A3(n1205), .A4(n1204), .ZN(n1213)
         );
  AOI22_X1 U507 ( .A1(n2985), .A2(mem[323]), .B1(n2979), .B2(mem[3]), .ZN(
        n1211) );
  AOI22_X1 U508 ( .A1(n2968), .A2(mem[899]), .B1(n2798), .B2(mem[67]), .ZN(
        n1210) );
  AOI22_X1 U509 ( .A1(n2859), .A2(mem[131]), .B1(n2841), .B2(mem[707]), .ZN(
        n1209) );
  AOI22_X1 U510 ( .A1(n2989), .A2(mem[963]), .B1(n2803), .B2(mem[227]), .ZN(
        n1208) );
  NAND4_X1 U511 ( .A1(n1211), .A2(n1210), .A3(n1209), .A4(n1208), .ZN(n1212)
         );
  OR4_X1 U512 ( .A1(n1215), .A2(n1214), .A3(n1213), .A4(n1212), .ZN(
        rdata_b_o[3]) );
  AOI22_X1 U513 ( .A1(n2765), .A2(mem[578]), .B1(n2951), .B2(mem[130]), .ZN(
        n1219) );
  AOI22_X1 U514 ( .A1(n2989), .A2(mem[962]), .B1(n2976), .B2(mem[290]), .ZN(
        n1218) );
  AOI22_X1 U515 ( .A1(n2954), .A2(mem[354]), .B1(n2841), .B2(mem[706]), .ZN(
        n1217) );
  NAND2_X1 U516 ( .A1(n2848), .A2(mem[258]), .ZN(n1216) );
  NAND4_X1 U517 ( .A1(n1219), .A2(n1218), .A3(n1217), .A4(n1216), .ZN(n1236)
         );
  AOI22_X1 U518 ( .A1(n2852), .A2(mem[770]), .B1(n2803), .B2(mem[226]), .ZN(
        n1223) );
  AOI22_X1 U519 ( .A1(n2849), .A2(mem[482]), .B1(n2955), .B2(mem[802]), .ZN(
        n1222) );
  AOI22_X1 U520 ( .A1(n2775), .A2(mem[34]), .B1(n2977), .B2(mem[194]), .ZN(
        n1221) );
  AOI22_X1 U521 ( .A1(n2988), .A2(mem[514]), .B1(n2834), .B2(mem[2]), .ZN(
        n1220) );
  NAND4_X1 U522 ( .A1(n1223), .A2(n1222), .A3(n1221), .A4(n1220), .ZN(n1235)
         );
  AOI22_X1 U523 ( .A1(n2956), .A2(mem[610]), .B1(n2785), .B2(mem[898]), .ZN(
        n1227) );
  AOI22_X1 U524 ( .A1(n2764), .A2(mem[738]), .B1(n2952), .B2(mem[450]), .ZN(
        n1226) );
  AOI22_X1 U525 ( .A1(n2974), .A2(mem[98]), .B1(n2786), .B2(mem[546]), .ZN(
        n1225) );
  AOI22_X1 U526 ( .A1(n2963), .A2(mem[930]), .B1(n2759), .B2(mem[322]), .ZN(
        n1224) );
  NAND4_X1 U527 ( .A1(n1227), .A2(n1226), .A3(n1225), .A4(n1224), .ZN(n1234)
         );
  AOI22_X1 U528 ( .A1(n2969), .A2(mem[674]), .B1(n2964), .B2(mem[418]), .ZN(
        n1232) );
  AOI22_X1 U529 ( .A1(n2992), .A2(mem[866]), .B1(n2860), .B2(mem[162]), .ZN(
        n1231) );
  AOI22_X1 U530 ( .A1(n2962), .A2(mem[834]), .B1(n2851), .B2(mem[386]), .ZN(
        n1230) );
  AOI22_X1 U531 ( .A1(n2796), .A2(mem[642]), .B1(n2966), .B2(mem[66]), .ZN(
        n1229) );
  NAND4_X1 U532 ( .A1(n1232), .A2(n1231), .A3(n1230), .A4(n1229), .ZN(n1233)
         );
  OR4_X1 U533 ( .A1(n1236), .A2(n1235), .A3(n1234), .A4(n1233), .ZN(
        rdata_b_o[2]) );
  AOI22_X1 U534 ( .A1(n2765), .A2(mem[585]), .B1(n2977), .B2(mem[201]), .ZN(
        n1240) );
  AOI22_X1 U535 ( .A1(n2955), .A2(mem[809]), .B1(n2954), .B2(mem[361]), .ZN(
        n1239) );
  AOI22_X1 U536 ( .A1(n2966), .A2(mem[73]), .B1(n2951), .B2(mem[137]), .ZN(
        n1238) );
  CLKBUF_X1 U537 ( .A(n2849), .Z(n2965) );
  NAND2_X1 U538 ( .A1(n2965), .A2(mem[489]), .ZN(n1237) );
  NAND4_X1 U539 ( .A1(n1240), .A2(n1239), .A3(n1238), .A4(n1237), .ZN(n1256)
         );
  AOI22_X1 U540 ( .A1(n2796), .A2(mem[649]), .B1(n2976), .B2(mem[297]), .ZN(
        n1244) );
  AOI22_X1 U541 ( .A1(n2850), .A2(mem[681]), .B1(n2770), .B2(mem[617]), .ZN(
        n1243) );
  AOI22_X1 U542 ( .A1(n2957), .A2(mem[233]), .B1(n2786), .B2(mem[553]), .ZN(
        n1242) );
  AOI22_X1 U543 ( .A1(n2968), .A2(mem[905]), .B1(n2835), .B2(mem[521]), .ZN(
        n1241) );
  NAND4_X1 U544 ( .A1(n1244), .A2(n1243), .A3(n1242), .A4(n1241), .ZN(n1255)
         );
  AOI22_X1 U545 ( .A1(n2775), .A2(mem[41]), .B1(n2979), .B2(mem[9]), .ZN(n1248) );
  AOI22_X1 U546 ( .A1(n2962), .A2(mem[841]), .B1(n2985), .B2(mem[329]), .ZN(
        n1247) );
  AOI22_X1 U547 ( .A1(n2833), .A2(mem[457]), .B1(n2791), .B2(mem[969]), .ZN(
        n1246) );
  AOI22_X1 U548 ( .A1(n2764), .A2(mem[745]), .B1(n2832), .B2(mem[425]), .ZN(
        n1245) );
  NAND4_X1 U549 ( .A1(n1248), .A2(n1247), .A3(n1246), .A4(n1245), .ZN(n1254)
         );
  AOI22_X1 U550 ( .A1(n2978), .A2(mem[265]), .B1(n2841), .B2(mem[713]), .ZN(
        n1252) );
  AOI22_X1 U551 ( .A1(n2853), .A2(mem[873]), .B1(n2851), .B2(mem[393]), .ZN(
        n1251) );
  AOI22_X1 U552 ( .A1(n2974), .A2(mem[105]), .B1(n1228), .B2(mem[169]), .ZN(
        n1250) );
  AOI22_X1 U553 ( .A1(n2797), .A2(mem[937]), .B1(n2852), .B2(mem[777]), .ZN(
        n1249) );
  NAND4_X1 U554 ( .A1(n1252), .A2(n1251), .A3(n1250), .A4(n1249), .ZN(n1253)
         );
  OR4_X1 U555 ( .A1(n1256), .A2(n1255), .A3(n1254), .A4(n1253), .ZN(
        rdata_b_o[9]) );
  AOI22_X1 U556 ( .A1(n2974), .A2(mem[104]), .B1(n2841), .B2(mem[712]), .ZN(
        n1260) );
  AOI22_X1 U557 ( .A1(n2962), .A2(mem[840]), .B1(n2965), .B2(mem[488]), .ZN(
        n1259) );
  AOI22_X1 U558 ( .A1(n2853), .A2(mem[872]), .B1(n2954), .B2(mem[360]), .ZN(
        n1258) );
  NAND2_X1 U559 ( .A1(n2963), .A2(mem[936]), .ZN(n1257) );
  NAND4_X1 U560 ( .A1(n1260), .A2(n1259), .A3(n1258), .A4(n1257), .ZN(n1276)
         );
  AOI22_X1 U561 ( .A1(n2833), .A2(mem[456]), .B1(n2786), .B2(mem[552]), .ZN(
        n1264) );
  AOI22_X1 U562 ( .A1(n2986), .A2(mem[584]), .B1(n2851), .B2(mem[392]), .ZN(
        n1263) );
  AOI22_X1 U563 ( .A1(n2764), .A2(mem[744]), .B1(n2989), .B2(mem[968]), .ZN(
        n1262) );
  AOI22_X1 U564 ( .A1(n2759), .A2(mem[328]), .B1(n2860), .B2(mem[168]), .ZN(
        n1261) );
  NAND4_X1 U565 ( .A1(n1264), .A2(n1263), .A3(n1262), .A4(n1261), .ZN(n1275)
         );
  AOI22_X1 U566 ( .A1(n2775), .A2(mem[40]), .B1(n2832), .B2(mem[424]), .ZN(
        n1268) );
  AOI22_X1 U567 ( .A1(n2852), .A2(mem[776]), .B1(n2957), .B2(mem[232]), .ZN(
        n1267) );
  AOI22_X1 U568 ( .A1(n2858), .A2(mem[296]), .B1(n2835), .B2(mem[520]), .ZN(
        n1266) );
  AOI22_X1 U569 ( .A1(n2770), .A2(mem[616]), .B1(n2840), .B2(mem[808]), .ZN(
        n1265) );
  NAND4_X1 U570 ( .A1(n1268), .A2(n1267), .A3(n1266), .A4(n1265), .ZN(n1274)
         );
  AOI22_X1 U571 ( .A1(n2850), .A2(mem[680]), .B1(n2979), .B2(mem[8]), .ZN(
        n1272) );
  AOI22_X1 U572 ( .A1(n2798), .A2(mem[72]), .B1(n2848), .B2(mem[264]), .ZN(
        n1271) );
  AOI22_X1 U573 ( .A1(n2968), .A2(mem[904]), .B1(n2951), .B2(mem[136]), .ZN(
        n1270) );
  AOI22_X1 U574 ( .A1(n2796), .A2(mem[648]), .B1(n2776), .B2(mem[200]), .ZN(
        n1269) );
  NAND4_X1 U575 ( .A1(n1272), .A2(n1271), .A3(n1270), .A4(n1269), .ZN(n1273)
         );
  OR4_X1 U576 ( .A1(n1276), .A2(n1275), .A3(n1274), .A4(n1273), .ZN(
        rdata_b_o[8]) );
  AOI22_X1 U577 ( .A1(n2803), .A2(mem[235]), .B1(n2976), .B2(mem[299]), .ZN(
        n1280) );
  AOI22_X1 U578 ( .A1(n2985), .A2(mem[331]), .B1(n2954), .B2(mem[363]), .ZN(
        n1279) );
  AOI22_X1 U579 ( .A1(n2765), .A2(mem[587]), .B1(n2835), .B2(mem[523]), .ZN(
        n1278) );
  NAND2_X1 U580 ( .A1(n2775), .A2(mem[43]), .ZN(n1277) );
  NAND4_X1 U581 ( .A1(n1280), .A2(n1279), .A3(n1278), .A4(n1277), .ZN(n1296)
         );
  AOI22_X1 U582 ( .A1(n2977), .A2(mem[203]), .B1(n2841), .B2(mem[715]), .ZN(
        n1284) );
  AOI22_X1 U583 ( .A1(n2764), .A2(mem[747]), .B1(n1228), .B2(mem[171]), .ZN(
        n1283) );
  AOI22_X1 U584 ( .A1(n2796), .A2(mem[651]), .B1(n2978), .B2(mem[267]), .ZN(
        n1282) );
  AOI22_X1 U585 ( .A1(n2849), .A2(mem[491]), .B1(n2955), .B2(mem[811]), .ZN(
        n1281) );
  NAND4_X1 U586 ( .A1(n1284), .A2(n1283), .A3(n1282), .A4(n1281), .ZN(n1295)
         );
  AOI22_X1 U587 ( .A1(n2850), .A2(mem[683]), .B1(n2851), .B2(mem[395]), .ZN(
        n1288) );
  AOI22_X1 U588 ( .A1(n2791), .A2(mem[971]), .B1(n2785), .B2(mem[907]), .ZN(
        n1287) );
  AOI22_X1 U589 ( .A1(n2852), .A2(mem[779]), .B1(n2843), .B2(mem[107]), .ZN(
        n1286) );
  AOI22_X1 U590 ( .A1(n2770), .A2(mem[619]), .B1(n2834), .B2(mem[11]), .ZN(
        n1285) );
  NAND4_X1 U591 ( .A1(n1288), .A2(n1287), .A3(n1286), .A4(n1285), .ZN(n1294)
         );
  AOI22_X1 U592 ( .A1(n2853), .A2(mem[875]), .B1(n2952), .B2(mem[459]), .ZN(
        n1292) );
  AOI22_X1 U593 ( .A1(n2859), .A2(mem[139]), .B1(n2964), .B2(mem[427]), .ZN(
        n1291) );
  AOI22_X1 U594 ( .A1(n2797), .A2(mem[939]), .B1(n2798), .B2(mem[75]), .ZN(
        n1290) );
  AOI22_X1 U595 ( .A1(n2639), .A2(mem[843]), .B1(n2991), .B2(mem[555]), .ZN(
        n1289) );
  NAND4_X1 U596 ( .A1(n1292), .A2(n1291), .A3(n1290), .A4(n1289), .ZN(n1293)
         );
  OR4_X1 U597 ( .A1(n1296), .A2(n1295), .A3(n1294), .A4(n1293), .ZN(
        rdata_b_o[11]) );
  AOI22_X1 U598 ( .A1(n2832), .A2(mem[422]), .B1(n2835), .B2(mem[518]), .ZN(
        n1300) );
  AOI22_X1 U599 ( .A1(n2850), .A2(mem[678]), .B1(n2989), .B2(mem[966]), .ZN(
        n1299) );
  AOI22_X1 U600 ( .A1(n2985), .A2(mem[326]), .B1(n2954), .B2(mem[358]), .ZN(
        n1298) );
  NAND2_X1 U601 ( .A1(n2966), .A2(mem[70]), .ZN(n1297) );
  NAND4_X1 U602 ( .A1(n1300), .A2(n1299), .A3(n1298), .A4(n1297), .ZN(n1316)
         );
  AOI22_X1 U603 ( .A1(n2775), .A2(mem[38]), .B1(n2965), .B2(mem[486]), .ZN(
        n1304) );
  AOI22_X1 U604 ( .A1(n2974), .A2(mem[102]), .B1(n2955), .B2(mem[806]), .ZN(
        n1303) );
  AOI22_X1 U605 ( .A1(n2796), .A2(mem[646]), .B1(n2848), .B2(mem[262]), .ZN(
        n1302) );
  AOI22_X1 U606 ( .A1(n2977), .A2(mem[198]), .B1(n2976), .B2(mem[294]), .ZN(
        n1301) );
  NAND4_X1 U607 ( .A1(n1304), .A2(n1303), .A3(n1302), .A4(n1301), .ZN(n1315)
         );
  AOI22_X1 U608 ( .A1(n2962), .A2(mem[838]), .B1(n2765), .B2(mem[582]), .ZN(
        n1308) );
  AOI22_X1 U609 ( .A1(n2852), .A2(mem[774]), .B1(n2851), .B2(mem[390]), .ZN(
        n1307) );
  AOI22_X1 U610 ( .A1(n2963), .A2(mem[934]), .B1(n2764), .B2(mem[742]), .ZN(
        n1306) );
  AOI22_X1 U611 ( .A1(n2968), .A2(mem[902]), .B1(n2951), .B2(mem[134]), .ZN(
        n1305) );
  NAND4_X1 U612 ( .A1(n1308), .A2(n1307), .A3(n1306), .A4(n1305), .ZN(n1314)
         );
  AOI22_X1 U613 ( .A1(n2833), .A2(mem[454]), .B1(n2957), .B2(mem[230]), .ZN(
        n1312) );
  AOI22_X1 U614 ( .A1(n2770), .A2(mem[614]), .B1(n2979), .B2(mem[6]), .ZN(
        n1311) );
  AOI22_X1 U615 ( .A1(n2860), .A2(mem[166]), .B1(n2841), .B2(mem[710]), .ZN(
        n1310) );
  AOI22_X1 U616 ( .A1(n2853), .A2(mem[870]), .B1(n2786), .B2(mem[550]), .ZN(
        n1309) );
  NAND4_X1 U617 ( .A1(n1312), .A2(n1311), .A3(n1310), .A4(n1309), .ZN(n1313)
         );
  OR4_X1 U618 ( .A1(n1316), .A2(n1315), .A3(n1314), .A4(n1313), .ZN(
        rdata_b_o[6]) );
  AOI22_X1 U619 ( .A1(n2853), .A2(mem[880]), .B1(n2979), .B2(mem[16]), .ZN(
        n1320) );
  AOI22_X1 U620 ( .A1(n2860), .A2(mem[176]), .B1(n2991), .B2(mem[560]), .ZN(
        n1319) );
  AOI22_X1 U621 ( .A1(n2765), .A2(mem[592]), .B1(n2835), .B2(mem[528]), .ZN(
        n1318) );
  NAND2_X1 U622 ( .A1(n2951), .A2(mem[144]), .ZN(n1317) );
  NAND4_X1 U623 ( .A1(n1320), .A2(n1319), .A3(n1318), .A4(n1317), .ZN(n1336)
         );
  AOI22_X1 U624 ( .A1(n2963), .A2(mem[944]), .B1(n2764), .B2(mem[752]), .ZN(
        n1324) );
  AOI22_X1 U625 ( .A1(n2989), .A2(mem[976]), .B1(n2976), .B2(mem[304]), .ZN(
        n1323) );
  AOI22_X1 U626 ( .A1(n2990), .A2(mem[48]), .B1(n2964), .B2(mem[432]), .ZN(
        n1322) );
  AOI22_X1 U627 ( .A1(n2957), .A2(mem[240]), .B1(n2841), .B2(mem[720]), .ZN(
        n1321) );
  NAND4_X1 U628 ( .A1(n1324), .A2(n1323), .A3(n1322), .A4(n1321), .ZN(n1335)
         );
  AOI22_X1 U629 ( .A1(n2849), .A2(mem[496]), .B1(n2851), .B2(mem[400]), .ZN(
        n1328) );
  AOI22_X1 U630 ( .A1(n2759), .A2(mem[336]), .B1(n2842), .B2(mem[368]), .ZN(
        n1327) );
  AOI22_X1 U631 ( .A1(n2967), .A2(mem[656]), .B1(n2785), .B2(mem[912]), .ZN(
        n1326) );
  AOI22_X1 U632 ( .A1(n2770), .A2(mem[624]), .B1(n2962), .B2(mem[848]), .ZN(
        n1325) );
  NAND4_X1 U633 ( .A1(n1328), .A2(n1327), .A3(n1326), .A4(n1325), .ZN(n1334)
         );
  AOI22_X1 U634 ( .A1(n2843), .A2(mem[112]), .B1(n2966), .B2(mem[80]), .ZN(
        n1332) );
  AOI22_X1 U635 ( .A1(n2850), .A2(mem[688]), .B1(n2852), .B2(mem[784]), .ZN(
        n1331) );
  AOI22_X1 U636 ( .A1(n2833), .A2(mem[464]), .B1(n2848), .B2(mem[272]), .ZN(
        n1330) );
  AOI22_X1 U637 ( .A1(n2776), .A2(mem[208]), .B1(n2955), .B2(mem[816]), .ZN(
        n1329) );
  NAND4_X1 U638 ( .A1(n1332), .A2(n1331), .A3(n1330), .A4(n1329), .ZN(n1333)
         );
  OR4_X1 U639 ( .A1(n1336), .A2(n1335), .A3(n1334), .A4(n1333), .ZN(
        rdata_b_o[16]) );
  INV_X1 U640 ( .A(raddr_c_i[0]), .ZN(n1344) );
  NAND3_X1 U641 ( .A1(raddr_c_i[4]), .A2(raddr_c_i[3]), .A3(raddr_c_i[2]), 
        .ZN(n1345) );
  NOR2_X1 U642 ( .A1(n1362), .A2(n1345), .ZN(n1403) );
  INV_X1 U643 ( .A(raddr_c_i[4]), .ZN(n1343) );
  INV_X1 U644 ( .A(raddr_c_i[3]), .ZN(n1346) );
  NAND3_X1 U645 ( .A1(raddr_c_i[2]), .A2(n1343), .A3(n1346), .ZN(n1351) );
  NOR2_X1 U646 ( .A1(n1358), .A2(n1351), .ZN(n1408) );
  AOI22_X1 U647 ( .A1(n2869), .A2(mem[912]), .B1(n1043), .B2(mem[112]), .ZN(
        n1341) );
  INV_X1 U648 ( .A(raddr_c_i[2]), .ZN(n1342) );
  NAND3_X1 U649 ( .A1(raddr_c_i[3]), .A2(raddr_c_i[4]), .A3(n1342), .ZN(n1363)
         );
  NAND2_X1 U650 ( .A1(raddr_c_i[1]), .A2(raddr_c_i[0]), .ZN(n1361) );
  NOR2_X1 U651 ( .A1(n1363), .A2(n1361), .ZN(n1516) );
  NOR2_X1 U652 ( .A1(raddr_c_i[3]), .A2(raddr_c_i[2]), .ZN(n1337) );
  NAND2_X1 U653 ( .A1(n1337), .A2(n1343), .ZN(n1360) );
  NOR2_X1 U654 ( .A1(n1360), .A2(n1362), .ZN(n1751) );
  AOI22_X1 U655 ( .A1(n1050), .A2(mem[848]), .B1(n1045), .B2(mem[16]), .ZN(
        n1340) );
  NAND2_X1 U656 ( .A1(raddr_c_i[4]), .A2(n1337), .ZN(n1365) );
  NOR2_X1 U657 ( .A1(n1358), .A2(n1365), .ZN(n1740) );
  NOR2_X1 U658 ( .A1(n1361), .A2(n1365), .ZN(n1752) );
  AOI22_X1 U659 ( .A1(n2062), .A2(mem[496]), .B1(n2433), .B2(mem[592]), .ZN(
        n1339) );
  NOR2_X1 U660 ( .A1(n1361), .A2(n1345), .ZN(n1750) );
  NAND2_X1 U661 ( .A1(n1055), .A2(mem[976]), .ZN(n1338) );
  NAND4_X1 U662 ( .A1(n1341), .A2(n1340), .A3(n1339), .A4(n1338), .ZN(n1373)
         );
  NAND3_X1 U663 ( .A1(raddr_c_i[3]), .A2(raddr_c_i[2]), .A3(n1343), .ZN(n1352)
         );
  NOR2_X1 U664 ( .A1(n1361), .A2(n1352), .ZN(n1776) );
  NAND3_X1 U665 ( .A1(raddr_c_i[3]), .A2(n1343), .A3(n1342), .ZN(n1359) );
  NOR2_X1 U666 ( .A1(n1362), .A2(n1359), .ZN(n1738) );
  AOI22_X1 U667 ( .A1(n1046), .A2(mem[464]), .B1(n1049), .B2(mem[272]), .ZN(
        n1350) );
  NOR2_X1 U668 ( .A1(n1361), .A2(n1351), .ZN(n1511) );
  NOR2_X1 U669 ( .A1(n1358), .A2(n1345), .ZN(n1415) );
  AOI22_X1 U670 ( .A1(n1040), .A2(mem[208]), .B1(n1415), .B2(mem[880]), .ZN(
        n1349) );
  NOR2_X1 U671 ( .A1(n1364), .A2(n1360), .ZN(n1414) );
  NOR2_X1 U672 ( .A1(n1364), .A2(n1345), .ZN(n1402) );
  AOI22_X1 U673 ( .A1(n3001), .A2(mem[48]), .B1(n1402), .B2(mem[944]), .ZN(
        n1348) );
  NAND3_X1 U674 ( .A1(raddr_c_i[4]), .A2(raddr_c_i[2]), .A3(n1346), .ZN(n1357)
         );
  NOR2_X1 U675 ( .A1(n1357), .A2(n1364), .ZN(n1431) );
  NOR2_X1 U676 ( .A1(n1362), .A2(n1351), .ZN(n1396) );
  AOI22_X1 U677 ( .A1(n1052), .A2(mem[688]), .B1(n1051), .B2(mem[144]), .ZN(
        n1347) );
  NAND4_X1 U678 ( .A1(n1350), .A2(n1349), .A3(n1348), .A4(n1347), .ZN(n1372)
         );
  NOR2_X1 U679 ( .A1(n1357), .A2(n1362), .ZN(n2067) );
  NOR2_X1 U680 ( .A1(n1363), .A2(n1358), .ZN(n1461) );
  AOI22_X1 U681 ( .A1(n2578), .A2(mem[656]), .B1(n2705), .B2(mem[752]), .ZN(
        n1356) );
  NOR2_X1 U682 ( .A1(n1358), .A2(n1352), .ZN(n1424) );
  NOR2_X1 U683 ( .A1(n1361), .A2(n1357), .ZN(n1452) );
  AOI22_X1 U684 ( .A1(n2874), .A2(mem[368]), .B1(n3015), .B2(mem[720]), .ZN(
        n1355) );
  NOR2_X1 U685 ( .A1(n1362), .A2(n1352), .ZN(n1786) );
  NOR2_X1 U686 ( .A1(n1365), .A2(n1362), .ZN(n1474) );
  AOI22_X1 U687 ( .A1(n1033), .A2(mem[400]), .B1(n2750), .B2(mem[528]), .ZN(
        n1354) );
  NOR2_X1 U688 ( .A1(n1364), .A2(n1351), .ZN(n1430) );
  NOR2_X1 U689 ( .A1(n1364), .A2(n1352), .ZN(n1521) );
  AOI22_X1 U690 ( .A1(n1041), .A2(mem[176]), .B1(n1053), .B2(mem[432]), .ZN(
        n1353) );
  NAND4_X1 U691 ( .A1(n1356), .A2(n1355), .A3(n1354), .A4(n1353), .ZN(n1371)
         );
  NOR2_X1 U692 ( .A1(n1357), .A2(n1358), .ZN(n1745) );
  NOR2_X1 U693 ( .A1(n1358), .A2(n1359), .ZN(n1781) );
  AOI22_X1 U694 ( .A1(n2668), .A2(mem[624]), .B1(n1042), .B2(mem[240]), .ZN(
        n1369) );
  NOR2_X1 U695 ( .A1(n1364), .A2(n1359), .ZN(n1395) );
  NOR2_X1 U696 ( .A1(n1363), .A2(n1364), .ZN(n1401) );
  AOI22_X1 U697 ( .A1(n3016), .A2(mem[304]), .B1(n1044), .B2(mem[816]), .ZN(
        n1368) );
  NOR2_X1 U698 ( .A1(n1361), .A2(n1359), .ZN(n1409) );
  NOR2_X1 U699 ( .A1(n1361), .A2(n1360), .ZN(n1429) );
  AOI22_X1 U700 ( .A1(n1054), .A2(mem[336]), .B1(n1047), .B2(mem[80]), .ZN(
        n1367) );
  NOR2_X1 U701 ( .A1(n1363), .A2(n1362), .ZN(n1739) );
  NOR2_X1 U702 ( .A1(n1365), .A2(n1364), .ZN(n1394) );
  AOI22_X1 U703 ( .A1(n1048), .A2(mem[784]), .B1(n3010), .B2(mem[560]), .ZN(
        n1366) );
  NAND4_X1 U704 ( .A1(n1369), .A2(n1368), .A3(n1367), .A4(n1366), .ZN(n1370)
         );
  OR4_X1 U705 ( .A1(n1373), .A2(n1372), .A3(n1371), .A4(n1370), .ZN(
        rdata_c_o[16]) );
  AOI22_X1 U706 ( .A1(mem[608]), .A2(n2668), .B1(mem[480]), .B2(n2062), .ZN(
        n1377) );
  AOI22_X1 U707 ( .A1(mem[576]), .A2(n2433), .B1(mem[32]), .B2(n1414), .ZN(
        n1376) );
  AOI22_X1 U708 ( .A1(mem[0]), .A2(n1045), .B1(mem[288]), .B2(n1395), .ZN(
        n1375) );
  NAND2_X1 U709 ( .A1(mem[832]), .A2(n1050), .ZN(n1374) );
  NAND4_X1 U710 ( .A1(n1377), .A2(n1376), .A3(n1375), .A4(n1374), .ZN(n1393)
         );
  AOI22_X1 U711 ( .A1(mem[352]), .A2(n1424), .B1(mem[384]), .B2(n1033), .ZN(
        n1381) );
  AOI22_X1 U712 ( .A1(mem[960]), .A2(n1055), .B1(mem[928]), .B2(n1039), .ZN(
        n1380) );
  AOI22_X1 U713 ( .A1(mem[160]), .A2(n1041), .B1(mem[896]), .B2(n2869), .ZN(
        n1379) );
  AOI22_X1 U714 ( .A1(mem[224]), .A2(n1042), .B1(mem[192]), .B2(n1040), .ZN(
        n1378) );
  NAND4_X1 U715 ( .A1(n1381), .A2(n1380), .A3(n1379), .A4(n1378), .ZN(n1392)
         );
  AOI22_X1 U716 ( .A1(mem[704]), .A2(n3015), .B1(mem[320]), .B2(n1054), .ZN(
        n1385) );
  AOI22_X1 U717 ( .A1(mem[416]), .A2(n1053), .B1(mem[640]), .B2(n2578), .ZN(
        n1384) );
  AOI22_X1 U718 ( .A1(mem[736]), .A2(n2705), .B1(mem[672]), .B2(n1052), .ZN(
        n1383) );
  AOI22_X1 U719 ( .A1(mem[512]), .A2(n2750), .B1(mem[768]), .B2(n1048), .ZN(
        n1382) );
  NAND4_X1 U720 ( .A1(n1385), .A2(n1384), .A3(n1383), .A4(n1382), .ZN(n1391)
         );
  AOI22_X1 U721 ( .A1(mem[64]), .A2(n1047), .B1(mem[448]), .B2(n1046), .ZN(
        n1389) );
  AOI22_X1 U722 ( .A1(mem[800]), .A2(n1044), .B1(mem[544]), .B2(n3010), .ZN(
        n1388) );
  AOI22_X1 U723 ( .A1(mem[96]), .A2(n1043), .B1(mem[864]), .B2(n1056), .ZN(
        n1387) );
  AOI22_X1 U724 ( .A1(mem[256]), .A2(n1049), .B1(mem[128]), .B2(n1051), .ZN(
        n1386) );
  NAND4_X1 U725 ( .A1(n1389), .A2(n1388), .A3(n1387), .A4(n1386), .ZN(n1390)
         );
  OR4_X1 U726 ( .A1(n1393), .A2(n1392), .A3(n1391), .A4(n1390), .ZN(
        rdata_c_o[0]) );
  AOI22_X1 U727 ( .A1(n2874), .A2(mem[357]), .B1(n3010), .B2(mem[549]), .ZN(
        n1400) );
  AOI22_X1 U728 ( .A1(n1050), .A2(mem[837]), .B1(n1395), .B2(mem[293]), .ZN(
        n1399) );
  AOI22_X1 U729 ( .A1(n2433), .A2(mem[581]), .B1(n1049), .B2(mem[261]), .ZN(
        n1398) );
  NAND2_X1 U730 ( .A1(n1051), .A2(mem[133]), .ZN(n1397) );
  NAND4_X1 U731 ( .A1(n1400), .A2(n1399), .A3(n1398), .A4(n1397), .ZN(n1423)
         );
  AOI22_X1 U732 ( .A1(n1055), .A2(mem[965]), .B1(n1044), .B2(mem[805]), .ZN(
        n1407) );
  AOI22_X1 U733 ( .A1(n1039), .A2(mem[933]), .B1(n2705), .B2(mem[741]), .ZN(
        n1406) );
  AOI22_X1 U734 ( .A1(n2668), .A2(mem[613]), .B1(n2869), .B2(mem[901]), .ZN(
        n1405) );
  AOI22_X1 U735 ( .A1(n2062), .A2(mem[485]), .B1(n1041), .B2(mem[165]), .ZN(
        n1404) );
  NAND4_X1 U736 ( .A1(n1407), .A2(n1406), .A3(n1405), .A4(n1404), .ZN(n1422)
         );
  AOI22_X1 U737 ( .A1(n1047), .A2(mem[69]), .B1(n1408), .B2(mem[101]), .ZN(
        n1413) );
  AOI22_X1 U738 ( .A1(n1042), .A2(mem[229]), .B1(n1054), .B2(mem[325]), .ZN(
        n1412) );
  AOI22_X1 U739 ( .A1(n2750), .A2(mem[517]), .B1(n1046), .B2(mem[453]), .ZN(
        n1411) );
  AOI22_X1 U740 ( .A1(n3015), .A2(mem[709]), .B1(n1053), .B2(mem[421]), .ZN(
        n1410) );
  NAND4_X1 U741 ( .A1(n1413), .A2(n1412), .A3(n1411), .A4(n1410), .ZN(n1421)
         );
  AOI22_X1 U742 ( .A1(n1040), .A2(mem[197]), .B1(n2578), .B2(mem[645]), .ZN(
        n1419) );
  AOI22_X1 U743 ( .A1(n3001), .A2(mem[37]), .B1(n1045), .B2(mem[5]), .ZN(n1418) );
  AOI22_X1 U744 ( .A1(n1033), .A2(mem[389]), .B1(n1052), .B2(mem[677]), .ZN(
        n1417) );
  AOI22_X1 U745 ( .A1(n1048), .A2(mem[773]), .B1(n1056), .B2(mem[869]), .ZN(
        n1416) );
  NAND4_X1 U746 ( .A1(n1419), .A2(n1418), .A3(n1417), .A4(n1416), .ZN(n1420)
         );
  OR4_X1 U747 ( .A1(n1423), .A2(n1422), .A3(n1421), .A4(n1420), .ZN(
        rdata_c_o[5]) );
  AOI22_X1 U748 ( .A1(n1053), .A2(mem[427]), .B1(n3010), .B2(mem[555]), .ZN(
        n1428) );
  AOI22_X1 U749 ( .A1(n1055), .A2(mem[971]), .B1(n1054), .B2(mem[331]), .ZN(
        n1427) );
  AOI22_X1 U750 ( .A1(n1050), .A2(mem[843]), .B1(n1402), .B2(mem[939]), .ZN(
        n1426) );
  NAND2_X1 U751 ( .A1(n2874), .A2(mem[363]), .ZN(n1425) );
  NAND4_X1 U752 ( .A1(n1428), .A2(n1427), .A3(n1426), .A4(n1425), .ZN(n1447)
         );
  AOI22_X1 U753 ( .A1(n1033), .A2(mem[395]), .B1(n1040), .B2(mem[203]), .ZN(
        n1435) );
  AOI22_X1 U754 ( .A1(n1752), .A2(mem[587]), .B1(n1056), .B2(mem[875]), .ZN(
        n1434) );
  AOI22_X1 U755 ( .A1(n1452), .A2(mem[715]), .B1(n1047), .B2(mem[75]), .ZN(
        n1433) );
  AOI22_X1 U756 ( .A1(n1041), .A2(mem[171]), .B1(n1052), .B2(mem[683]), .ZN(
        n1432) );
  NAND4_X1 U757 ( .A1(n1435), .A2(n1434), .A3(n1433), .A4(n1432), .ZN(n1446)
         );
  AOI22_X1 U758 ( .A1(n2705), .A2(mem[747]), .B1(n1046), .B2(mem[459]), .ZN(
        n1439) );
  AOI22_X1 U759 ( .A1(n2750), .A2(mem[523]), .B1(n1043), .B2(mem[107]), .ZN(
        n1438) );
  AOI22_X1 U760 ( .A1(n1740), .A2(mem[491]), .B1(n3001), .B2(mem[43]), .ZN(
        n1437) );
  AOI22_X1 U761 ( .A1(n1042), .A2(mem[235]), .B1(n2578), .B2(mem[651]), .ZN(
        n1436) );
  NAND4_X1 U762 ( .A1(n1439), .A2(n1438), .A3(n1437), .A4(n1436), .ZN(n1445)
         );
  AOI22_X1 U763 ( .A1(n1045), .A2(mem[11]), .B1(n1044), .B2(mem[811]), .ZN(
        n1443) );
  AOI22_X1 U764 ( .A1(n2668), .A2(mem[619]), .B1(n1051), .B2(mem[139]), .ZN(
        n1442) );
  AOI22_X1 U765 ( .A1(n2869), .A2(mem[907]), .B1(n1048), .B2(mem[779]), .ZN(
        n1441) );
  AOI22_X1 U766 ( .A1(n3016), .A2(mem[299]), .B1(n1049), .B2(mem[267]), .ZN(
        n1440) );
  NAND4_X1 U767 ( .A1(n1443), .A2(n1442), .A3(n1441), .A4(n1440), .ZN(n1444)
         );
  OR4_X1 U768 ( .A1(n1447), .A2(n1446), .A3(n1445), .A4(n1444), .ZN(
        rdata_c_o[11]) );
  AOI22_X1 U769 ( .A1(n2433), .A2(mem[578]), .B1(n2578), .B2(mem[642]), .ZN(
        n1451) );
  AOI22_X1 U770 ( .A1(n1414), .A2(mem[34]), .B1(n3010), .B2(mem[546]), .ZN(
        n1450) );
  AOI22_X1 U771 ( .A1(n1045), .A2(mem[2]), .B1(n1403), .B2(mem[898]), .ZN(
        n1449) );
  NAND2_X1 U772 ( .A1(n2874), .A2(mem[354]), .ZN(n1448) );
  NAND4_X1 U773 ( .A1(n1451), .A2(n1450), .A3(n1449), .A4(n1448), .ZN(n1469)
         );
  AOI22_X1 U774 ( .A1(n1053), .A2(mem[418]), .B1(n2750), .B2(mem[514]), .ZN(
        n1456) );
  AOI22_X1 U775 ( .A1(n3016), .A2(mem[290]), .B1(n1056), .B2(mem[866]), .ZN(
        n1455) );
  AOI22_X1 U776 ( .A1(n1042), .A2(mem[226]), .B1(n1452), .B2(mem[706]), .ZN(
        n1454) );
  AOI22_X1 U777 ( .A1(n2668), .A2(mem[610]), .B1(n1049), .B2(mem[258]), .ZN(
        n1453) );
  NAND4_X1 U778 ( .A1(n1456), .A2(n1455), .A3(n1454), .A4(n1453), .ZN(n1468)
         );
  AOI22_X1 U779 ( .A1(n1033), .A2(mem[386]), .B1(n1044), .B2(mem[802]), .ZN(
        n1460) );
  AOI22_X1 U780 ( .A1(n1046), .A2(mem[450]), .B1(n1051), .B2(mem[130]), .ZN(
        n1459) );
  AOI22_X1 U781 ( .A1(n1041), .A2(mem[162]), .B1(n1054), .B2(mem[322]), .ZN(
        n1458) );
  AOI22_X1 U782 ( .A1(n1516), .A2(mem[834]), .B1(n1048), .B2(mem[770]), .ZN(
        n1457) );
  NAND4_X1 U783 ( .A1(n1460), .A2(n1459), .A3(n1458), .A4(n1457), .ZN(n1467)
         );
  AOI22_X1 U784 ( .A1(n1052), .A2(mem[674]), .B1(n1408), .B2(mem[98]), .ZN(
        n1465) );
  AOI22_X1 U785 ( .A1(n2062), .A2(mem[482]), .B1(n1750), .B2(mem[962]), .ZN(
        n1464) );
  AOI22_X1 U786 ( .A1(n1040), .A2(mem[194]), .B1(n1047), .B2(mem[66]), .ZN(
        n1463) );
  AOI22_X1 U787 ( .A1(n1039), .A2(mem[930]), .B1(n1461), .B2(mem[738]), .ZN(
        n1462) );
  NAND4_X1 U788 ( .A1(n1465), .A2(n1464), .A3(n1463), .A4(n1462), .ZN(n1466)
         );
  OR4_X1 U789 ( .A1(n1469), .A2(n1468), .A3(n1467), .A4(n1466), .ZN(
        rdata_c_o[2]) );
  AOI22_X1 U790 ( .A1(n1740), .A2(mem[486]), .B1(n2578), .B2(mem[646]), .ZN(
        n1473) );
  AOI22_X1 U791 ( .A1(n1055), .A2(mem[966]), .B1(n2705), .B2(mem[742]), .ZN(
        n1472) );
  AOI22_X1 U792 ( .A1(n2869), .A2(mem[902]), .B1(n1053), .B2(mem[422]), .ZN(
        n1471) );
  NAND2_X1 U793 ( .A1(n3010), .A2(mem[550]), .ZN(n1470) );
  NAND4_X1 U794 ( .A1(n1473), .A2(n1472), .A3(n1471), .A4(n1470), .ZN(n1490)
         );
  AOI22_X1 U795 ( .A1(n1752), .A2(mem[582]), .B1(n1054), .B2(mem[326]), .ZN(
        n1478) );
  AOI22_X1 U796 ( .A1(n1040), .A2(mem[198]), .B1(n1048), .B2(mem[774]), .ZN(
        n1477) );
  AOI22_X1 U797 ( .A1(n1414), .A2(mem[38]), .B1(n1395), .B2(mem[294]), .ZN(
        n1476) );
  AOI22_X1 U798 ( .A1(n1045), .A2(mem[6]), .B1(n2750), .B2(mem[518]), .ZN(
        n1475) );
  NAND4_X1 U799 ( .A1(n1478), .A2(n1477), .A3(n1476), .A4(n1475), .ZN(n1489)
         );
  AOI22_X1 U800 ( .A1(n1452), .A2(mem[710]), .B1(n1047), .B2(mem[70]), .ZN(
        n1482) );
  AOI22_X1 U801 ( .A1(n1033), .A2(mem[390]), .B1(n1052), .B2(mem[678]), .ZN(
        n1481) );
  AOI22_X1 U802 ( .A1(n1044), .A2(mem[806]), .B1(n1051), .B2(mem[134]), .ZN(
        n1480) );
  AOI22_X1 U803 ( .A1(n1516), .A2(mem[838]), .B1(n1424), .B2(mem[358]), .ZN(
        n1479) );
  NAND4_X1 U804 ( .A1(n1482), .A2(n1481), .A3(n1480), .A4(n1479), .ZN(n1488)
         );
  AOI22_X1 U805 ( .A1(n1041), .A2(mem[166]), .B1(n1042), .B2(mem[230]), .ZN(
        n1486) );
  AOI22_X1 U806 ( .A1(n1039), .A2(mem[934]), .B1(n1408), .B2(mem[102]), .ZN(
        n1485) );
  AOI22_X1 U807 ( .A1(n2668), .A2(mem[614]), .B1(n1049), .B2(mem[262]), .ZN(
        n1484) );
  AOI22_X1 U808 ( .A1(n1046), .A2(mem[454]), .B1(n1056), .B2(mem[870]), .ZN(
        n1483) );
  NAND4_X1 U809 ( .A1(n1486), .A2(n1485), .A3(n1484), .A4(n1483), .ZN(n1487)
         );
  OR4_X1 U810 ( .A1(n1490), .A2(n1489), .A3(n1488), .A4(n1487), .ZN(
        rdata_c_o[6]) );
  AOI22_X1 U811 ( .A1(n2668), .A2(mem[612]), .B1(n1402), .B2(mem[932]), .ZN(
        n1494) );
  AOI22_X1 U812 ( .A1(n1516), .A2(mem[836]), .B1(n1044), .B2(mem[804]), .ZN(
        n1493) );
  AOI22_X1 U813 ( .A1(n1042), .A2(mem[228]), .B1(n1046), .B2(mem[452]), .ZN(
        n1492) );
  NAND2_X1 U814 ( .A1(n1055), .A2(mem[964]), .ZN(n1491) );
  NAND4_X1 U815 ( .A1(n1494), .A2(n1493), .A3(n1492), .A4(n1491), .ZN(n1510)
         );
  AOI22_X1 U816 ( .A1(n1424), .A2(mem[356]), .B1(n1403), .B2(mem[900]), .ZN(
        n1498) );
  AOI22_X1 U817 ( .A1(n3016), .A2(mem[292]), .B1(n2578), .B2(mem[644]), .ZN(
        n1497) );
  AOI22_X1 U818 ( .A1(n1053), .A2(mem[420]), .B1(n1056), .B2(mem[868]), .ZN(
        n1496) );
  AOI22_X1 U819 ( .A1(n1045), .A2(mem[4]), .B1(n1051), .B2(mem[132]), .ZN(
        n1495) );
  NAND4_X1 U820 ( .A1(n1498), .A2(n1497), .A3(n1496), .A4(n1495), .ZN(n1509)
         );
  AOI22_X1 U821 ( .A1(n2705), .A2(mem[740]), .B1(n2750), .B2(mem[516]), .ZN(
        n1502) );
  AOI22_X1 U822 ( .A1(n1052), .A2(mem[676]), .B1(n3010), .B2(mem[548]), .ZN(
        n1501) );
  AOI22_X1 U823 ( .A1(n2062), .A2(mem[484]), .B1(n1041), .B2(mem[164]), .ZN(
        n1500) );
  AOI22_X1 U824 ( .A1(n1040), .A2(mem[196]), .B1(n1054), .B2(mem[324]), .ZN(
        n1499) );
  NAND4_X1 U825 ( .A1(n1502), .A2(n1501), .A3(n1500), .A4(n1499), .ZN(n1508)
         );
  AOI22_X1 U826 ( .A1(n1033), .A2(mem[388]), .B1(n1049), .B2(mem[260]), .ZN(
        n1506) );
  AOI22_X1 U827 ( .A1(n1414), .A2(mem[36]), .B1(n1408), .B2(mem[100]), .ZN(
        n1505) );
  AOI22_X1 U828 ( .A1(n2433), .A2(mem[580]), .B1(n1047), .B2(mem[68]), .ZN(
        n1504) );
  AOI22_X1 U829 ( .A1(n1452), .A2(mem[708]), .B1(n1048), .B2(mem[772]), .ZN(
        n1503) );
  NAND4_X1 U830 ( .A1(n1506), .A2(n1505), .A3(n1504), .A4(n1503), .ZN(n1507)
         );
  OR4_X1 U831 ( .A1(n1510), .A2(n1509), .A3(n1508), .A4(n1507), .ZN(
        rdata_c_o[4]) );
  AOI22_X1 U832 ( .A1(n2668), .A2(mem[611]), .B1(n1040), .B2(mem[195]), .ZN(
        n1515) );
  AOI22_X1 U833 ( .A1(n1045), .A2(mem[3]), .B1(n1042), .B2(mem[227]), .ZN(
        n1514) );
  AOI22_X1 U834 ( .A1(n2433), .A2(mem[579]), .B1(n2750), .B2(mem[515]), .ZN(
        n1513) );
  NAND2_X1 U835 ( .A1(n1452), .A2(mem[707]), .ZN(n1512) );
  NAND4_X1 U836 ( .A1(n1515), .A2(n1514), .A3(n1513), .A4(n1512), .ZN(n1533)
         );
  AOI22_X1 U837 ( .A1(n1039), .A2(mem[931]), .B1(n1049), .B2(mem[259]), .ZN(
        n1520) );
  AOI22_X1 U838 ( .A1(n1516), .A2(mem[835]), .B1(n1046), .B2(mem[451]), .ZN(
        n1519) );
  AOI22_X1 U839 ( .A1(n1044), .A2(mem[803]), .B1(n3010), .B2(mem[547]), .ZN(
        n1518) );
  AOI22_X1 U840 ( .A1(n2705), .A2(mem[739]), .B1(n1408), .B2(mem[99]), .ZN(
        n1517) );
  NAND4_X1 U841 ( .A1(n1520), .A2(n1519), .A3(n1518), .A4(n1517), .ZN(n1532)
         );
  AOI22_X1 U842 ( .A1(n2062), .A2(mem[483]), .B1(n1395), .B2(mem[291]), .ZN(
        n1525) );
  AOI22_X1 U843 ( .A1(n1414), .A2(mem[35]), .B1(n1033), .B2(mem[387]), .ZN(
        n1524) );
  AOI22_X1 U844 ( .A1(n1055), .A2(mem[963]), .B1(n2869), .B2(mem[899]), .ZN(
        n1523) );
  AOI22_X1 U845 ( .A1(n1424), .A2(mem[355]), .B1(n1053), .B2(mem[419]), .ZN(
        n1522) );
  NAND4_X1 U846 ( .A1(n1525), .A2(n1524), .A3(n1523), .A4(n1522), .ZN(n1531)
         );
  AOI22_X1 U847 ( .A1(n1041), .A2(mem[163]), .B1(n1051), .B2(mem[131]), .ZN(
        n1529) );
  AOI22_X1 U848 ( .A1(n1047), .A2(mem[67]), .B1(n1056), .B2(mem[867]), .ZN(
        n1528) );
  AOI22_X1 U849 ( .A1(n1052), .A2(mem[675]), .B1(n1048), .B2(mem[771]), .ZN(
        n1527) );
  AOI22_X1 U850 ( .A1(n1054), .A2(mem[323]), .B1(n2578), .B2(mem[643]), .ZN(
        n1526) );
  NAND4_X1 U851 ( .A1(n1529), .A2(n1528), .A3(n1527), .A4(n1526), .ZN(n1530)
         );
  OR4_X1 U852 ( .A1(n1533), .A2(n1532), .A3(n1531), .A4(n1530), .ZN(
        rdata_c_o[3]) );
  INV_X1 U853 ( .A(wdata_b_i[3]), .ZN(n4414) );
  INV_X1 U855 ( .A(waddr_b_i[0]), .ZN(n1534) );
  NAND2_X1 U856 ( .A1(we_b_i), .A2(n1534), .ZN(n1560) );
  INV_X1 U857 ( .A(waddr_b_i[3]), .ZN(n2468) );
  NOR2_X1 U859 ( .A1(n2532), .A2(n2527), .ZN(n3771) );
  INV_X1 U860 ( .A(n3771), .ZN(n1565) );
  INV_X1 U861 ( .A(waddr_a_i[4]), .ZN(n1536) );
  NOR2_X1 U862 ( .A1(n1536), .A2(waddr_a_i[3]), .ZN(n1554) );
  NAND2_X1 U863 ( .A1(n1554), .A2(n2533), .ZN(n1596) );
  NOR2_X1 U864 ( .A1(n1565), .A2(n1596), .ZN(n1539) );
  INV_X1 U865 ( .A(n1539), .ZN(n1537) );
  NOR2_X1 U870 ( .A1(waddr_b_i[1]), .A2(waddr_b_i[3]), .ZN(n2478) );
  NOR2_X1 U872 ( .A1(n2532), .A2(waddr_a_i[1]), .ZN(n3848) );
  INV_X1 U873 ( .A(n3848), .ZN(n1603) );
  NOR2_X1 U874 ( .A1(n1603), .A2(n1596), .ZN(n1543) );
  INV_X1 U875 ( .A(n1543), .ZN(n1541) );
  AND2_X1 U880 ( .A1(n3770), .A2(n3768), .ZN(n2259) );
  INV_X1 U881 ( .A(n2259), .ZN(n1585) );
  INV_X1 U883 ( .A(waddr_a_i[3]), .ZN(n1545) );
  NOR2_X1 U884 ( .A1(n1545), .A2(waddr_a_i[4]), .ZN(n2262) );
  NAND2_X1 U885 ( .A1(n2262), .A2(n2533), .ZN(n1602) );
  NOR2_X1 U886 ( .A1(n1565), .A2(n1602), .ZN(n1548) );
  INV_X1 U887 ( .A(n1548), .ZN(n1546) );
  NOR2_X1 U892 ( .A1(n2468), .A2(waddr_b_i[1]), .ZN(n3845) );
  NAND2_X1 U893 ( .A1(waddr_b_i[0]), .A2(we_b_i), .ZN(n1614) );
  OR2_X1 U894 ( .A1(n1614), .A2(waddr_b_i[2]), .ZN(n2479) );
  NOR2_X1 U896 ( .A1(n1602), .A2(n2480), .ZN(n1551) );
  INV_X1 U897 ( .A(n1551), .ZN(n1550) );
  INV_X1 U903 ( .A(waddr_b_i[2]), .ZN(n1559) );
  NAND2_X1 U905 ( .A1(n1554), .A2(waddr_a_i[2]), .ZN(n1609) );
  NOR2_X1 U906 ( .A1(n1609), .A2(n2480), .ZN(n1556) );
  INV_X1 U907 ( .A(n1556), .ZN(n1555) );
  OR2_X1 U912 ( .A1(n1560), .A2(n1559), .ZN(n2547) );
  NOR2_X1 U914 ( .A1(n1603), .A2(n1609), .ZN(n1563) );
  INV_X1 U915 ( .A(n1563), .ZN(n1561) );
  NOR2_X1 U921 ( .A1(n1565), .A2(n1609), .ZN(n1568) );
  INV_X1 U922 ( .A(n1568), .ZN(n1566) );
  NOR3_X1 U928 ( .A1(waddr_a_i[1]), .A2(waddr_a_i[4]), .A3(n1586), .ZN(n1570)
         );
  NAND3_X1 U929 ( .A1(waddr_a_i[2]), .A2(waddr_a_i[3]), .A3(n1570), .ZN(n1571)
         );
  NOR2_X1 U936 ( .A1(n2532), .A2(n2533), .ZN(n2549) );
  INV_X1 U937 ( .A(n2549), .ZN(n1576) );
  INV_X1 U938 ( .A(n2262), .ZN(n1575) );
  NOR3_X1 U939 ( .A1(n1576), .A2(waddr_a_i[1]), .A3(n1575), .ZN(n1579) );
  INV_X1 U940 ( .A(n1579), .ZN(n1577) );
  AND3_X1 U946 ( .A1(n2549), .A2(waddr_a_i[1]), .A3(n2262), .ZN(n1582) );
  INV_X1 U947 ( .A(n1582), .ZN(n1581) );
  INV_X1 U953 ( .A(n1586), .ZN(n2473) );
  AND2_X1 U954 ( .A1(waddr_a_i[1]), .A2(n2473), .ZN(n2261) );
  INV_X1 U955 ( .A(n2261), .ZN(n1615) );
  OR2_X1 U956 ( .A1(n1602), .A2(n1615), .ZN(n1587) );
  NOR2_X1 U963 ( .A1(n1596), .A2(n2480), .ZN(n1593) );
  INV_X1 U964 ( .A(n1593), .ZN(n1592) );
  NOR2_X1 U970 ( .A1(n1596), .A2(n1615), .ZN(n1598) );
  INV_X1 U971 ( .A(n1598), .ZN(n1597) );
  NOR2_X1 U977 ( .A1(n1603), .A2(n1602), .ZN(n1606) );
  INV_X1 U978 ( .A(n1606), .ZN(n1604) );
  NOR2_X1 U984 ( .A1(n1609), .A2(n1615), .ZN(n1611) );
  INV_X1 U985 ( .A(n1611), .ZN(n1610) );
  OR2_X1 U990 ( .A1(n3768), .A2(n1614), .ZN(n1620) );
  NOR2_X1 U991 ( .A1(waddr_b_i[2]), .A2(n1620), .ZN(n1643) );
  NAND2_X1 U993 ( .A1(waddr_a_i[3]), .A2(waddr_a_i[4]), .ZN(n1622) );
  OR2_X1 U994 ( .A1(n1622), .A2(waddr_a_i[2]), .ZN(n1644) );
  NOR2_X1 U995 ( .A1(n1644), .A2(n1615), .ZN(n1618) );
  INV_X1 U996 ( .A(n1618), .ZN(n1616) );
  INV_X1 U1001 ( .A(n1620), .ZN(n1621) );
  AND2_X1 U1002 ( .A1(waddr_b_i[2]), .A2(n1621), .ZN(n1636) );
  NAND2_X1 U1004 ( .A1(n1637), .A2(n2261), .ZN(n1623) );
  INV_X1 U1006 ( .A(n1623), .ZN(n1625) );
  NOR2_X1 U1010 ( .A1(n2547), .A2(n3768), .ZN(n1631) );
  NAND2_X1 U1012 ( .A1(n3771), .A2(n1637), .ZN(n1627) );
  NAND2_X1 U1019 ( .A1(n3848), .A2(n1637), .ZN(n1632) );
  INV_X1 U1026 ( .A(n1637), .ZN(n1638) );
  NOR2_X1 U1027 ( .A1(n1638), .A2(n2480), .ZN(n1641) );
  INV_X1 U1028 ( .A(n1641), .ZN(n1639) );
  INV_X1 U1034 ( .A(n1644), .ZN(n3847) );
  INV_X1 U1035 ( .A(n2480), .ZN(n1645) );
  NAND2_X1 U1036 ( .A1(n3847), .A2(n1645), .ZN(n1646) );
  INV_X1 U1038 ( .A(n1646), .ZN(n1648) );
  AOI22_X1 U1075 ( .A1(n2852), .A2(mem[796]), .B1(n2841), .B2(mem[732]), .ZN(
        n1668) );
  AOI22_X1 U1076 ( .A1(n2980), .A2(mem[764]), .B1(n2786), .B2(mem[572]), .ZN(
        n1667) );
  AOI22_X1 U1077 ( .A1(n2978), .A2(mem[284]), .B1(n2860), .B2(mem[188]), .ZN(
        n1666) );
  NAND2_X1 U1078 ( .A1(n2963), .A2(mem[956]), .ZN(n1665) );
  NAND4_X1 U1079 ( .A1(n1668), .A2(n1667), .A3(n1666), .A4(n1665), .ZN(n1684)
         );
  AOI22_X1 U1080 ( .A1(n2853), .A2(mem[892]), .B1(n2974), .B2(mem[124]), .ZN(
        n1672) );
  AOI22_X1 U1081 ( .A1(n2969), .A2(mem[700]), .B1(n2965), .B2(mem[508]), .ZN(
        n1671) );
  AOI22_X1 U1082 ( .A1(n2957), .A2(mem[252]), .B1(n2776), .B2(mem[220]), .ZN(
        n1670) );
  AOI22_X1 U1083 ( .A1(n2833), .A2(mem[476]), .B1(n2979), .B2(mem[28]), .ZN(
        n1669) );
  NAND4_X1 U1084 ( .A1(n1672), .A2(n1671), .A3(n1670), .A4(n1669), .ZN(n1683)
         );
  AOI22_X1 U1085 ( .A1(n2951), .A2(mem[156]), .B1(n2988), .B2(mem[540]), .ZN(
        n1676) );
  AOI22_X1 U1086 ( .A1(n2832), .A2(mem[444]), .B1(n2842), .B2(mem[380]), .ZN(
        n1675) );
  AOI22_X1 U1087 ( .A1(n2770), .A2(mem[636]), .B1(n2765), .B2(mem[604]), .ZN(
        n1674) );
  AOI22_X1 U1088 ( .A1(n2990), .A2(mem[60]), .B1(n2639), .B2(mem[860]), .ZN(
        n1673) );
  NAND4_X1 U1089 ( .A1(n1676), .A2(n1675), .A3(n1674), .A4(n1673), .ZN(n1682)
         );
  AOI22_X1 U1090 ( .A1(n2967), .A2(mem[668]), .B1(n2987), .B2(mem[412]), .ZN(
        n1680) );
  AOI22_X1 U1091 ( .A1(n2798), .A2(mem[92]), .B1(n2976), .B2(mem[316]), .ZN(
        n1679) );
  AOI22_X1 U1092 ( .A1(n2791), .A2(mem[988]), .B1(n2840), .B2(mem[828]), .ZN(
        n1678) );
  AOI22_X1 U1093 ( .A1(n2968), .A2(mem[924]), .B1(n2985), .B2(mem[348]), .ZN(
        n1677) );
  NAND4_X1 U1094 ( .A1(n1680), .A2(n1679), .A3(n1678), .A4(n1677), .ZN(n1681)
         );
  OR4_X1 U1095 ( .A1(n1684), .A2(n1683), .A3(n1682), .A4(n1681), .ZN(
        rdata_b_o[28]) );
  INV_X1 U1096 ( .A(raddr_a_i[3]), .ZN(n1685) );
  OR2_X1 U1097 ( .A1(n1685), .A2(raddr_a_i[4]), .ZN(n1686) );
  INV_X1 U1098 ( .A(raddr_a_i[2]), .ZN(n1719) );
  NOR2_X1 U1099 ( .A1(n1686), .A2(n1719), .ZN(n1704) );
  NOR2_X1 U1100 ( .A1(raddr_a_i[1]), .A2(raddr_a_i[0]), .ZN(n1710) );
  NOR2_X1 U1101 ( .A1(n1686), .A2(n997), .ZN(n1705) );
  BUF_X1 U1104 ( .A(n2162), .Z(n3577) );
  AOI22_X1 U1105 ( .A1(mem[380]), .A2(n1023), .B1(n3577), .B2(mem[316]), .ZN(
        n1695) );
  INV_X1 U1106 ( .A(raddr_a_i[4]), .ZN(n1688) );
  NOR2_X1 U1108 ( .A1(n1696), .A2(n997), .ZN(n1718) );
  OR2_X1 U1109 ( .A1(raddr_a_i[4]), .A2(raddr_a_i[3]), .ZN(n1697) );
  NOR2_X1 U1110 ( .A1(n1697), .A2(raddr_a_i[2]), .ZN(n1691) );
  AOI22_X1 U1111 ( .A1(n1092), .A2(mem[508]), .B1(mem[60]), .B2(n4730), .ZN(
        n1694) );
  INV_X1 U1112 ( .A(n1724), .ZN(n1689) );
  AOI22_X1 U1116 ( .A1(mem[92]), .A2(n3512), .B1(n3578), .B2(mem[28]), .ZN(
        n1693) );
  NAND2_X1 U1117 ( .A1(raddr_a_i[4]), .A2(raddr_a_i[3]), .ZN(n1720) );
  OR2_X1 U1118 ( .A1(n1720), .A2(raddr_a_i[2]), .ZN(n1725) );
  INV_X1 U1119 ( .A(n1717), .ZN(n1722) );
  NOR2_X1 U1120 ( .A1(n1725), .A2(n1722), .ZN(n1811) );
  NAND2_X1 U1121 ( .A1(n1027), .A2(mem[796]), .ZN(n1692) );
  NAND4_X1 U1122 ( .A1(n1695), .A2(n1694), .A3(n1693), .A4(n1692), .ZN(n1733)
         );
  AND2_X1 U1123 ( .A1(n1706), .A2(n1708), .ZN(n3188) );
  AND2_X1 U1124 ( .A1(n1717), .A2(n1704), .ZN(n2153) );
  BUF_X1 U1125 ( .A(n2153), .Z(n3585) );
  AOI22_X1 U1126 ( .A1(mem[700]), .A2(n1070), .B1(n3585), .B2(mem[412]), .ZN(
        n1702) );
  NOR2_X1 U1127 ( .A1(n1697), .A2(n1719), .ZN(n1698) );
  INV_X1 U1128 ( .A(n1698), .ZN(n1712) );
  NOR2_X1 U1129 ( .A1(n1712), .A2(n1724), .ZN(n2156) );
  AOI22_X1 U1130 ( .A1(n1018), .A2(mem[220]), .B1(mem[124]), .B2(n1029), .ZN(
        n1701) );
  AND2_X1 U1131 ( .A1(n1710), .A2(n1706), .ZN(n3189) );
  AND2_X1 U1132 ( .A1(n1718), .A2(n1708), .ZN(n2154) );
  BUF_X1 U1133 ( .A(n2154), .Z(n3586) );
  AOI22_X1 U1134 ( .A1(mem[636]), .A2(n1071), .B1(n3586), .B2(mem[572]), .ZN(
        n1700) );
  AND2_X1 U1135 ( .A1(n1706), .A2(n1717), .ZN(n3061) );
  AND2_X1 U1136 ( .A1(n1698), .A2(n1708), .ZN(n3114) );
  AOI22_X1 U1137 ( .A1(n3587), .A2(mem[668]), .B1(mem[188]), .B2(n1072), .ZN(
        n1699) );
  NAND4_X1 U1138 ( .A1(n1702), .A2(n1701), .A3(n1700), .A4(n1699), .ZN(n1732)
         );
  INV_X1 U1139 ( .A(n1718), .ZN(n1703) );
  NOR2_X1 U1140 ( .A1(n1703), .A2(n1724), .ZN(n3078) );
  INV_X1 U1141 ( .A(n1704), .ZN(n1709) );
  NOR2_X1 U1142 ( .A1(n1709), .A2(n1724), .ZN(n3207) );
  AOI22_X1 U1143 ( .A1(mem[604]), .A2(n1016), .B1(n994), .B2(mem[476]), .ZN(
        n1716) );
  INV_X1 U1144 ( .A(n1705), .ZN(n1711) );
  NOR2_X1 U1145 ( .A1(n1711), .A2(n1724), .ZN(n3075) );
  NOR2_X1 U1146 ( .A1(n1711), .A2(n1722), .ZN(n3176) );
  AOI22_X1 U1147 ( .A1(mem[348]), .A2(n1007), .B1(n1084), .B2(mem[284]), .ZN(
        n1715) );
  INV_X1 U1148 ( .A(n1706), .ZN(n1707) );
  NOR2_X1 U1149 ( .A1(n1707), .A2(n1724), .ZN(n2146) );
  AOI22_X1 U1150 ( .A1(mem[732]), .A2(n1080), .B1(n1013), .B2(mem[444]), .ZN(
        n1714) );
  INV_X1 U1151 ( .A(n1710), .ZN(n1721) );
  NOR2_X1 U1152 ( .A1(n1711), .A2(n1721), .ZN(n2148) );
  NOR2_X1 U1153 ( .A1(n1712), .A2(n1722), .ZN(n3102) );
  AOI22_X1 U1154 ( .A1(n1010), .A2(mem[252]), .B1(mem[156]), .B2(n1022), .ZN(
        n1713) );
  NAND4_X1 U1155 ( .A1(n1716), .A2(n1715), .A3(n1714), .A4(n1713), .ZN(n1731)
         );
  AND2_X1 U1156 ( .A1(n1717), .A2(n1718), .ZN(n3194) );
  NOR2_X1 U1157 ( .A1(n1723), .A2(n1095), .ZN(n3040) );
  AOI22_X1 U1158 ( .A1(n1068), .A2(mem[540]), .B1(mem[956]), .B2(n3592), .ZN(
        n1729) );
  NOR2_X1 U1159 ( .A1(n1723), .A2(n1724), .ZN(n2169) );
  BUF_X1 U1160 ( .A(n2169), .Z(n3564) );
  NOR2_X1 U1161 ( .A1(n1725), .A2(n1721), .ZN(n3195) );
  AOI22_X1 U1162 ( .A1(mem[988]), .A2(n3564), .B1(n1087), .B2(mem[764]), .ZN(
        n1728) );
  NOR2_X1 U1163 ( .A1(n1723), .A2(n1721), .ZN(n3092) );
  NOR2_X1 U1164 ( .A1(n1725), .A2(n1095), .ZN(n3196) );
  AOI22_X1 U1165 ( .A1(mem[892]), .A2(n3593), .B1(n1069), .B2(mem[828]), .ZN(
        n1727) );
  NOR2_X1 U1166 ( .A1(n1722), .A2(n1723), .ZN(n2170) );
  NOR2_X1 U1167 ( .A1(n1725), .A2(n1724), .ZN(n3222) );
  AOI22_X1 U1168 ( .A1(mem[924]), .A2(n3594), .B1(n1090), .B2(mem[860]), .ZN(
        n1726) );
  NAND4_X1 U1169 ( .A1(n1729), .A2(n1728), .A3(n1727), .A4(n1726), .ZN(n1730)
         );
  OR4_X1 U1170 ( .A1(n1733), .A2(n1732), .A3(n1731), .A4(n1730), .ZN(
        rdata_a_o[28]) );
  AOI22_X1 U1171 ( .A1(n1050), .A2(mem[860]), .B1(n1046), .B2(mem[476]), .ZN(
        n1737) );
  AOI22_X1 U1172 ( .A1(n2869), .A2(mem[924]), .B1(n1043), .B2(mem[124]), .ZN(
        n1736) );
  AOI22_X1 U1173 ( .A1(n1044), .A2(mem[828]), .B1(n3010), .B2(mem[572]), .ZN(
        n1735) );
  NAND2_X1 U1174 ( .A1(n1040), .A2(mem[220]), .ZN(n1734) );
  NAND4_X1 U1175 ( .A1(n1737), .A2(n1736), .A3(n1735), .A4(n1734), .ZN(n1760)
         );
  AOI22_X1 U1176 ( .A1(n1041), .A2(mem[188]), .B1(n1049), .B2(mem[284]), .ZN(
        n1744) );
  AOI22_X1 U1177 ( .A1(n1054), .A2(mem[348]), .B1(n1048), .B2(mem[796]), .ZN(
        n1743) );
  AOI22_X1 U1178 ( .A1(n1740), .A2(mem[508]), .B1(n1056), .B2(mem[892]), .ZN(
        n1742) );
  AOI22_X1 U1179 ( .A1(n3001), .A2(mem[60]), .B1(n3015), .B2(mem[732]), .ZN(
        n1741) );
  NAND4_X1 U1180 ( .A1(n1744), .A2(n1743), .A3(n1742), .A4(n1741), .ZN(n1759)
         );
  AOI22_X1 U1181 ( .A1(n1745), .A2(mem[636]), .B1(n1047), .B2(mem[92]), .ZN(
        n1749) );
  AOI22_X1 U1182 ( .A1(n1053), .A2(mem[444]), .B1(n2578), .B2(mem[668]), .ZN(
        n1748) );
  AOI22_X1 U1183 ( .A1(n2874), .A2(mem[380]), .B1(n1052), .B2(mem[700]), .ZN(
        n1747) );
  AOI22_X1 U1184 ( .A1(n1039), .A2(mem[956]), .B1(n1461), .B2(mem[764]), .ZN(
        n1746) );
  NAND4_X1 U1185 ( .A1(n1749), .A2(n1748), .A3(n1747), .A4(n1746), .ZN(n1758)
         );
  AOI22_X1 U1186 ( .A1(n1055), .A2(mem[988]), .B1(n2750), .B2(mem[540]), .ZN(
        n1756) );
  AOI22_X1 U1187 ( .A1(n3016), .A2(mem[316]), .B1(n1042), .B2(mem[252]), .ZN(
        n1755) );
  AOI22_X1 U1188 ( .A1(n1045), .A2(mem[28]), .B1(n1051), .B2(mem[156]), .ZN(
        n1754) );
  AOI22_X1 U1189 ( .A1(n2433), .A2(mem[604]), .B1(n1033), .B2(mem[412]), .ZN(
        n1753) );
  NAND4_X1 U1190 ( .A1(n1756), .A2(n1755), .A3(n1754), .A4(n1753), .ZN(n1757)
         );
  OR4_X1 U1191 ( .A1(n1760), .A2(n1759), .A3(n1758), .A4(n1757), .ZN(
        rdata_c_o[28]) );
  AOI22_X1 U1222 ( .A1(n1055), .A2(mem[990]), .B1(n1452), .B2(mem[734]), .ZN(
        n1780) );
  AOI22_X1 U1223 ( .A1(n1050), .A2(mem[862]), .B1(n1046), .B2(mem[478]), .ZN(
        n1779) );
  AOI22_X1 U1224 ( .A1(n3001), .A2(mem[62]), .B1(n1047), .B2(mem[94]), .ZN(
        n1778) );
  NAND2_X1 U1225 ( .A1(n1056), .A2(mem[894]), .ZN(n1777) );
  NAND4_X1 U1226 ( .A1(n1780), .A2(n1779), .A3(n1778), .A4(n1777), .ZN(n1798)
         );
  AOI22_X1 U1227 ( .A1(n1041), .A2(mem[190]), .B1(n1044), .B2(mem[830]), .ZN(
        n1785) );
  AOI22_X1 U1228 ( .A1(n1042), .A2(mem[254]), .B1(n1053), .B2(mem[446]), .ZN(
        n1784) );
  AOI22_X1 U1229 ( .A1(n1052), .A2(mem[702]), .B1(n3010), .B2(mem[574]), .ZN(
        n1783) );
  AOI22_X1 U1230 ( .A1(n2705), .A2(mem[766]), .B1(n1048), .B2(mem[798]), .ZN(
        n1782) );
  NAND4_X1 U1231 ( .A1(n1785), .A2(n1784), .A3(n1783), .A4(n1782), .ZN(n1797)
         );
  AOI22_X1 U1232 ( .A1(n2433), .A2(mem[606]), .B1(n2750), .B2(mem[542]), .ZN(
        n1790) );
  AOI22_X1 U1233 ( .A1(n1745), .A2(mem[638]), .B1(n1043), .B2(mem[126]), .ZN(
        n1789) );
  AOI22_X1 U1234 ( .A1(n1045), .A2(mem[30]), .B1(n2874), .B2(mem[382]), .ZN(
        n1788) );
  AOI22_X1 U1235 ( .A1(n1033), .A2(mem[414]), .B1(n1040), .B2(mem[222]), .ZN(
        n1787) );
  NAND4_X1 U1236 ( .A1(n1790), .A2(n1789), .A3(n1788), .A4(n1787), .ZN(n1796)
         );
  AOI22_X1 U1237 ( .A1(n2578), .A2(mem[670]), .B1(n1051), .B2(mem[158]), .ZN(
        n1794) );
  AOI22_X1 U1238 ( .A1(n3016), .A2(mem[318]), .B1(n1054), .B2(mem[350]), .ZN(
        n1793) );
  AOI22_X1 U1239 ( .A1(n2062), .A2(mem[510]), .B1(n1403), .B2(mem[926]), .ZN(
        n1792) );
  AOI22_X1 U1240 ( .A1(n1039), .A2(mem[958]), .B1(n1049), .B2(mem[286]), .ZN(
        n1791) );
  NAND4_X1 U1241 ( .A1(n1794), .A2(n1793), .A3(n1792), .A4(n1791), .ZN(n1795)
         );
  OR4_X1 U1242 ( .A1(n1798), .A2(n1797), .A3(n1796), .A4(n1795), .ZN(
        rdata_c_o[30]) );
  AOI22_X1 U1243 ( .A1(mem[382]), .A2(n1023), .B1(n3577), .B2(mem[318]), .ZN(
        n1802) );
  AOI22_X1 U1244 ( .A1(n1092), .A2(mem[510]), .B1(mem[30]), .B2(n3131), .ZN(
        n1801) );
  AOI22_X1 U1245 ( .A1(n1008), .A2(mem[254]), .B1(mem[158]), .B2(n1020), .ZN(
        n1800) );
  NAND2_X1 U1246 ( .A1(n3592), .A2(mem[958]), .ZN(n1799) );
  NAND4_X1 U1247 ( .A1(n1802), .A2(n1801), .A3(n1800), .A4(n1799), .ZN(n1819)
         );
  AOI22_X1 U1248 ( .A1(mem[478]), .A2(n994), .B1(n1085), .B2(mem[286]), .ZN(
        n1806) );
  AOI22_X1 U1249 ( .A1(mem[734]), .A2(n1082), .B1(n1007), .B2(mem[350]), .ZN(
        n1805) );
  AOI22_X1 U1250 ( .A1(n1014), .A2(mem[606]), .B1(n3234), .B2(mem[94]), .ZN(
        n1804) );
  AOI22_X1 U1251 ( .A1(mem[990]), .A2(n1073), .B1(n1086), .B2(mem[766]), .ZN(
        n1803) );
  NAND4_X1 U1252 ( .A1(n1806), .A2(n1805), .A3(n1804), .A4(n1803), .ZN(n1818)
         );
  BUF_X1 U1253 ( .A(n3188), .Z(n3161) );
  AOI22_X1 U1254 ( .A1(mem[702]), .A2(n3161), .B1(n3585), .B2(mem[414]), .ZN(
        n1810) );
  AOI22_X1 U1255 ( .A1(mem[638]), .A2(n3162), .B1(n3586), .B2(mem[574]), .ZN(
        n1809) );
  AOI22_X1 U1256 ( .A1(n1013), .A2(mem[446]), .B1(n4729), .B2(mem[62]), .ZN(
        n1808) );
  AOI22_X1 U1257 ( .A1(mem[126]), .A2(n4736), .B1(n3066), .B2(mem[894]), .ZN(
        n1807) );
  NAND4_X1 U1258 ( .A1(n1810), .A2(n1809), .A3(n1808), .A4(n1807), .ZN(n1817)
         );
  AOI22_X1 U1259 ( .A1(n3587), .A2(mem[670]), .B1(mem[222]), .B2(n1018), .ZN(
        n1815) );
  AOI22_X1 U1260 ( .A1(n3167), .A2(mem[542]), .B1(mem[190]), .B2(n3517), .ZN(
        n1814) );
  BUF_X1 U1261 ( .A(n3196), .Z(n3168) );
  AOI22_X1 U1262 ( .A1(mem[862]), .A2(n1091), .B1(n3168), .B2(mem[830]), .ZN(
        n1813) );
  AOI22_X1 U1263 ( .A1(mem[926]), .A2(n3455), .B1(n1026), .B2(mem[798]), .ZN(
        n1812) );
  NAND4_X1 U1264 ( .A1(n1815), .A2(n1814), .A3(n1813), .A4(n1812), .ZN(n1816)
         );
  OR4_X1 U1265 ( .A1(n1819), .A2(n1818), .A3(n1817), .A4(n1816), .ZN(
        rdata_a_o[30]) );
  AOI22_X1 U1266 ( .A1(n2759), .A2(mem[350]), .B1(n2841), .B2(mem[734]), .ZN(
        n1823) );
  AOI22_X1 U1267 ( .A1(n2853), .A2(mem[894]), .B1(n2835), .B2(mem[542]), .ZN(
        n1822) );
  AOI22_X1 U1268 ( .A1(n2954), .A2(mem[382]), .B1(n2851), .B2(mem[414]), .ZN(
        n1821) );
  NAND2_X1 U1269 ( .A1(n2765), .A2(mem[606]), .ZN(n1820) );
  NAND4_X1 U1270 ( .A1(n1823), .A2(n1822), .A3(n1821), .A4(n1820), .ZN(n1839)
         );
  AOI22_X1 U1271 ( .A1(n2966), .A2(mem[94]), .B1(n2965), .B2(mem[510]), .ZN(
        n1827) );
  AOI22_X1 U1272 ( .A1(n2957), .A2(mem[254]), .B1(n2786), .B2(mem[574]), .ZN(
        n1826) );
  AOI22_X1 U1273 ( .A1(n2977), .A2(mem[222]), .B1(n2951), .B2(mem[158]), .ZN(
        n1825) );
  AOI22_X1 U1274 ( .A1(n2955), .A2(mem[830]), .B1(n1228), .B2(mem[190]), .ZN(
        n1824) );
  NAND4_X1 U1275 ( .A1(n1827), .A2(n1826), .A3(n1825), .A4(n1824), .ZN(n1838)
         );
  AOI22_X1 U1276 ( .A1(n2833), .A2(mem[478]), .B1(n2964), .B2(mem[446]), .ZN(
        n1831) );
  AOI22_X1 U1277 ( .A1(n2764), .A2(mem[766]), .B1(n2989), .B2(mem[990]), .ZN(
        n1830) );
  AOI22_X1 U1278 ( .A1(n2969), .A2(mem[702]), .B1(n2978), .B2(mem[286]), .ZN(
        n1829) );
  AOI22_X1 U1279 ( .A1(n2990), .A2(mem[62]), .B1(n2639), .B2(mem[862]), .ZN(
        n1828) );
  NAND4_X1 U1280 ( .A1(n1831), .A2(n1830), .A3(n1829), .A4(n1828), .ZN(n1837)
         );
  AOI22_X1 U1281 ( .A1(n2797), .A2(mem[958]), .B1(n2975), .B2(mem[798]), .ZN(
        n1835) );
  AOI22_X1 U1282 ( .A1(n2967), .A2(mem[670]), .B1(n2979), .B2(mem[30]), .ZN(
        n1834) );
  AOI22_X1 U1283 ( .A1(n2956), .A2(mem[638]), .B1(n2968), .B2(mem[926]), .ZN(
        n1833) );
  AOI22_X1 U1284 ( .A1(n2974), .A2(mem[126]), .B1(n2858), .B2(mem[318]), .ZN(
        n1832) );
  NAND4_X1 U1285 ( .A1(n1835), .A2(n1834), .A3(n1833), .A4(n1832), .ZN(n1836)
         );
  OR4_X1 U1286 ( .A1(n1839), .A2(n1838), .A3(n1837), .A4(n1836), .ZN(
        rdata_b_o[30]) );
  AOI22_X1 U1287 ( .A1(n2869), .A2(mem[923]), .B1(n1048), .B2(mem[795]), .ZN(
        n1843) );
  AOI22_X1 U1288 ( .A1(n2668), .A2(mem[635]), .B1(n1452), .B2(mem[731]), .ZN(
        n1842) );
  AOI22_X1 U1289 ( .A1(n1033), .A2(mem[411]), .B1(n1054), .B2(mem[347]), .ZN(
        n1841) );
  NAND2_X1 U1290 ( .A1(n2062), .A2(mem[507]), .ZN(n1840) );
  NAND4_X1 U1291 ( .A1(n1843), .A2(n1842), .A3(n1841), .A4(n1840), .ZN(n1859)
         );
  AOI22_X1 U1292 ( .A1(n1055), .A2(mem[987]), .B1(n1041), .B2(mem[187]), .ZN(
        n1847) );
  AOI22_X1 U1293 ( .A1(n1053), .A2(mem[443]), .B1(n1052), .B2(mem[699]), .ZN(
        n1846) );
  AOI22_X1 U1294 ( .A1(n1047), .A2(mem[91]), .B1(n1049), .B2(mem[283]), .ZN(
        n1845) );
  AOI22_X1 U1295 ( .A1(n2578), .A2(mem[667]), .B1(n1461), .B2(mem[763]), .ZN(
        n1844) );
  NAND4_X1 U1296 ( .A1(n1847), .A2(n1846), .A3(n1845), .A4(n1844), .ZN(n1858)
         );
  AOI22_X1 U1297 ( .A1(n3010), .A2(mem[571]), .B1(n1051), .B2(mem[155]), .ZN(
        n1851) );
  AOI22_X1 U1298 ( .A1(n1045), .A2(mem[27]), .B1(n1044), .B2(mem[827]), .ZN(
        n1850) );
  AOI22_X1 U1299 ( .A1(n2874), .A2(mem[379]), .B1(n2750), .B2(mem[539]), .ZN(
        n1849) );
  AOI22_X1 U1300 ( .A1(n2433), .A2(mem[603]), .B1(n3001), .B2(mem[59]), .ZN(
        n1848) );
  NAND4_X1 U1301 ( .A1(n1851), .A2(n1850), .A3(n1849), .A4(n1848), .ZN(n1857)
         );
  AOI22_X1 U1302 ( .A1(n1043), .A2(mem[123]), .B1(n1056), .B2(mem[891]), .ZN(
        n1855) );
  AOI22_X1 U1303 ( .A1(n1050), .A2(mem[859]), .B1(n1040), .B2(mem[219]), .ZN(
        n1854) );
  AOI22_X1 U1304 ( .A1(n3016), .A2(mem[315]), .B1(n1039), .B2(mem[955]), .ZN(
        n1853) );
  AOI22_X1 U1305 ( .A1(n1042), .A2(mem[251]), .B1(n1046), .B2(mem[475]), .ZN(
        n1852) );
  NAND4_X1 U1306 ( .A1(n1855), .A2(n1854), .A3(n1853), .A4(n1852), .ZN(n1856)
         );
  OR4_X1 U1307 ( .A1(n1859), .A2(n1858), .A3(n1857), .A4(n1856), .ZN(
        rdata_c_o[27]) );
  AOI22_X1 U1308 ( .A1(n2968), .A2(mem[923]), .B1(n2976), .B2(mem[315]), .ZN(
        n1863) );
  AOI22_X1 U1309 ( .A1(n2764), .A2(mem[763]), .B1(n2965), .B2(mem[507]), .ZN(
        n1862) );
  AOI22_X1 U1310 ( .A1(n2860), .A2(mem[187]), .B1(n2954), .B2(mem[379]), .ZN(
        n1861) );
  NAND2_X1 U1311 ( .A1(n2850), .A2(mem[699]), .ZN(n1860) );
  NAND4_X1 U1312 ( .A1(n1863), .A2(n1862), .A3(n1861), .A4(n1860), .ZN(n1879)
         );
  AOI22_X1 U1313 ( .A1(n2952), .A2(mem[475]), .B1(n2966), .B2(mem[91]), .ZN(
        n1867) );
  AOI22_X1 U1314 ( .A1(n2992), .A2(mem[891]), .B1(n2991), .B2(mem[571]), .ZN(
        n1866) );
  AOI22_X1 U1315 ( .A1(n2796), .A2(mem[667]), .B1(n2957), .B2(mem[251]), .ZN(
        n1865) );
  AOI22_X1 U1316 ( .A1(n2977), .A2(mem[219]), .B1(n2951), .B2(mem[155]), .ZN(
        n1864) );
  NAND4_X1 U1317 ( .A1(n1867), .A2(n1866), .A3(n1865), .A4(n1864), .ZN(n1878)
         );
  AOI22_X1 U1318 ( .A1(n2978), .A2(mem[283]), .B1(n2987), .B2(mem[411]), .ZN(
        n1871) );
  AOI22_X1 U1319 ( .A1(n2956), .A2(mem[635]), .B1(n2988), .B2(mem[539]), .ZN(
        n1870) );
  AOI22_X1 U1320 ( .A1(n2990), .A2(mem[59]), .B1(n2975), .B2(mem[795]), .ZN(
        n1869) );
  AOI22_X1 U1321 ( .A1(n2797), .A2(mem[955]), .B1(n2986), .B2(mem[603]), .ZN(
        n1868) );
  NAND4_X1 U1322 ( .A1(n1871), .A2(n1870), .A3(n1869), .A4(n1868), .ZN(n1877)
         );
  AOI22_X1 U1323 ( .A1(n2791), .A2(mem[987]), .B1(n2953), .B2(mem[731]), .ZN(
        n1875) );
  AOI22_X1 U1324 ( .A1(n2639), .A2(mem[859]), .B1(n2834), .B2(mem[27]), .ZN(
        n1874) );
  AOI22_X1 U1325 ( .A1(n2843), .A2(mem[123]), .B1(n2985), .B2(mem[347]), .ZN(
        n1873) );
  AOI22_X1 U1326 ( .A1(n2840), .A2(mem[827]), .B1(n2832), .B2(mem[443]), .ZN(
        n1872) );
  NAND4_X1 U1327 ( .A1(n1875), .A2(n1874), .A3(n1873), .A4(n1872), .ZN(n1876)
         );
  OR4_X1 U1328 ( .A1(n1879), .A2(n1878), .A3(n1877), .A4(n1876), .ZN(
        rdata_b_o[27]) );
  AOI22_X1 U1329 ( .A1(n2968), .A2(mem[922]), .B1(n2848), .B2(mem[282]), .ZN(
        n1883) );
  AOI22_X1 U1330 ( .A1(n2955), .A2(mem[826]), .B1(n2835), .B2(mem[538]), .ZN(
        n1882) );
  AOI22_X1 U1331 ( .A1(n2786), .A2(mem[570]), .B1(n2953), .B2(mem[730]), .ZN(
        n1881) );
  NAND2_X1 U1332 ( .A1(n2853), .A2(mem[890]), .ZN(n1880) );
  NAND4_X1 U1333 ( .A1(n1883), .A2(n1882), .A3(n1881), .A4(n1880), .ZN(n1899)
         );
  AOI22_X1 U1334 ( .A1(n2770), .A2(mem[634]), .B1(n2966), .B2(mem[90]), .ZN(
        n1887) );
  AOI22_X1 U1335 ( .A1(n2775), .A2(mem[58]), .B1(n2976), .B2(mem[314]), .ZN(
        n1886) );
  AOI22_X1 U1336 ( .A1(n2977), .A2(mem[218]), .B1(n2849), .B2(mem[506]), .ZN(
        n1885) );
  AOI22_X1 U1337 ( .A1(n2986), .A2(mem[602]), .B1(n2860), .B2(mem[186]), .ZN(
        n1884) );
  NAND4_X1 U1338 ( .A1(n1887), .A2(n1886), .A3(n1885), .A4(n1884), .ZN(n1898)
         );
  AOI22_X1 U1339 ( .A1(n2969), .A2(mem[698]), .B1(n2834), .B2(mem[26]), .ZN(
        n1891) );
  AOI22_X1 U1340 ( .A1(n2952), .A2(mem[474]), .B1(n2639), .B2(mem[858]), .ZN(
        n1890) );
  AOI22_X1 U1341 ( .A1(n2980), .A2(mem[762]), .B1(n2803), .B2(mem[250]), .ZN(
        n1889) );
  AOI22_X1 U1342 ( .A1(n2975), .A2(mem[794]), .B1(n2859), .B2(mem[154]), .ZN(
        n1888) );
  NAND4_X1 U1343 ( .A1(n1891), .A2(n1890), .A3(n1889), .A4(n1888), .ZN(n1897)
         );
  AOI22_X1 U1344 ( .A1(n2797), .A2(mem[954]), .B1(n2759), .B2(mem[346]), .ZN(
        n1895) );
  AOI22_X1 U1345 ( .A1(n2989), .A2(mem[986]), .B1(n2987), .B2(mem[410]), .ZN(
        n1894) );
  AOI22_X1 U1346 ( .A1(n2843), .A2(mem[122]), .B1(n2832), .B2(mem[442]), .ZN(
        n1893) );
  AOI22_X1 U1347 ( .A1(n2967), .A2(mem[666]), .B1(n2842), .B2(mem[378]), .ZN(
        n1892) );
  NAND4_X1 U1348 ( .A1(n1895), .A2(n1894), .A3(n1893), .A4(n1892), .ZN(n1896)
         );
  OR4_X1 U1349 ( .A1(n1899), .A2(n1898), .A3(n1897), .A4(n1896), .ZN(
        rdata_b_o[26]) );
  AOI22_X1 U1350 ( .A1(n1052), .A2(mem[698]), .B1(n1047), .B2(mem[90]), .ZN(
        n1903) );
  AOI22_X1 U1351 ( .A1(n2750), .A2(mem[538]), .B1(n1056), .B2(mem[890]), .ZN(
        n1902) );
  AOI22_X1 U1352 ( .A1(n1054), .A2(mem[346]), .B1(n1046), .B2(mem[474]), .ZN(
        n1901) );
  NAND2_X1 U1353 ( .A1(n1042), .A2(mem[250]), .ZN(n1900) );
  NAND4_X1 U1354 ( .A1(n1903), .A2(n1902), .A3(n1901), .A4(n1900), .ZN(n1919)
         );
  AOI22_X1 U1355 ( .A1(n1055), .A2(mem[986]), .B1(n2705), .B2(mem[762]), .ZN(
        n1907) );
  AOI22_X1 U1356 ( .A1(n2668), .A2(mem[634]), .B1(n1048), .B2(mem[794]), .ZN(
        n1906) );
  AOI22_X1 U1357 ( .A1(n1033), .A2(mem[410]), .B1(n3015), .B2(mem[730]), .ZN(
        n1905) );
  AOI22_X1 U1358 ( .A1(n2874), .A2(mem[378]), .B1(n1043), .B2(mem[122]), .ZN(
        n1904) );
  NAND4_X1 U1359 ( .A1(n1907), .A2(n1906), .A3(n1905), .A4(n1904), .ZN(n1918)
         );
  AOI22_X1 U1360 ( .A1(n2433), .A2(mem[602]), .B1(n1051), .B2(mem[154]), .ZN(
        n1911) );
  AOI22_X1 U1361 ( .A1(n3001), .A2(mem[58]), .B1(n1040), .B2(mem[218]), .ZN(
        n1910) );
  AOI22_X1 U1362 ( .A1(n1039), .A2(mem[954]), .B1(n1041), .B2(mem[186]), .ZN(
        n1909) );
  AOI22_X1 U1363 ( .A1(n1050), .A2(mem[858]), .B1(n1395), .B2(mem[314]), .ZN(
        n1908) );
  NAND4_X1 U1364 ( .A1(n1911), .A2(n1910), .A3(n1909), .A4(n1908), .ZN(n1917)
         );
  AOI22_X1 U1365 ( .A1(n1045), .A2(mem[26]), .B1(n1049), .B2(mem[282]), .ZN(
        n1915) );
  AOI22_X1 U1366 ( .A1(n2062), .A2(mem[506]), .B1(n1044), .B2(mem[826]), .ZN(
        n1914) );
  AOI22_X1 U1367 ( .A1(n1403), .A2(mem[922]), .B1(n3010), .B2(mem[570]), .ZN(
        n1913) );
  AOI22_X1 U1368 ( .A1(n1053), .A2(mem[442]), .B1(n2578), .B2(mem[666]), .ZN(
        n1912) );
  NAND4_X1 U1369 ( .A1(n1915), .A2(n1914), .A3(n1913), .A4(n1912), .ZN(n1916)
         );
  OR4_X1 U1370 ( .A1(n1919), .A2(n1918), .A3(n1917), .A4(n1916), .ZN(
        rdata_c_o[26]) );
  AOI22_X1 U1371 ( .A1(n2853), .A2(mem[893]), .B1(n2968), .B2(mem[925]), .ZN(
        n1923) );
  AOI22_X1 U1372 ( .A1(n2956), .A2(mem[637]), .B1(n2962), .B2(mem[861]), .ZN(
        n1922) );
  AOI22_X1 U1373 ( .A1(n2843), .A2(mem[125]), .B1(n2953), .B2(mem[733]), .ZN(
        n1921) );
  NAND2_X1 U1374 ( .A1(n2966), .A2(mem[93]), .ZN(n1920) );
  NAND4_X1 U1375 ( .A1(n1923), .A2(n1922), .A3(n1921), .A4(n1920), .ZN(n1939)
         );
  AOI22_X1 U1376 ( .A1(n2963), .A2(mem[957]), .B1(n2832), .B2(mem[445]), .ZN(
        n1927) );
  AOI22_X1 U1377 ( .A1(n2957), .A2(mem[253]), .B1(n2955), .B2(mem[829]), .ZN(
        n1926) );
  AOI22_X1 U1378 ( .A1(n2969), .A2(mem[701]), .B1(n2848), .B2(mem[285]), .ZN(
        n1925) );
  AOI22_X1 U1379 ( .A1(n2990), .A2(mem[61]), .B1(n2951), .B2(mem[157]), .ZN(
        n1924) );
  NAND4_X1 U1380 ( .A1(n1927), .A2(n1926), .A3(n1925), .A4(n1924), .ZN(n1938)
         );
  AOI22_X1 U1381 ( .A1(n2975), .A2(mem[797]), .B1(n2965), .B2(mem[509]), .ZN(
        n1931) );
  AOI22_X1 U1382 ( .A1(n2791), .A2(mem[989]), .B1(n2979), .B2(mem[29]), .ZN(
        n1930) );
  AOI22_X1 U1383 ( .A1(n2977), .A2(mem[221]), .B1(n2860), .B2(mem[189]), .ZN(
        n1929) );
  AOI22_X1 U1384 ( .A1(n2980), .A2(mem[765]), .B1(n2796), .B2(mem[669]), .ZN(
        n1928) );
  NAND4_X1 U1385 ( .A1(n1931), .A2(n1930), .A3(n1929), .A4(n1928), .ZN(n1937)
         );
  AOI22_X1 U1386 ( .A1(n2991), .A2(mem[573]), .B1(n2988), .B2(mem[541]), .ZN(
        n1935) );
  AOI22_X1 U1387 ( .A1(n2985), .A2(mem[349]), .B1(n2987), .B2(mem[413]), .ZN(
        n1934) );
  AOI22_X1 U1388 ( .A1(n2952), .A2(mem[477]), .B1(n2858), .B2(mem[317]), .ZN(
        n1933) );
  AOI22_X1 U1389 ( .A1(n2986), .A2(mem[605]), .B1(n2842), .B2(mem[381]), .ZN(
        n1932) );
  NAND4_X1 U1390 ( .A1(n1935), .A2(n1934), .A3(n1933), .A4(n1932), .ZN(n1936)
         );
  OR4_X1 U1391 ( .A1(n1939), .A2(n1938), .A3(n1937), .A4(n1936), .ZN(
        rdata_b_o[29]) );
  AOI22_X1 U1392 ( .A1(mem[381]), .A2(n1024), .B1(n3350), .B2(mem[317]), .ZN(
        n1943) );
  AOI22_X1 U1393 ( .A1(n1092), .A2(mem[509]), .B1(mem[61]), .B2(n4729), .ZN(
        n1942) );
  AOI22_X1 U1394 ( .A1(mem[93]), .A2(n3512), .B1(n3578), .B2(mem[29]), .ZN(
        n1941) );
  NAND2_X1 U1395 ( .A1(n1025), .A2(mem[797]), .ZN(n1940) );
  NAND4_X1 U1396 ( .A1(n1943), .A2(n1942), .A3(n1941), .A4(n1940), .ZN(n1959)
         );
  BUF_X1 U1397 ( .A(n2153), .Z(n3382) );
  AOI22_X1 U1398 ( .A1(mem[701]), .A2(n1070), .B1(n3382), .B2(mem[413]), .ZN(
        n1947) );
  AOI22_X1 U1399 ( .A1(n1017), .A2(mem[221]), .B1(mem[125]), .B2(n1031), .ZN(
        n1946) );
  AOI22_X1 U1400 ( .A1(mem[637]), .A2(n1071), .B1(n3383), .B2(mem[573]), .ZN(
        n1945) );
  AOI22_X1 U1401 ( .A1(n3358), .A2(mem[669]), .B1(mem[189]), .B2(n1072), .ZN(
        n1944) );
  NAND4_X1 U1402 ( .A1(n1947), .A2(n1946), .A3(n1945), .A4(n1944), .ZN(n1958)
         );
  AOI22_X1 U1403 ( .A1(mem[605]), .A2(n1016), .B1(n994), .B2(mem[477]), .ZN(
        n1951) );
  AOI22_X1 U1404 ( .A1(mem[349]), .A2(n1007), .B1(n1084), .B2(mem[285]), .ZN(
        n1950) );
  AOI22_X1 U1405 ( .A1(mem[733]), .A2(n1081), .B1(n1011), .B2(mem[445]), .ZN(
        n1949) );
  AOI22_X1 U1406 ( .A1(n1009), .A2(mem[253]), .B1(mem[157]), .B2(n1021), .ZN(
        n1948) );
  NAND4_X1 U1407 ( .A1(n1951), .A2(n1950), .A3(n1949), .A4(n1948), .ZN(n1957)
         );
  AOI22_X1 U1408 ( .A1(n1068), .A2(mem[541]), .B1(mem[957]), .B2(n3592), .ZN(
        n1955) );
  AOI22_X1 U1409 ( .A1(mem[989]), .A2(n3564), .B1(n1086), .B2(mem[765]), .ZN(
        n1954) );
  AOI22_X1 U1410 ( .A1(mem[893]), .A2(n3593), .B1(n1069), .B2(mem[829]), .ZN(
        n1953) );
  AOI22_X1 U1411 ( .A1(mem[925]), .A2(n3594), .B1(n1091), .B2(mem[861]), .ZN(
        n1952) );
  NAND4_X1 U1412 ( .A1(n1955), .A2(n1954), .A3(n1953), .A4(n1952), .ZN(n1956)
         );
  OR4_X1 U1413 ( .A1(n1959), .A2(n1958), .A3(n1957), .A4(n1956), .ZN(
        rdata_a_o[29]) );
  AOI22_X1 U1414 ( .A1(n1033), .A2(mem[413]), .B1(n1051), .B2(mem[157]), .ZN(
        n1963) );
  AOI22_X1 U1415 ( .A1(n1740), .A2(mem[509]), .B1(n1055), .B2(mem[989]), .ZN(
        n1962) );
  AOI22_X1 U1416 ( .A1(n1052), .A2(mem[701]), .B1(n3010), .B2(mem[573]), .ZN(
        n1961) );
  NAND2_X1 U1417 ( .A1(n1395), .A2(mem[317]), .ZN(n1960) );
  NAND4_X1 U1418 ( .A1(n1963), .A2(n1962), .A3(n1961), .A4(n1960), .ZN(n1979)
         );
  AOI22_X1 U1419 ( .A1(n1752), .A2(mem[605]), .B1(n1040), .B2(mem[221]), .ZN(
        n1967) );
  AOI22_X1 U1420 ( .A1(n1042), .A2(mem[253]), .B1(n1046), .B2(mem[477]), .ZN(
        n1966) );
  AOI22_X1 U1421 ( .A1(n1751), .A2(mem[29]), .B1(n1049), .B2(mem[285]), .ZN(
        n1965) );
  AOI22_X1 U1422 ( .A1(n2750), .A2(mem[541]), .B1(n1048), .B2(mem[797]), .ZN(
        n1964) );
  NAND4_X1 U1423 ( .A1(n1967), .A2(n1966), .A3(n1965), .A4(n1964), .ZN(n1978)
         );
  AOI22_X1 U1424 ( .A1(n1054), .A2(mem[349]), .B1(n1461), .B2(mem[765]), .ZN(
        n1971) );
  AOI22_X1 U1425 ( .A1(n1041), .A2(mem[189]), .B1(n1056), .B2(mem[893]), .ZN(
        n1970) );
  AOI22_X1 U1426 ( .A1(n1403), .A2(mem[925]), .B1(n1047), .B2(mem[93]), .ZN(
        n1969) );
  AOI22_X1 U1427 ( .A1(n1452), .A2(mem[733]), .B1(n1043), .B2(mem[125]), .ZN(
        n1968) );
  NAND4_X1 U1428 ( .A1(n1971), .A2(n1970), .A3(n1969), .A4(n1968), .ZN(n1977)
         );
  AOI22_X1 U1429 ( .A1(n1745), .A2(mem[637]), .B1(n1044), .B2(mem[829]), .ZN(
        n1975) );
  AOI22_X1 U1430 ( .A1(n3001), .A2(mem[61]), .B1(n2578), .B2(mem[669]), .ZN(
        n1974) );
  AOI22_X1 U1431 ( .A1(n1039), .A2(mem[957]), .B1(n1053), .B2(mem[445]), .ZN(
        n1973) );
  AOI22_X1 U1432 ( .A1(n1050), .A2(mem[861]), .B1(n2874), .B2(mem[381]), .ZN(
        n1972) );
  NAND4_X1 U1433 ( .A1(n1975), .A2(n1974), .A3(n1973), .A4(n1972), .ZN(n1976)
         );
  OR4_X1 U1434 ( .A1(n1979), .A2(n1978), .A3(n1977), .A4(n1976), .ZN(
        rdata_c_o[29]) );
  INV_X1 U1435 ( .A(wdata_b_i[4]), .ZN(n4416) );
  INV_X1 U1480 ( .A(wdata_b_i[5]), .ZN(n4418) );
  AOI22_X1 U1486 ( .A1(n1045), .A2(mem[1]), .B1(n1054), .B2(mem[321]), .ZN(
        n2006) );
  AOI22_X1 U1487 ( .A1(n1033), .A2(mem[385]), .B1(n1042), .B2(mem[225]), .ZN(
        n2005) );
  AOI22_X1 U1488 ( .A1(n1040), .A2(mem[193]), .B1(n1056), .B2(mem[865]), .ZN(
        n2004) );
  NAND2_X1 U1489 ( .A1(n2433), .A2(mem[577]), .ZN(n2003) );
  NAND4_X1 U1490 ( .A1(n2006), .A2(n2005), .A3(n2004), .A4(n2003), .ZN(n2022)
         );
  AOI22_X1 U1491 ( .A1(n3016), .A2(mem[289]), .B1(n1049), .B2(mem[257]), .ZN(
        n2010) );
  AOI22_X1 U1492 ( .A1(n2869), .A2(mem[897]), .B1(n1047), .B2(mem[65]), .ZN(
        n2009) );
  AOI22_X1 U1493 ( .A1(n1039), .A2(mem[929]), .B1(n1431), .B2(mem[673]), .ZN(
        n2008) );
  AOI22_X1 U1494 ( .A1(n2062), .A2(mem[481]), .B1(n2874), .B2(mem[353]), .ZN(
        n2007) );
  NAND4_X1 U1495 ( .A1(n2010), .A2(n2009), .A3(n2008), .A4(n2007), .ZN(n2021)
         );
  AOI22_X1 U1496 ( .A1(n2668), .A2(mem[609]), .B1(n2578), .B2(mem[641]), .ZN(
        n2014) );
  AOI22_X1 U1497 ( .A1(n3001), .A2(mem[33]), .B1(n1046), .B2(mem[449]), .ZN(
        n2013) );
  AOI22_X1 U1498 ( .A1(n1055), .A2(mem[961]), .B1(n1044), .B2(mem[801]), .ZN(
        n2012) );
  AOI22_X1 U1499 ( .A1(n1050), .A2(mem[833]), .B1(n1041), .B2(mem[161]), .ZN(
        n2011) );
  NAND4_X1 U1500 ( .A1(n2014), .A2(n2013), .A3(n2012), .A4(n2011), .ZN(n2020)
         );
  AOI22_X1 U1501 ( .A1(n3015), .A2(mem[705]), .B1(n2705), .B2(mem[737]), .ZN(
        n2018) );
  AOI22_X1 U1502 ( .A1(n1048), .A2(mem[769]), .B1(n1043), .B2(mem[97]), .ZN(
        n2017) );
  AOI22_X1 U1503 ( .A1(n1053), .A2(mem[417]), .B1(n3010), .B2(mem[545]), .ZN(
        n2016) );
  AOI22_X1 U1504 ( .A1(n2750), .A2(mem[513]), .B1(n1051), .B2(mem[129]), .ZN(
        n2015) );
  NAND4_X1 U1505 ( .A1(n2018), .A2(n2017), .A3(n2016), .A4(n2015), .ZN(n2019)
         );
  OR4_X1 U1506 ( .A1(n2022), .A2(n2021), .A3(n2020), .A4(n2019), .ZN(
        rdata_c_o[1]) );
  AOI22_X1 U1546 ( .A1(n2852), .A2(mem[788]), .B1(n2965), .B2(mem[500]), .ZN(
        n2045) );
  AOI22_X1 U1547 ( .A1(n2759), .A2(mem[340]), .B1(n2841), .B2(mem[724]), .ZN(
        n2044) );
  AOI22_X1 U1548 ( .A1(n2989), .A2(mem[980]), .B1(n2776), .B2(mem[212]), .ZN(
        n2043) );
  NAND2_X1 U1549 ( .A1(n2848), .A2(mem[276]), .ZN(n2042) );
  NAND4_X1 U1550 ( .A1(n2045), .A2(n2044), .A3(n2043), .A4(n2042), .ZN(n2061)
         );
  AOI22_X1 U1551 ( .A1(n2832), .A2(mem[436]), .B1(n2979), .B2(mem[20]), .ZN(
        n2049) );
  AOI22_X1 U1552 ( .A1(n2976), .A2(mem[308]), .B1(n2835), .B2(mem[532]), .ZN(
        n2048) );
  AOI22_X1 U1553 ( .A1(n2765), .A2(mem[596]), .B1(n2966), .B2(mem[84]), .ZN(
        n2047) );
  AOI22_X1 U1554 ( .A1(n2992), .A2(mem[884]), .B1(n2833), .B2(mem[468]), .ZN(
        n2046) );
  NAND4_X1 U1555 ( .A1(n2049), .A2(n2048), .A3(n2047), .A4(n2046), .ZN(n2060)
         );
  AOI22_X1 U1556 ( .A1(n2860), .A2(mem[180]), .B1(n2786), .B2(mem[564]), .ZN(
        n2053) );
  AOI22_X1 U1557 ( .A1(n2797), .A2(mem[948]), .B1(n2968), .B2(mem[916]), .ZN(
        n2052) );
  AOI22_X1 U1558 ( .A1(n2969), .A2(mem[692]), .B1(n2796), .B2(mem[660]), .ZN(
        n2051) );
  AOI22_X1 U1559 ( .A1(n2803), .A2(mem[244]), .B1(n2951), .B2(mem[148]), .ZN(
        n2050) );
  NAND4_X1 U1560 ( .A1(n2053), .A2(n2052), .A3(n2051), .A4(n2050), .ZN(n2059)
         );
  AOI22_X1 U1561 ( .A1(n2770), .A2(mem[628]), .B1(n2955), .B2(mem[820]), .ZN(
        n2057) );
  AOI22_X1 U1562 ( .A1(n2639), .A2(mem[852]), .B1(n2842), .B2(mem[372]), .ZN(
        n2056) );
  AOI22_X1 U1563 ( .A1(n2974), .A2(mem[116]), .B1(n2987), .B2(mem[404]), .ZN(
        n2055) );
  AOI22_X1 U1564 ( .A1(n2980), .A2(mem[756]), .B1(n2775), .B2(mem[52]), .ZN(
        n2054) );
  NAND4_X1 U1565 ( .A1(n2057), .A2(n2056), .A3(n2055), .A4(n2054), .ZN(n2058)
         );
  OR4_X1 U1566 ( .A1(n2061), .A2(n2060), .A3(n2059), .A4(n2058), .ZN(
        rdata_b_o[20]) );
  AOI22_X1 U1567 ( .A1(n2668), .A2(mem[628]), .B1(n1044), .B2(mem[820]), .ZN(
        n2066) );
  AOI22_X1 U1568 ( .A1(n2750), .A2(mem[532]), .B1(n1056), .B2(mem[884]), .ZN(
        n2065) );
  AOI22_X1 U1569 ( .A1(n3001), .A2(mem[52]), .B1(n1053), .B2(mem[436]), .ZN(
        n2064) );
  NAND2_X1 U1570 ( .A1(n2062), .A2(mem[500]), .ZN(n2063) );
  NAND4_X1 U1571 ( .A1(n2066), .A2(n2065), .A3(n2064), .A4(n2063), .ZN(n2083)
         );
  AOI22_X1 U1572 ( .A1(n1040), .A2(mem[212]), .B1(n1043), .B2(mem[116]), .ZN(
        n2071) );
  AOI22_X1 U1573 ( .A1(n1751), .A2(mem[20]), .B1(n2578), .B2(mem[660]), .ZN(
        n2070) );
  AOI22_X1 U1574 ( .A1(n2874), .A2(mem[372]), .B1(n1049), .B2(mem[276]), .ZN(
        n2069) );
  AOI22_X1 U1575 ( .A1(n1039), .A2(mem[948]), .B1(n1461), .B2(mem[756]), .ZN(
        n2068) );
  NAND4_X1 U1576 ( .A1(n2071), .A2(n2070), .A3(n2069), .A4(n2068), .ZN(n2082)
         );
  AOI22_X1 U1577 ( .A1(n1752), .A2(mem[596]), .B1(n1046), .B2(mem[468]), .ZN(
        n2075) );
  AOI22_X1 U1578 ( .A1(n1055), .A2(mem[980]), .B1(n3010), .B2(mem[564]), .ZN(
        n2074) );
  AOI22_X1 U1579 ( .A1(n1042), .A2(mem[244]), .B1(n1051), .B2(mem[148]), .ZN(
        n2073) );
  AOI22_X1 U1580 ( .A1(n3016), .A2(mem[308]), .B1(n1054), .B2(mem[340]), .ZN(
        n2072) );
  NAND4_X1 U1581 ( .A1(n2075), .A2(n2074), .A3(n2073), .A4(n2072), .ZN(n2081)
         );
  AOI22_X1 U1582 ( .A1(n1050), .A2(mem[852]), .B1(n1047), .B2(mem[84]), .ZN(
        n2079) );
  AOI22_X1 U1583 ( .A1(n1041), .A2(mem[180]), .B1(n1048), .B2(mem[788]), .ZN(
        n2078) );
  AOI22_X1 U1584 ( .A1(n1403), .A2(mem[916]), .B1(n3015), .B2(mem[724]), .ZN(
        n2077) );
  AOI22_X1 U1585 ( .A1(n1033), .A2(mem[404]), .B1(n1052), .B2(mem[692]), .ZN(
        n2076) );
  NAND4_X1 U1586 ( .A1(n2079), .A2(n2078), .A3(n2077), .A4(n2076), .ZN(n2080)
         );
  OR4_X1 U1587 ( .A1(n2083), .A2(n2082), .A3(n2081), .A4(n2080), .ZN(
        rdata_c_o[20]) );
  INV_X1 U1588 ( .A(wdata_b_i[2]), .ZN(n4412) );
  AOI22_X1 U1594 ( .A1(n2433), .A2(mem[588]), .B1(n1043), .B2(mem[108]), .ZN(
        n2089) );
  AOI22_X1 U1595 ( .A1(n1047), .A2(mem[76]), .B1(n1049), .B2(mem[268]), .ZN(
        n2088) );
  AOI22_X1 U1596 ( .A1(n2874), .A2(mem[364]), .B1(n3015), .B2(mem[716]), .ZN(
        n2087) );
  NAND2_X1 U1597 ( .A1(n1055), .A2(mem[972]), .ZN(n2086) );
  NAND4_X1 U1598 ( .A1(n2089), .A2(n2088), .A3(n2087), .A4(n2086), .ZN(n2105)
         );
  AOI22_X1 U1599 ( .A1(n1053), .A2(mem[428]), .B1(n1046), .B2(mem[460]), .ZN(
        n2093) );
  AOI22_X1 U1600 ( .A1(n1048), .A2(mem[780]), .B1(n3010), .B2(mem[556]), .ZN(
        n2092) );
  AOI22_X1 U1601 ( .A1(n2062), .A2(mem[492]), .B1(n2869), .B2(mem[908]), .ZN(
        n2091) );
  AOI22_X1 U1602 ( .A1(n1033), .A2(mem[396]), .B1(n2578), .B2(mem[652]), .ZN(
        n2090) );
  NAND4_X1 U1603 ( .A1(n2093), .A2(n2092), .A3(n2091), .A4(n2090), .ZN(n2104)
         );
  AOI22_X1 U1604 ( .A1(n2705), .A2(mem[748]), .B1(n1051), .B2(mem[140]), .ZN(
        n2097) );
  AOI22_X1 U1605 ( .A1(n3016), .A2(mem[300]), .B1(n1041), .B2(mem[172]), .ZN(
        n2096) );
  AOI22_X1 U1606 ( .A1(n1045), .A2(mem[12]), .B1(n1040), .B2(mem[204]), .ZN(
        n2095) );
  AOI22_X1 U1607 ( .A1(n1745), .A2(mem[620]), .B1(n3001), .B2(mem[44]), .ZN(
        n2094) );
  NAND4_X1 U1608 ( .A1(n2097), .A2(n2096), .A3(n2095), .A4(n2094), .ZN(n2103)
         );
  AOI22_X1 U1609 ( .A1(n1042), .A2(mem[236]), .B1(n2750), .B2(mem[524]), .ZN(
        n2101) );
  AOI22_X1 U1610 ( .A1(n1054), .A2(mem[332]), .B1(n1056), .B2(mem[876]), .ZN(
        n2100) );
  AOI22_X1 U1611 ( .A1(n1039), .A2(mem[940]), .B1(n1044), .B2(mem[812]), .ZN(
        n2099) );
  AOI22_X1 U1612 ( .A1(n1050), .A2(mem[844]), .B1(n1052), .B2(mem[684]), .ZN(
        n2098) );
  NAND4_X1 U1613 ( .A1(n2101), .A2(n2100), .A3(n2099), .A4(n2098), .ZN(n2102)
         );
  OR4_X1 U1614 ( .A1(n2105), .A2(n2104), .A3(n2103), .A4(n2102), .ZN(
        rdata_c_o[12]) );
  AOI22_X1 U1615 ( .A1(n2764), .A2(mem[748]), .B1(n2786), .B2(mem[556]), .ZN(
        n2109) );
  AOI22_X1 U1616 ( .A1(n2963), .A2(mem[940]), .B1(n2775), .B2(mem[44]), .ZN(
        n2108) );
  AOI22_X1 U1617 ( .A1(n2759), .A2(mem[332]), .B1(n2851), .B2(mem[396]), .ZN(
        n2107) );
  NAND2_X1 U1618 ( .A1(n2860), .A2(mem[172]), .ZN(n2106) );
  NAND4_X1 U1619 ( .A1(n2109), .A2(n2108), .A3(n2107), .A4(n2106), .ZN(n2125)
         );
  AOI22_X1 U1620 ( .A1(n2989), .A2(mem[972]), .B1(n2966), .B2(mem[76]), .ZN(
        n2113) );
  AOI22_X1 U1621 ( .A1(n2965), .A2(mem[492]), .B1(n2955), .B2(mem[812]), .ZN(
        n2112) );
  AOI22_X1 U1622 ( .A1(n2853), .A2(mem[876]), .B1(n2852), .B2(mem[780]), .ZN(
        n2111) );
  AOI22_X1 U1623 ( .A1(n2848), .A2(mem[268]), .B1(n2953), .B2(mem[716]), .ZN(
        n2110) );
  NAND4_X1 U1624 ( .A1(n2113), .A2(n2112), .A3(n2111), .A4(n2110), .ZN(n2124)
         );
  AOI22_X1 U1625 ( .A1(n2962), .A2(mem[844]), .B1(n2977), .B2(mem[204]), .ZN(
        n2117) );
  AOI22_X1 U1626 ( .A1(n2858), .A2(mem[300]), .B1(n2964), .B2(mem[428]), .ZN(
        n2116) );
  AOI22_X1 U1627 ( .A1(n2765), .A2(mem[588]), .B1(n2951), .B2(mem[140]), .ZN(
        n2115) );
  AOI22_X1 U1628 ( .A1(n2770), .A2(mem[620]), .B1(n2785), .B2(mem[908]), .ZN(
        n2114) );
  NAND4_X1 U1629 ( .A1(n2117), .A2(n2116), .A3(n2115), .A4(n2114), .ZN(n2123)
         );
  AOI22_X1 U1630 ( .A1(n2954), .A2(mem[364]), .B1(n2979), .B2(mem[12]), .ZN(
        n2121) );
  AOI22_X1 U1631 ( .A1(n2957), .A2(mem[236]), .B1(n2835), .B2(mem[524]), .ZN(
        n2120) );
  AOI22_X1 U1632 ( .A1(n2833), .A2(mem[460]), .B1(n2974), .B2(mem[108]), .ZN(
        n2119) );
  AOI22_X1 U1633 ( .A1(n2850), .A2(mem[684]), .B1(n2796), .B2(mem[652]), .ZN(
        n2118) );
  NAND4_X1 U1634 ( .A1(n2121), .A2(n2120), .A3(n2119), .A4(n2118), .ZN(n2122)
         );
  OR4_X1 U1635 ( .A1(n2125), .A2(n2124), .A3(n2123), .A4(n2122), .ZN(
        rdata_b_o[12]) );
  AOI22_X1 U1636 ( .A1(n1053), .A2(mem[424]), .B1(n1046), .B2(mem[456]), .ZN(
        n2129) );
  AOI22_X1 U1637 ( .A1(n1055), .A2(mem[968]), .B1(n1054), .B2(mem[328]), .ZN(
        n2128) );
  AOI22_X1 U1638 ( .A1(n1047), .A2(mem[72]), .B1(n1049), .B2(mem[264]), .ZN(
        n2127) );
  NAND2_X1 U1639 ( .A1(n1042), .A2(mem[232]), .ZN(n2126) );
  NAND4_X1 U1640 ( .A1(n2129), .A2(n2128), .A3(n2127), .A4(n2126), .ZN(n2145)
         );
  AOI22_X1 U1641 ( .A1(n2668), .A2(mem[616]), .B1(n2705), .B2(mem[744]), .ZN(
        n2133) );
  AOI22_X1 U1642 ( .A1(n2578), .A2(mem[648]), .B1(n2750), .B2(mem[520]), .ZN(
        n2132) );
  AOI22_X1 U1643 ( .A1(n1052), .A2(mem[680]), .B1(n1051), .B2(mem[136]), .ZN(
        n2131) );
  AOI22_X1 U1644 ( .A1(n1045), .A2(mem[8]), .B1(n1041), .B2(mem[168]), .ZN(
        n2130) );
  NAND4_X1 U1645 ( .A1(n2133), .A2(n2132), .A3(n2131), .A4(n2130), .ZN(n2144)
         );
  AOI22_X1 U1646 ( .A1(n1044), .A2(mem[808]), .B1(n1408), .B2(mem[104]), .ZN(
        n2137) );
  AOI22_X1 U1647 ( .A1(n1424), .A2(mem[360]), .B1(n2869), .B2(mem[904]), .ZN(
        n2136) );
  AOI22_X1 U1648 ( .A1(n1033), .A2(mem[392]), .B1(n1048), .B2(mem[776]), .ZN(
        n2135) );
  AOI22_X1 U1649 ( .A1(n2433), .A2(mem[584]), .B1(n1395), .B2(mem[296]), .ZN(
        n2134) );
  NAND4_X1 U1650 ( .A1(n2137), .A2(n2136), .A3(n2135), .A4(n2134), .ZN(n2143)
         );
  AOI22_X1 U1651 ( .A1(n1039), .A2(mem[936]), .B1(n3010), .B2(mem[552]), .ZN(
        n2141) );
  AOI22_X1 U1652 ( .A1(n1414), .A2(mem[40]), .B1(n1056), .B2(mem[872]), .ZN(
        n2140) );
  AOI22_X1 U1653 ( .A1(n1050), .A2(mem[840]), .B1(n3015), .B2(mem[712]), .ZN(
        n2139) );
  AOI22_X1 U1654 ( .A1(n2062), .A2(mem[488]), .B1(n1040), .B2(mem[200]), .ZN(
        n2138) );
  NAND4_X1 U1655 ( .A1(n2141), .A2(n2140), .A3(n2139), .A4(n2138), .ZN(n2142)
         );
  OR4_X1 U1656 ( .A1(n2145), .A2(n2144), .A3(n2143), .A4(n2142), .ZN(
        rdata_c_o[8]) );
  AOI22_X1 U1657 ( .A1(mem[581]), .A2(n1016), .B1(n995), .B2(mem[453]), .ZN(
        n2152) );
  AOI22_X1 U1658 ( .A1(mem[325]), .A2(n1007), .B1(n1084), .B2(mem[261]), .ZN(
        n2151) );
  AOI22_X1 U1659 ( .A1(mem[709]), .A2(n1081), .B1(n1012), .B2(mem[421]), .ZN(
        n2150) );
  AOI22_X1 U1660 ( .A1(n1009), .A2(mem[229]), .B1(mem[133]), .B2(n1022), .ZN(
        n2149) );
  BUF_X1 U1661 ( .A(n2153), .Z(n3112) );
  AOI22_X1 U1662 ( .A1(mem[677]), .A2(n3161), .B1(n3112), .B2(mem[389]), .ZN(
        n2160) );
  BUF_X1 U1663 ( .A(n2154), .Z(n3113) );
  AOI22_X1 U1664 ( .A1(mem[613]), .A2(n3162), .B1(n3113), .B2(mem[549]), .ZN(
        n2159) );
  AOI22_X1 U1665 ( .A1(mem[101]), .A2(n1029), .B1(n1017), .B2(mem[197]), .ZN(
        n2158) );
  AOI22_X1 U1666 ( .A1(n3587), .A2(mem[645]), .B1(mem[165]), .B2(n1072), .ZN(
        n2157) );
  AOI22_X1 U1667 ( .A1(mem[357]), .A2(n1024), .B1(n2162), .B2(mem[293]), .ZN(
        n2168) );
  AOI22_X1 U1668 ( .A1(mem[69]), .A2(n3234), .B1(n3131), .B2(mem[5]), .ZN(
        n2167) );
  AOI22_X1 U1669 ( .A1(n1092), .A2(mem[485]), .B1(mem[37]), .B2(n4729), .ZN(
        n2166) );
  NAND2_X1 U1670 ( .A1(n1025), .A2(mem[773]), .ZN(n2165) );
  BUF_X1 U1671 ( .A(n3040), .Z(n3221) );
  AOI22_X1 U1672 ( .A1(n3167), .A2(mem[517]), .B1(mem[933]), .B2(n3221), .ZN(
        n2174) );
  AOI22_X1 U1673 ( .A1(mem[965]), .A2(n1073), .B1(n1086), .B2(mem[741]), .ZN(
        n2173) );
  AOI22_X1 U1674 ( .A1(mem[869]), .A2(n3066), .B1(n1069), .B2(mem[805]), .ZN(
        n2172) );
  AOI22_X1 U1675 ( .A1(mem[901]), .A2(n3269), .B1(n1089), .B2(mem[837]), .ZN(
        n2171) );
  AOI22_X1 U1676 ( .A1(mem[580]), .A2(n1015), .B1(n994), .B2(mem[452]), .ZN(
        n2178) );
  AOI22_X1 U1677 ( .A1(mem[324]), .A2(n1006), .B1(n1084), .B2(mem[260]), .ZN(
        n2177) );
  AOI22_X1 U1678 ( .A1(mem[708]), .A2(n1082), .B1(n1013), .B2(mem[420]), .ZN(
        n2176) );
  AOI22_X1 U1679 ( .A1(n1009), .A2(mem[228]), .B1(mem[132]), .B2(n1021), .ZN(
        n2175) );
  NAND4_X1 U1680 ( .A1(n2178), .A2(n2177), .A3(n2176), .A4(n2175), .ZN(n2194)
         );
  AOI22_X1 U1681 ( .A1(mem[676]), .A2(n3161), .B1(n3112), .B2(mem[388]), .ZN(
        n2182) );
  AOI22_X1 U1682 ( .A1(mem[612]), .A2(n3162), .B1(n3113), .B2(mem[548]), .ZN(
        n2181) );
  AOI22_X1 U1683 ( .A1(mem[100]), .A2(n1029), .B1(n1017), .B2(mem[196]), .ZN(
        n2180) );
  AOI22_X1 U1684 ( .A1(n3358), .A2(mem[644]), .B1(mem[164]), .B2(n3517), .ZN(
        n2179) );
  NAND4_X1 U1685 ( .A1(n2182), .A2(n2181), .A3(n2180), .A4(n2179), .ZN(n2193)
         );
  AOI22_X1 U1686 ( .A1(mem[356]), .A2(n1023), .B1(n2162), .B2(mem[292]), .ZN(
        n2186) );
  AOI22_X1 U1687 ( .A1(mem[68]), .A2(n3234), .B1(n3131), .B2(mem[4]), .ZN(
        n2185) );
  AOI22_X1 U1688 ( .A1(n1093), .A2(mem[484]), .B1(mem[36]), .B2(n4729), .ZN(
        n2184) );
  NAND2_X1 U1689 ( .A1(n1025), .A2(mem[772]), .ZN(n2183) );
  NAND4_X1 U1690 ( .A1(n2186), .A2(n2185), .A3(n2184), .A4(n2183), .ZN(n2192)
         );
  AOI22_X1 U1691 ( .A1(n3167), .A2(mem[516]), .B1(mem[932]), .B2(n3221), .ZN(
        n2190) );
  AOI22_X1 U1692 ( .A1(mem[964]), .A2(n1073), .B1(n1087), .B2(mem[740]), .ZN(
        n2189) );
  AOI22_X1 U1693 ( .A1(mem[868]), .A2(n3066), .B1(n3168), .B2(mem[804]), .ZN(
        n2188) );
  AOI22_X1 U1694 ( .A1(mem[900]), .A2(n3269), .B1(n1090), .B2(mem[836]), .ZN(
        n2187) );
  NAND4_X1 U1695 ( .A1(n2190), .A2(n2189), .A3(n2188), .A4(n2187), .ZN(n2191)
         );
  AOI22_X1 U1697 ( .A1(n1045), .A2(mem[9]), .B1(n1044), .B2(mem[809]), .ZN(
        n2198) );
  AOI22_X1 U1698 ( .A1(n1033), .A2(mem[393]), .B1(n1053), .B2(mem[425]), .ZN(
        n2197) );
  AOI22_X1 U1699 ( .A1(n3016), .A2(mem[297]), .B1(n1056), .B2(mem[873]), .ZN(
        n2196) );
  NAND2_X1 U1700 ( .A1(n1452), .A2(mem[713]), .ZN(n2195) );
  NAND4_X1 U1701 ( .A1(n2198), .A2(n2197), .A3(n2196), .A4(n2195), .ZN(n2214)
         );
  AOI22_X1 U1702 ( .A1(n1414), .A2(mem[41]), .B1(n2750), .B2(mem[521]), .ZN(
        n2202) );
  AOI22_X1 U1703 ( .A1(n1752), .A2(mem[585]), .B1(n1046), .B2(mem[457]), .ZN(
        n2201) );
  AOI22_X1 U1704 ( .A1(n1054), .A2(mem[329]), .B1(n3010), .B2(mem[553]), .ZN(
        n2200) );
  AOI22_X1 U1705 ( .A1(n1740), .A2(mem[489]), .B1(n1052), .B2(mem[681]), .ZN(
        n2199) );
  NAND4_X1 U1706 ( .A1(n2202), .A2(n2201), .A3(n2200), .A4(n2199), .ZN(n2213)
         );
  AOI22_X1 U1707 ( .A1(n1055), .A2(mem[969]), .B1(n1049), .B2(mem[265]), .ZN(
        n2206) );
  AOI22_X1 U1708 ( .A1(n1050), .A2(mem[841]), .B1(n1039), .B2(mem[937]), .ZN(
        n2205) );
  AOI22_X1 U1709 ( .A1(n2578), .A2(mem[649]), .B1(n1051), .B2(mem[137]), .ZN(
        n2204) );
  AOI22_X1 U1710 ( .A1(n2668), .A2(mem[617]), .B1(n1040), .B2(mem[201]), .ZN(
        n2203) );
  NAND4_X1 U1711 ( .A1(n2206), .A2(n2205), .A3(n2204), .A4(n2203), .ZN(n2212)
         );
  AOI22_X1 U1712 ( .A1(n1041), .A2(mem[169]), .B1(n1042), .B2(mem[233]), .ZN(
        n2210) );
  AOI22_X1 U1713 ( .A1(n2869), .A2(mem[905]), .B1(n1043), .B2(mem[105]), .ZN(
        n2209) );
  AOI22_X1 U1714 ( .A1(n1424), .A2(mem[361]), .B1(n1047), .B2(mem[73]), .ZN(
        n2208) );
  AOI22_X1 U1715 ( .A1(n2705), .A2(mem[745]), .B1(n1048), .B2(mem[777]), .ZN(
        n2207) );
  NAND4_X1 U1716 ( .A1(n2210), .A2(n2209), .A3(n2208), .A4(n2207), .ZN(n2211)
         );
  OR4_X1 U1717 ( .A1(n2214), .A2(n2213), .A3(n2212), .A4(n2211), .ZN(
        rdata_c_o[9]) );
  AOI22_X1 U1723 ( .A1(n2869), .A2(mem[909]), .B1(n1042), .B2(mem[237]), .ZN(
        n2220) );
  AOI22_X1 U1724 ( .A1(n3016), .A2(mem[301]), .B1(n1048), .B2(mem[781]), .ZN(
        n2219) );
  AOI22_X1 U1725 ( .A1(n1052), .A2(mem[685]), .B1(n1043), .B2(mem[109]), .ZN(
        n2218) );
  NAND2_X1 U1726 ( .A1(n3001), .A2(mem[45]), .ZN(n2217) );
  NAND4_X1 U1727 ( .A1(n2220), .A2(n2219), .A3(n2218), .A4(n2217), .ZN(n2236)
         );
  AOI22_X1 U1728 ( .A1(n2874), .A2(mem[365]), .B1(n1046), .B2(mem[461]), .ZN(
        n2224) );
  AOI22_X1 U1729 ( .A1(n1044), .A2(mem[813]), .B1(n1049), .B2(mem[269]), .ZN(
        n2223) );
  AOI22_X1 U1730 ( .A1(n1040), .A2(mem[205]), .B1(n1056), .B2(mem[877]), .ZN(
        n2222) );
  AOI22_X1 U1731 ( .A1(n1054), .A2(mem[333]), .B1(n1461), .B2(mem[749]), .ZN(
        n2221) );
  NAND4_X1 U1732 ( .A1(n2224), .A2(n2223), .A3(n2222), .A4(n2221), .ZN(n2235)
         );
  AOI22_X1 U1733 ( .A1(n1050), .A2(mem[845]), .B1(n1051), .B2(mem[141]), .ZN(
        n2228) );
  AOI22_X1 U1734 ( .A1(n2433), .A2(mem[589]), .B1(n2578), .B2(mem[653]), .ZN(
        n2227) );
  AOI22_X1 U1735 ( .A1(n2750), .A2(mem[525]), .B1(n3010), .B2(mem[557]), .ZN(
        n2226) );
  AOI22_X1 U1736 ( .A1(n1033), .A2(mem[397]), .B1(n1039), .B2(mem[941]), .ZN(
        n2225) );
  NAND4_X1 U1737 ( .A1(n2228), .A2(n2227), .A3(n2226), .A4(n2225), .ZN(n2234)
         );
  AOI22_X1 U1738 ( .A1(n1045), .A2(mem[13]), .B1(n1055), .B2(mem[973]), .ZN(
        n2232) );
  AOI22_X1 U1739 ( .A1(n1745), .A2(mem[621]), .B1(n1053), .B2(mem[429]), .ZN(
        n2231) );
  AOI22_X1 U1740 ( .A1(n1041), .A2(mem[173]), .B1(n1047), .B2(mem[77]), .ZN(
        n2230) );
  AOI22_X1 U1741 ( .A1(n2062), .A2(mem[493]), .B1(n3015), .B2(mem[717]), .ZN(
        n2229) );
  NAND4_X1 U1742 ( .A1(n2232), .A2(n2231), .A3(n2230), .A4(n2229), .ZN(n2233)
         );
  OR4_X1 U1743 ( .A1(n2236), .A2(n2235), .A3(n2234), .A4(n2233), .ZN(
        rdata_c_o[13]) );
  AOI22_X1 U1744 ( .A1(n2832), .A2(mem[429]), .B1(n2841), .B2(mem[717]), .ZN(
        n2240) );
  AOI22_X1 U1745 ( .A1(n2957), .A2(mem[237]), .B1(n2835), .B2(mem[525]), .ZN(
        n2239) );
  AOI22_X1 U1746 ( .A1(n2965), .A2(mem[493]), .B1(n2786), .B2(mem[557]), .ZN(
        n2238) );
  NAND2_X1 U1747 ( .A1(n2968), .A2(mem[909]), .ZN(n2237) );
  NAND4_X1 U1748 ( .A1(n2240), .A2(n2239), .A3(n2238), .A4(n2237), .ZN(n2256)
         );
  AOI22_X1 U1749 ( .A1(n2951), .A2(mem[141]), .B1(n2955), .B2(mem[813]), .ZN(
        n2244) );
  AOI22_X1 U1750 ( .A1(n2989), .A2(mem[973]), .B1(n2765), .B2(mem[589]), .ZN(
        n2243) );
  AOI22_X1 U1751 ( .A1(n2853), .A2(mem[877]), .B1(n1228), .B2(mem[173]), .ZN(
        n2242) );
  AOI22_X1 U1752 ( .A1(n2833), .A2(mem[461]), .B1(n2954), .B2(mem[365]), .ZN(
        n2241) );
  NAND4_X1 U1753 ( .A1(n2244), .A2(n2243), .A3(n2242), .A4(n2241), .ZN(n2255)
         );
  AOI22_X1 U1754 ( .A1(n2850), .A2(mem[685]), .B1(n2851), .B2(mem[397]), .ZN(
        n2248) );
  AOI22_X1 U1755 ( .A1(n2764), .A2(mem[749]), .B1(n2985), .B2(mem[333]), .ZN(
        n2247) );
  AOI22_X1 U1756 ( .A1(n2852), .A2(mem[781]), .B1(n2976), .B2(mem[301]), .ZN(
        n2246) );
  AOI22_X1 U1757 ( .A1(n2775), .A2(mem[45]), .B1(n2966), .B2(mem[77]), .ZN(
        n2245) );
  NAND4_X1 U1758 ( .A1(n2248), .A2(n2247), .A3(n2246), .A4(n2245), .ZN(n2254)
         );
  AOI22_X1 U1759 ( .A1(n2796), .A2(mem[653]), .B1(n2776), .B2(mem[205]), .ZN(
        n2252) );
  AOI22_X1 U1760 ( .A1(n2963), .A2(mem[941]), .B1(n2979), .B2(mem[13]), .ZN(
        n2251) );
  AOI22_X1 U1761 ( .A1(n2770), .A2(mem[621]), .B1(n2848), .B2(mem[269]), .ZN(
        n2250) );
  AOI22_X1 U1762 ( .A1(n2962), .A2(mem[845]), .B1(n2974), .B2(mem[109]), .ZN(
        n2249) );
  NAND4_X1 U1763 ( .A1(n2252), .A2(n2251), .A3(n2250), .A4(n2249), .ZN(n2253)
         );
  OR4_X1 U1764 ( .A1(n2256), .A2(n2255), .A3(n2254), .A4(n2253), .ZN(
        rdata_b_o[13]) );
  INV_X1 U1765 ( .A(wdata_b_i[11]), .ZN(n4430) );
  INV_X1 U1772 ( .A(n2540), .ZN(n2260) );
  NAND3_X1 U1775 ( .A1(n2262), .A2(n2261), .A3(waddr_a_i[2]), .ZN(n2264) );
  AOI22_X1 U1813 ( .A1(n2843), .A2(mem[113]), .B1(n2966), .B2(mem[81]), .ZN(
        n2284) );
  AOI22_X1 U1814 ( .A1(n2850), .A2(mem[689]), .B1(n2835), .B2(mem[529]), .ZN(
        n2283) );
  AOI22_X1 U1815 ( .A1(n2833), .A2(mem[465]), .B1(n2786), .B2(mem[561]), .ZN(
        n2282) );
  NAND2_X1 U1816 ( .A1(n2764), .A2(mem[753]), .ZN(n2281) );
  NAND4_X1 U1817 ( .A1(n2284), .A2(n2283), .A3(n2282), .A4(n2281), .ZN(n2300)
         );
  AOI22_X1 U1818 ( .A1(n2791), .A2(mem[977]), .B1(n2965), .B2(mem[497]), .ZN(
        n2288) );
  AOI22_X1 U1819 ( .A1(n2860), .A2(mem[177]), .B1(n2954), .B2(mem[369]), .ZN(
        n2287) );
  AOI22_X1 U1820 ( .A1(n2770), .A2(mem[625]), .B1(n2775), .B2(mem[49]), .ZN(
        n2286) );
  AOI22_X1 U1821 ( .A1(n2803), .A2(mem[241]), .B1(n2848), .B2(mem[273]), .ZN(
        n2285) );
  NAND4_X1 U1822 ( .A1(n2288), .A2(n2287), .A3(n2286), .A4(n2285), .ZN(n2299)
         );
  AOI22_X1 U1823 ( .A1(n2796), .A2(mem[657]), .B1(n2979), .B2(mem[17]), .ZN(
        n2292) );
  AOI22_X1 U1824 ( .A1(n2992), .A2(mem[881]), .B1(n2977), .B2(mem[209]), .ZN(
        n2291) );
  AOI22_X1 U1825 ( .A1(n2859), .A2(mem[145]), .B1(n2953), .B2(mem[721]), .ZN(
        n2290) );
  AOI22_X1 U1826 ( .A1(n2963), .A2(mem[945]), .B1(n2858), .B2(mem[305]), .ZN(
        n2289) );
  NAND4_X1 U1827 ( .A1(n2292), .A2(n2291), .A3(n2290), .A4(n2289), .ZN(n2298)
         );
  AOI22_X1 U1828 ( .A1(n2968), .A2(mem[913]), .B1(n2986), .B2(mem[593]), .ZN(
        n2296) );
  AOI22_X1 U1829 ( .A1(n2759), .A2(mem[337]), .B1(n2832), .B2(mem[433]), .ZN(
        n2295) );
  AOI22_X1 U1830 ( .A1(n2639), .A2(mem[849]), .B1(n2987), .B2(mem[401]), .ZN(
        n2294) );
  AOI22_X1 U1831 ( .A1(n2975), .A2(mem[785]), .B1(n2840), .B2(mem[817]), .ZN(
        n2293) );
  NAND4_X1 U1832 ( .A1(n2296), .A2(n2295), .A3(n2294), .A4(n2293), .ZN(n2297)
         );
  OR4_X1 U1833 ( .A1(n2300), .A2(n2299), .A3(n2298), .A4(n2297), .ZN(
        rdata_b_o[17]) );
  AOI22_X1 U1834 ( .A1(n1050), .A2(mem[849]), .B1(n1395), .B2(mem[305]), .ZN(
        n2304) );
  AOI22_X1 U1835 ( .A1(n2668), .A2(mem[625]), .B1(n2578), .B2(mem[657]), .ZN(
        n2303) );
  AOI22_X1 U1836 ( .A1(n2750), .A2(mem[529]), .B1(n1051), .B2(mem[145]), .ZN(
        n2302) );
  NAND2_X1 U1837 ( .A1(n1053), .A2(mem[433]), .ZN(n2301) );
  NAND4_X1 U1838 ( .A1(n2304), .A2(n2303), .A3(n2302), .A4(n2301), .ZN(n2320)
         );
  AOI22_X1 U1839 ( .A1(n1033), .A2(mem[401]), .B1(n1040), .B2(mem[209]), .ZN(
        n2308) );
  AOI22_X1 U1840 ( .A1(n1055), .A2(mem[977]), .B1(n1039), .B2(mem[945]), .ZN(
        n2307) );
  AOI22_X1 U1841 ( .A1(n1054), .A2(mem[337]), .B1(n3010), .B2(mem[561]), .ZN(
        n2306) );
  AOI22_X1 U1842 ( .A1(n2433), .A2(mem[593]), .B1(n1415), .B2(mem[881]), .ZN(
        n2305) );
  NAND4_X1 U1843 ( .A1(n2308), .A2(n2307), .A3(n2306), .A4(n2305), .ZN(n2319)
         );
  AOI22_X1 U1844 ( .A1(n1740), .A2(mem[497]), .B1(n1044), .B2(mem[817]), .ZN(
        n2312) );
  AOI22_X1 U1845 ( .A1(n2705), .A2(mem[753]), .B1(n1047), .B2(mem[81]), .ZN(
        n2311) );
  AOI22_X1 U1846 ( .A1(n1048), .A2(mem[785]), .B1(n1049), .B2(mem[273]), .ZN(
        n2310) );
  AOI22_X1 U1847 ( .A1(n1041), .A2(mem[177]), .B1(n1042), .B2(mem[241]), .ZN(
        n2309) );
  NAND4_X1 U1848 ( .A1(n2312), .A2(n2311), .A3(n2310), .A4(n2309), .ZN(n2318)
         );
  AOI22_X1 U1849 ( .A1(n2869), .A2(mem[913]), .B1(n1052), .B2(mem[689]), .ZN(
        n2316) );
  AOI22_X1 U1850 ( .A1(n3001), .A2(mem[49]), .B1(n1043), .B2(mem[113]), .ZN(
        n2315) );
  AOI22_X1 U1851 ( .A1(n3015), .A2(mem[721]), .B1(n1046), .B2(mem[465]), .ZN(
        n2314) );
  AOI22_X1 U1852 ( .A1(n1045), .A2(mem[17]), .B1(n2874), .B2(mem[369]), .ZN(
        n2313) );
  NAND4_X1 U1853 ( .A1(n2316), .A2(n2315), .A3(n2314), .A4(n2313), .ZN(n2317)
         );
  OR4_X1 U1854 ( .A1(n2320), .A2(n2319), .A3(n2318), .A4(n2317), .ZN(
        rdata_c_o[17]) );
  AOI22_X1 U1855 ( .A1(n2963), .A2(mem[947]), .B1(n2957), .B2(mem[243]), .ZN(
        n2324) );
  AOI22_X1 U1856 ( .A1(n2967), .A2(mem[659]), .B1(n2841), .B2(mem[723]), .ZN(
        n2323) );
  AOI22_X1 U1857 ( .A1(n2965), .A2(mem[499]), .B1(n2851), .B2(mem[403]), .ZN(
        n2322) );
  NAND2_X1 U1858 ( .A1(n2850), .A2(mem[691]), .ZN(n2321) );
  NAND4_X1 U1859 ( .A1(n2324), .A2(n2323), .A3(n2322), .A4(n2321), .ZN(n2340)
         );
  AOI22_X1 U1860 ( .A1(n2764), .A2(mem[755]), .B1(n2976), .B2(mem[307]), .ZN(
        n2328) );
  AOI22_X1 U1861 ( .A1(n2785), .A2(mem[915]), .B1(n2765), .B2(mem[595]), .ZN(
        n2327) );
  AOI22_X1 U1862 ( .A1(n2966), .A2(mem[83]), .B1(n2835), .B2(mem[531]), .ZN(
        n2326) );
  AOI22_X1 U1863 ( .A1(n2853), .A2(mem[883]), .B1(n2955), .B2(mem[819]), .ZN(
        n2325) );
  NAND4_X1 U1864 ( .A1(n2328), .A2(n2327), .A3(n2326), .A4(n2325), .ZN(n2339)
         );
  AOI22_X1 U1865 ( .A1(n2791), .A2(mem[979]), .B1(n2964), .B2(mem[435]), .ZN(
        n2332) );
  AOI22_X1 U1866 ( .A1(n2975), .A2(mem[787]), .B1(n2951), .B2(mem[147]), .ZN(
        n2331) );
  AOI22_X1 U1867 ( .A1(n2956), .A2(mem[627]), .B1(n2776), .B2(mem[211]), .ZN(
        n2330) );
  AOI22_X1 U1868 ( .A1(n2985), .A2(mem[339]), .B1(n1228), .B2(mem[179]), .ZN(
        n2329) );
  NAND4_X1 U1869 ( .A1(n2332), .A2(n2331), .A3(n2330), .A4(n2329), .ZN(n2338)
         );
  AOI22_X1 U1870 ( .A1(n2954), .A2(mem[371]), .B1(n2979), .B2(mem[19]), .ZN(
        n2336) );
  AOI22_X1 U1871 ( .A1(n2974), .A2(mem[115]), .B1(n2848), .B2(mem[275]), .ZN(
        n2335) );
  AOI22_X1 U1872 ( .A1(n2775), .A2(mem[51]), .B1(n2991), .B2(mem[563]), .ZN(
        n2334) );
  AOI22_X1 U1873 ( .A1(n2952), .A2(mem[467]), .B1(n2962), .B2(mem[851]), .ZN(
        n2333) );
  NAND4_X1 U1874 ( .A1(n2336), .A2(n2335), .A3(n2334), .A4(n2333), .ZN(n2337)
         );
  OR4_X1 U1875 ( .A1(n2340), .A2(n2339), .A3(n2338), .A4(n2337), .ZN(
        rdata_b_o[19]) );
  AOI22_X1 U1876 ( .A1(n1033), .A2(mem[403]), .B1(n1049), .B2(mem[275]), .ZN(
        n2344) );
  AOI22_X1 U1877 ( .A1(n2869), .A2(mem[915]), .B1(n1048), .B2(mem[787]), .ZN(
        n2343) );
  AOI22_X1 U1878 ( .A1(n1053), .A2(mem[435]), .B1(n3010), .B2(mem[563]), .ZN(
        n2342) );
  NAND2_X1 U1879 ( .A1(n1051), .A2(mem[147]), .ZN(n2341) );
  NAND4_X1 U1880 ( .A1(n2344), .A2(n2343), .A3(n2342), .A4(n2341), .ZN(n2360)
         );
  AOI22_X1 U1881 ( .A1(n1751), .A2(mem[19]), .B1(n1043), .B2(mem[115]), .ZN(
        n2348) );
  AOI22_X1 U1882 ( .A1(n1055), .A2(mem[979]), .B1(n1047), .B2(mem[83]), .ZN(
        n2347) );
  AOI22_X1 U1883 ( .A1(n3001), .A2(mem[51]), .B1(n1040), .B2(mem[211]), .ZN(
        n2346) );
  AOI22_X1 U1884 ( .A1(n1039), .A2(mem[947]), .B1(n1046), .B2(mem[467]), .ZN(
        n2345) );
  NAND4_X1 U1885 ( .A1(n2348), .A2(n2347), .A3(n2346), .A4(n2345), .ZN(n2359)
         );
  AOI22_X1 U1886 ( .A1(n3016), .A2(mem[307]), .B1(n3015), .B2(mem[723]), .ZN(
        n2352) );
  AOI22_X1 U1887 ( .A1(n2062), .A2(mem[499]), .B1(n1052), .B2(mem[691]), .ZN(
        n2351) );
  AOI22_X1 U1888 ( .A1(n1050), .A2(mem[851]), .B1(n1056), .B2(mem[883]), .ZN(
        n2350) );
  AOI22_X1 U1889 ( .A1(n1745), .A2(mem[627]), .B1(n2874), .B2(mem[371]), .ZN(
        n2349) );
  NAND4_X1 U1890 ( .A1(n2352), .A2(n2351), .A3(n2350), .A4(n2349), .ZN(n2358)
         );
  AOI22_X1 U1891 ( .A1(n1042), .A2(mem[243]), .B1(n1054), .B2(mem[339]), .ZN(
        n2356) );
  AOI22_X1 U1892 ( .A1(n1041), .A2(mem[179]), .B1(n1461), .B2(mem[755]), .ZN(
        n2355) );
  AOI22_X1 U1893 ( .A1(n2433), .A2(mem[595]), .B1(n2578), .B2(mem[659]), .ZN(
        n2354) );
  AOI22_X1 U1894 ( .A1(n2750), .A2(mem[531]), .B1(n1044), .B2(mem[819]), .ZN(
        n2353) );
  NAND4_X1 U1895 ( .A1(n2356), .A2(n2355), .A3(n2354), .A4(n2353), .ZN(n2357)
         );
  OR4_X1 U1896 ( .A1(n2360), .A2(n2359), .A3(n2358), .A4(n2357), .ZN(
        rdata_c_o[19]) );
  AOI22_X1 U1897 ( .A1(n2803), .A2(mem[247]), .B1(n2841), .B2(mem[727]), .ZN(
        n2364) );
  AOI22_X1 U1898 ( .A1(n2965), .A2(mem[503]), .B1(n2964), .B2(mem[439]), .ZN(
        n2363) );
  AOI22_X1 U1899 ( .A1(n2956), .A2(mem[631]), .B1(n2986), .B2(mem[599]), .ZN(
        n2362) );
  NAND2_X1 U1900 ( .A1(n2985), .A2(mem[343]), .ZN(n2361) );
  NAND4_X1 U1901 ( .A1(n2364), .A2(n2363), .A3(n2362), .A4(n2361), .ZN(n2380)
         );
  AOI22_X1 U1902 ( .A1(n2850), .A2(mem[695]), .B1(n2785), .B2(mem[919]), .ZN(
        n2368) );
  AOI22_X1 U1903 ( .A1(n2853), .A2(mem[887]), .B1(n2852), .B2(mem[791]), .ZN(
        n2367) );
  AOI22_X1 U1904 ( .A1(n2775), .A2(mem[55]), .B1(n2991), .B2(mem[567]), .ZN(
        n2366) );
  AOI22_X1 U1905 ( .A1(n2764), .A2(mem[759]), .B1(n2833), .B2(mem[471]), .ZN(
        n2365) );
  NAND4_X1 U1906 ( .A1(n2368), .A2(n2367), .A3(n2366), .A4(n2365), .ZN(n2379)
         );
  AOI22_X1 U1907 ( .A1(n2951), .A2(mem[151]), .B1(n2976), .B2(mem[311]), .ZN(
        n2372) );
  AOI22_X1 U1908 ( .A1(n2840), .A2(mem[823]), .B1(n2851), .B2(mem[407]), .ZN(
        n2371) );
  AOI22_X1 U1909 ( .A1(n2966), .A2(mem[87]), .B1(n2977), .B2(mem[215]), .ZN(
        n2370) );
  AOI22_X1 U1910 ( .A1(n2639), .A2(mem[855]), .B1(n2989), .B2(mem[983]), .ZN(
        n2369) );
  NAND4_X1 U1911 ( .A1(n2372), .A2(n2371), .A3(n2370), .A4(n2369), .ZN(n2378)
         );
  AOI22_X1 U1912 ( .A1(n2797), .A2(mem[951]), .B1(n1228), .B2(mem[183]), .ZN(
        n2376) );
  AOI22_X1 U1913 ( .A1(n2796), .A2(mem[663]), .B1(n2842), .B2(mem[375]), .ZN(
        n2375) );
  AOI22_X1 U1914 ( .A1(n2988), .A2(mem[535]), .B1(n2834), .B2(mem[23]), .ZN(
        n2374) );
  AOI22_X1 U1915 ( .A1(n2974), .A2(mem[119]), .B1(n2848), .B2(mem[279]), .ZN(
        n2373) );
  NAND4_X1 U1916 ( .A1(n2376), .A2(n2375), .A3(n2374), .A4(n2373), .ZN(n2377)
         );
  OR4_X1 U1917 ( .A1(n2380), .A2(n2379), .A3(n2378), .A4(n2377), .ZN(
        rdata_b_o[23]) );
  AOI22_X1 U1918 ( .A1(n2874), .A2(mem[375]), .B1(n1053), .B2(mem[439]), .ZN(
        n2384) );
  AOI22_X1 U1919 ( .A1(n2668), .A2(mem[631]), .B1(n1041), .B2(mem[183]), .ZN(
        n2383) );
  AOI22_X1 U1920 ( .A1(n1039), .A2(mem[951]), .B1(n1049), .B2(mem[279]), .ZN(
        n2382) );
  NAND2_X1 U1921 ( .A1(n2578), .A2(mem[663]), .ZN(n2381) );
  NAND4_X1 U1922 ( .A1(n2384), .A2(n2383), .A3(n2382), .A4(n2381), .ZN(n2400)
         );
  AOI22_X1 U1923 ( .A1(n1752), .A2(mem[599]), .B1(n1048), .B2(mem[791]), .ZN(
        n2388) );
  AOI22_X1 U1924 ( .A1(n1033), .A2(mem[407]), .B1(n2705), .B2(mem[759]), .ZN(
        n2387) );
  AOI22_X1 U1925 ( .A1(n3001), .A2(mem[55]), .B1(n3010), .B2(mem[567]), .ZN(
        n2386) );
  AOI22_X1 U1926 ( .A1(n1042), .A2(mem[247]), .B1(n1043), .B2(mem[119]), .ZN(
        n2385) );
  NAND4_X1 U1927 ( .A1(n2388), .A2(n2387), .A3(n2386), .A4(n2385), .ZN(n2399)
         );
  AOI22_X1 U1928 ( .A1(n1055), .A2(mem[983]), .B1(n1044), .B2(mem[823]), .ZN(
        n2392) );
  AOI22_X1 U1929 ( .A1(n2062), .A2(mem[503]), .B1(n1395), .B2(mem[311]), .ZN(
        n2391) );
  AOI22_X1 U1930 ( .A1(n1403), .A2(mem[919]), .B1(n1054), .B2(mem[343]), .ZN(
        n2390) );
  AOI22_X1 U1931 ( .A1(n1050), .A2(mem[855]), .B1(n1045), .B2(mem[23]), .ZN(
        n2389) );
  NAND4_X1 U1932 ( .A1(n2392), .A2(n2391), .A3(n2390), .A4(n2389), .ZN(n2398)
         );
  AOI22_X1 U1933 ( .A1(n2750), .A2(mem[535]), .B1(n1046), .B2(mem[471]), .ZN(
        n2396) );
  AOI22_X1 U1934 ( .A1(n1052), .A2(mem[695]), .B1(n1051), .B2(mem[151]), .ZN(
        n2395) );
  AOI22_X1 U1935 ( .A1(n1040), .A2(mem[215]), .B1(n1047), .B2(mem[87]), .ZN(
        n2394) );
  AOI22_X1 U1936 ( .A1(n1452), .A2(mem[727]), .B1(n1056), .B2(mem[887]), .ZN(
        n2393) );
  NAND4_X1 U1937 ( .A1(n2396), .A2(n2395), .A3(n2394), .A4(n2393), .ZN(n2397)
         );
  OR4_X1 U1938 ( .A1(n2400), .A2(n2399), .A3(n2398), .A4(n2397), .ZN(
        rdata_c_o[23]) );
  AOI22_X1 U1939 ( .A1(n2853), .A2(mem[888]), .B1(n2951), .B2(mem[152]), .ZN(
        n2404) );
  AOI22_X1 U1940 ( .A1(n2843), .A2(mem[120]), .B1(n2834), .B2(mem[24]), .ZN(
        n2403) );
  AOI22_X1 U1941 ( .A1(n2963), .A2(mem[952]), .B1(n2976), .B2(mem[312]), .ZN(
        n2402) );
  NAND2_X1 U1942 ( .A1(n2852), .A2(mem[792]), .ZN(n2401) );
  NAND4_X1 U1943 ( .A1(n2404), .A2(n2403), .A3(n2402), .A4(n2401), .ZN(n2420)
         );
  AOI22_X1 U1944 ( .A1(n2833), .A2(mem[472]), .B1(n2953), .B2(mem[728]), .ZN(
        n2408) );
  AOI22_X1 U1945 ( .A1(n2967), .A2(mem[664]), .B1(n2965), .B2(mem[504]), .ZN(
        n2407) );
  AOI22_X1 U1946 ( .A1(n2770), .A2(mem[632]), .B1(n2985), .B2(mem[344]), .ZN(
        n2406) );
  AOI22_X1 U1947 ( .A1(n2989), .A2(mem[984]), .B1(n2954), .B2(mem[376]), .ZN(
        n2405) );
  NAND4_X1 U1948 ( .A1(n2408), .A2(n2407), .A3(n2406), .A4(n2405), .ZN(n2419)
         );
  AOI22_X1 U1949 ( .A1(n2968), .A2(mem[920]), .B1(n2765), .B2(mem[600]), .ZN(
        n2412) );
  AOI22_X1 U1950 ( .A1(n2764), .A2(mem[760]), .B1(n2639), .B2(mem[856]), .ZN(
        n2411) );
  AOI22_X1 U1951 ( .A1(n2775), .A2(mem[56]), .B1(n2848), .B2(mem[280]), .ZN(
        n2410) );
  AOI22_X1 U1952 ( .A1(n2969), .A2(mem[696]), .B1(n2860), .B2(mem[184]), .ZN(
        n2409) );
  NAND4_X1 U1953 ( .A1(n2412), .A2(n2411), .A3(n2410), .A4(n2409), .ZN(n2418)
         );
  AOI22_X1 U1954 ( .A1(n2957), .A2(mem[248]), .B1(n2991), .B2(mem[568]), .ZN(
        n2416) );
  AOI22_X1 U1955 ( .A1(n2798), .A2(mem[88]), .B1(n2840), .B2(mem[824]), .ZN(
        n2415) );
  AOI22_X1 U1956 ( .A1(n2977), .A2(mem[216]), .B1(n2988), .B2(mem[536]), .ZN(
        n2414) );
  AOI22_X1 U1957 ( .A1(n2832), .A2(mem[440]), .B1(n2987), .B2(mem[408]), .ZN(
        n2413) );
  NAND4_X1 U1958 ( .A1(n2416), .A2(n2415), .A3(n2414), .A4(n2413), .ZN(n2417)
         );
  OR4_X1 U1959 ( .A1(n2420), .A2(n2419), .A3(n2418), .A4(n2417), .ZN(
        rdata_b_o[24]) );
  AOI22_X1 U1960 ( .A1(n3015), .A2(mem[728]), .B1(n1049), .B2(mem[280]), .ZN(
        n2424) );
  AOI22_X1 U1961 ( .A1(n2874), .A2(mem[376]), .B1(n1047), .B2(mem[88]), .ZN(
        n2423) );
  AOI22_X1 U1962 ( .A1(n1055), .A2(mem[984]), .B1(n2705), .B2(mem[760]), .ZN(
        n2422) );
  NAND2_X1 U1963 ( .A1(n1053), .A2(mem[440]), .ZN(n2421) );
  NAND4_X1 U1964 ( .A1(n2424), .A2(n2423), .A3(n2422), .A4(n2421), .ZN(n2441)
         );
  AOI22_X1 U1965 ( .A1(n2578), .A2(mem[664]), .B1(n1052), .B2(mem[696]), .ZN(
        n2428) );
  AOI22_X1 U1966 ( .A1(n1751), .A2(mem[24]), .B1(n1041), .B2(mem[184]), .ZN(
        n2427) );
  AOI22_X1 U1967 ( .A1(n2869), .A2(mem[920]), .B1(n1040), .B2(mem[216]), .ZN(
        n2426) );
  AOI22_X1 U1968 ( .A1(n1050), .A2(mem[856]), .B1(n1042), .B2(mem[248]), .ZN(
        n2425) );
  NAND4_X1 U1969 ( .A1(n2428), .A2(n2427), .A3(n2426), .A4(n2425), .ZN(n2440)
         );
  AOI22_X1 U1970 ( .A1(n1043), .A2(mem[120]), .B1(n1056), .B2(mem[888]), .ZN(
        n2432) );
  AOI22_X1 U1971 ( .A1(n1039), .A2(mem[952]), .B1(n3010), .B2(mem[568]), .ZN(
        n2431) );
  AOI22_X1 U1972 ( .A1(n2062), .A2(mem[504]), .B1(n2750), .B2(mem[536]), .ZN(
        n2430) );
  AOI22_X1 U1973 ( .A1(n3001), .A2(mem[56]), .B1(n1033), .B2(mem[408]), .ZN(
        n2429) );
  NAND4_X1 U1974 ( .A1(n2432), .A2(n2431), .A3(n2430), .A4(n2429), .ZN(n2439)
         );
  AOI22_X1 U1975 ( .A1(n1745), .A2(mem[632]), .B1(n2433), .B2(mem[600]), .ZN(
        n2437) );
  AOI22_X1 U1976 ( .A1(n1054), .A2(mem[344]), .B1(n1046), .B2(mem[472]), .ZN(
        n2436) );
  AOI22_X1 U1977 ( .A1(n3016), .A2(mem[312]), .B1(n1048), .B2(mem[792]), .ZN(
        n2435) );
  AOI22_X1 U1978 ( .A1(n1044), .A2(mem[824]), .B1(n1051), .B2(mem[152]), .ZN(
        n2434) );
  NAND4_X1 U1979 ( .A1(n2437), .A2(n2436), .A3(n2435), .A4(n2434), .ZN(n2438)
         );
  OR4_X1 U1980 ( .A1(n2441), .A2(n2440), .A3(n2439), .A4(n2438), .ZN(
        rdata_c_o[24]) );
  INV_X1 U1981 ( .A(wdata_b_i[8]), .ZN(n4424) );
  NAND3_X1 U2035 ( .A1(n2468), .A2(n3768), .A3(waddr_b_i[1]), .ZN(n2546) );
  NOR2_X1 U2037 ( .A1(n2525), .A2(n2527), .ZN(n2548) );
  NAND3_X1 U2038 ( .A1(n2548), .A2(n2473), .A3(n2533), .ZN(n2469) );
  NAND3_X1 U2045 ( .A1(n2548), .A2(waddr_a_i[2]), .A3(n2473), .ZN(n2474) );
  NAND2_X1 U2051 ( .A1(n2478), .A2(n3768), .ZN(n2539) );
  NOR2_X1 U2053 ( .A1(n2525), .A2(n2480), .ZN(n2541) );
  NAND2_X1 U2054 ( .A1(n2541), .A2(n2533), .ZN(n2481) );
  AOI22_X1 U2060 ( .A1(n2869), .A2(mem[906]), .B1(n1047), .B2(mem[74]), .ZN(
        n2488) );
  AOI22_X1 U2061 ( .A1(n2062), .A2(mem[490]), .B1(n2578), .B2(mem[650]), .ZN(
        n2487) );
  AOI22_X1 U2062 ( .A1(n1045), .A2(mem[10]), .B1(n1395), .B2(mem[298]), .ZN(
        n2486) );
  NAND2_X1 U2063 ( .A1(n1051), .A2(mem[138]), .ZN(n2485) );
  NAND4_X1 U2064 ( .A1(n2488), .A2(n2487), .A3(n2486), .A4(n2485), .ZN(n2504)
         );
  AOI22_X1 U2065 ( .A1(n2668), .A2(mem[618]), .B1(n1049), .B2(mem[266]), .ZN(
        n2492) );
  AOI22_X1 U2066 ( .A1(n3001), .A2(mem[42]), .B1(n3010), .B2(mem[554]), .ZN(
        n2491) );
  AOI22_X1 U2067 ( .A1(n1039), .A2(mem[938]), .B1(n1041), .B2(mem[170]), .ZN(
        n2490) );
  AOI22_X1 U2068 ( .A1(n1033), .A2(mem[394]), .B1(n1052), .B2(mem[682]), .ZN(
        n2489) );
  NAND4_X1 U2069 ( .A1(n2492), .A2(n2491), .A3(n2490), .A4(n2489), .ZN(n2503)
         );
  AOI22_X1 U2070 ( .A1(n1050), .A2(mem[842]), .B1(n1054), .B2(mem[330]), .ZN(
        n2496) );
  AOI22_X1 U2071 ( .A1(n1424), .A2(mem[362]), .B1(n1040), .B2(mem[202]), .ZN(
        n2495) );
  AOI22_X1 U2072 ( .A1(n1752), .A2(mem[586]), .B1(n3015), .B2(mem[714]), .ZN(
        n2494) );
  AOI22_X1 U2073 ( .A1(n2705), .A2(mem[746]), .B1(n1048), .B2(mem[778]), .ZN(
        n2493) );
  NAND4_X1 U2074 ( .A1(n2496), .A2(n2495), .A3(n2494), .A4(n2493), .ZN(n2502)
         );
  AOI22_X1 U2075 ( .A1(n1055), .A2(mem[970]), .B1(n1056), .B2(mem[874]), .ZN(
        n2500) );
  AOI22_X1 U2076 ( .A1(n1042), .A2(mem[234]), .B1(n1046), .B2(mem[458]), .ZN(
        n2499) );
  AOI22_X1 U2077 ( .A1(n1044), .A2(mem[810]), .B1(n1043), .B2(mem[106]), .ZN(
        n2498) );
  AOI22_X1 U2078 ( .A1(n1053), .A2(mem[426]), .B1(n2750), .B2(mem[522]), .ZN(
        n2497) );
  NAND4_X1 U2079 ( .A1(n2500), .A2(n2499), .A3(n2498), .A4(n2497), .ZN(n2501)
         );
  OR4_X1 U2080 ( .A1(n2504), .A2(n2503), .A3(n2502), .A4(n2501), .ZN(
        rdata_c_o[10]) );
  AOI22_X1 U2081 ( .A1(n2852), .A2(mem[778]), .B1(n2835), .B2(mem[522]), .ZN(
        n2508) );
  AOI22_X1 U2082 ( .A1(n2803), .A2(mem[234]), .B1(n2978), .B2(mem[266]), .ZN(
        n2507) );
  AOI22_X1 U2083 ( .A1(n2989), .A2(mem[970]), .B1(n2977), .B2(mem[202]), .ZN(
        n2506) );
  NAND2_X1 U2084 ( .A1(n2796), .A2(mem[650]), .ZN(n2505) );
  NAND4_X1 U2085 ( .A1(n2508), .A2(n2507), .A3(n2506), .A4(n2505), .ZN(n2524)
         );
  AOI22_X1 U2086 ( .A1(n2843), .A2(mem[106]), .B1(n2955), .B2(mem[810]), .ZN(
        n2512) );
  AOI22_X1 U2087 ( .A1(n2962), .A2(mem[842]), .B1(n2841), .B2(mem[714]), .ZN(
        n2511) );
  AOI22_X1 U2088 ( .A1(n2963), .A2(mem[938]), .B1(n2860), .B2(mem[170]), .ZN(
        n2510) );
  AOI22_X1 U2089 ( .A1(n2853), .A2(mem[874]), .B1(n2770), .B2(mem[618]), .ZN(
        n2509) );
  NAND4_X1 U2090 ( .A1(n2512), .A2(n2511), .A3(n2510), .A4(n2509), .ZN(n2523)
         );
  AOI22_X1 U2091 ( .A1(n2966), .A2(mem[74]), .B1(n2954), .B2(mem[362]), .ZN(
        n2516) );
  AOI22_X1 U2092 ( .A1(n2951), .A2(mem[138]), .B1(n2786), .B2(mem[554]), .ZN(
        n2515) );
  AOI22_X1 U2093 ( .A1(n2765), .A2(mem[586]), .B1(n2979), .B2(mem[10]), .ZN(
        n2514) );
  AOI22_X1 U2094 ( .A1(n2850), .A2(mem[682]), .B1(n2851), .B2(mem[394]), .ZN(
        n2513) );
  NAND4_X1 U2095 ( .A1(n2516), .A2(n2515), .A3(n2514), .A4(n2513), .ZN(n2522)
         );
  AOI22_X1 U2096 ( .A1(n2764), .A2(mem[746]), .B1(n2832), .B2(mem[426]), .ZN(
        n2520) );
  AOI22_X1 U2097 ( .A1(n2968), .A2(mem[906]), .B1(n2976), .B2(mem[298]), .ZN(
        n2519) );
  AOI22_X1 U2098 ( .A1(n2759), .A2(mem[330]), .B1(n2965), .B2(mem[490]), .ZN(
        n2518) );
  AOI22_X1 U2099 ( .A1(n2833), .A2(mem[458]), .B1(n2775), .B2(mem[42]), .ZN(
        n2517) );
  NAND4_X1 U2100 ( .A1(n2520), .A2(n2519), .A3(n2518), .A4(n2517), .ZN(n2521)
         );
  OR4_X1 U2101 ( .A1(n2524), .A2(n2523), .A3(n2522), .A4(n2521), .ZN(
        rdata_b_o[10]) );
  INV_X1 U2103 ( .A(n2525), .ZN(n2526) );
  AND3_X1 U2104 ( .A1(n2549), .A2(n2527), .A3(n2526), .ZN(n2530) );
  INV_X1 U2105 ( .A(n2530), .ZN(n2528) );
  INV_X1 U2111 ( .A(n2532), .ZN(n2534) );
  NAND3_X1 U2112 ( .A1(n2534), .A2(n2548), .A3(n2533), .ZN(n2535) );
  NAND2_X1 U2119 ( .A1(n2541), .A2(waddr_a_i[2]), .ZN(n2542) );
  AND2_X1 U2126 ( .A1(n2549), .A2(n2548), .ZN(n2551) );
  INV_X1 U2127 ( .A(n2551), .ZN(n2550) );
  AOI22_X1 U2132 ( .A1(n2850), .A2(mem[694]), .B1(n2841), .B2(mem[726]), .ZN(
        n2557) );
  AOI22_X1 U2133 ( .A1(n2977), .A2(mem[214]), .B1(n2786), .B2(mem[566]), .ZN(
        n2556) );
  AOI22_X1 U2134 ( .A1(n2848), .A2(mem[278]), .B1(n2955), .B2(mem[822]), .ZN(
        n2555) );
  NAND2_X1 U2135 ( .A1(n2954), .A2(mem[374]), .ZN(n2554) );
  NAND4_X1 U2136 ( .A1(n2557), .A2(n2556), .A3(n2555), .A4(n2554), .ZN(n2573)
         );
  AOI22_X1 U2137 ( .A1(n2770), .A2(mem[630]), .B1(n2962), .B2(mem[854]), .ZN(
        n2561) );
  AOI22_X1 U2138 ( .A1(n2967), .A2(mem[662]), .B1(n2860), .B2(mem[182]), .ZN(
        n2560) );
  AOI22_X1 U2139 ( .A1(n2968), .A2(mem[918]), .B1(n2976), .B2(mem[310]), .ZN(
        n2559) );
  AOI22_X1 U2140 ( .A1(n2853), .A2(mem[886]), .B1(n2957), .B2(mem[246]), .ZN(
        n2558) );
  NAND4_X1 U2141 ( .A1(n2561), .A2(n2560), .A3(n2559), .A4(n2558), .ZN(n2572)
         );
  AOI22_X1 U2142 ( .A1(n2985), .A2(mem[342]), .B1(n2966), .B2(mem[86]), .ZN(
        n2565) );
  AOI22_X1 U2143 ( .A1(n2975), .A2(mem[790]), .B1(n2832), .B2(mem[438]), .ZN(
        n2564) );
  AOI22_X1 U2144 ( .A1(n2797), .A2(mem[950]), .B1(n2989), .B2(mem[982]), .ZN(
        n2563) );
  AOI22_X1 U2145 ( .A1(n2952), .A2(mem[470]), .B1(n2974), .B2(mem[118]), .ZN(
        n2562) );
  NAND4_X1 U2146 ( .A1(n2565), .A2(n2564), .A3(n2563), .A4(n2562), .ZN(n2571)
         );
  AOI22_X1 U2147 ( .A1(n2965), .A2(mem[502]), .B1(n2979), .B2(mem[22]), .ZN(
        n2569) );
  AOI22_X1 U2148 ( .A1(n2765), .A2(mem[598]), .B1(n2835), .B2(mem[534]), .ZN(
        n2568) );
  AOI22_X1 U2149 ( .A1(n2980), .A2(mem[758]), .B1(n2775), .B2(mem[54]), .ZN(
        n2567) );
  AOI22_X1 U2150 ( .A1(n2951), .A2(mem[150]), .B1(n2987), .B2(mem[406]), .ZN(
        n2566) );
  NAND4_X1 U2151 ( .A1(n2569), .A2(n2568), .A3(n2567), .A4(n2566), .ZN(n2570)
         );
  OR4_X1 U2152 ( .A1(n2573), .A2(n2572), .A3(n2571), .A4(n2570), .ZN(
        rdata_b_o[22]) );
  AOI22_X1 U2153 ( .A1(n1033), .A2(mem[406]), .B1(n2750), .B2(mem[534]), .ZN(
        n2577) );
  AOI22_X1 U2154 ( .A1(n1054), .A2(mem[342]), .B1(n1043), .B2(mem[118]), .ZN(
        n2576) );
  AOI22_X1 U2155 ( .A1(n1052), .A2(mem[694]), .B1(n1044), .B2(mem[822]), .ZN(
        n2575) );
  NAND2_X1 U2156 ( .A1(n1042), .A2(mem[246]), .ZN(n2574) );
  NAND4_X1 U2157 ( .A1(n2577), .A2(n2576), .A3(n2575), .A4(n2574), .ZN(n2594)
         );
  AOI22_X1 U2158 ( .A1(n1752), .A2(mem[598]), .B1(n3015), .B2(mem[726]), .ZN(
        n2582) );
  AOI22_X1 U2159 ( .A1(n1055), .A2(mem[982]), .B1(n1046), .B2(mem[470]), .ZN(
        n2581) );
  AOI22_X1 U2160 ( .A1(n1039), .A2(mem[950]), .B1(n1049), .B2(mem[278]), .ZN(
        n2580) );
  AOI22_X1 U2161 ( .A1(n3001), .A2(mem[54]), .B1(n2578), .B2(mem[662]), .ZN(
        n2579) );
  NAND4_X1 U2162 ( .A1(n2582), .A2(n2581), .A3(n2580), .A4(n2579), .ZN(n2593)
         );
  AOI22_X1 U2163 ( .A1(n2062), .A2(mem[502]), .B1(n1403), .B2(mem[918]), .ZN(
        n2586) );
  AOI22_X1 U2164 ( .A1(n1045), .A2(mem[22]), .B1(n1047), .B2(mem[86]), .ZN(
        n2585) );
  AOI22_X1 U2165 ( .A1(n1040), .A2(mem[214]), .B1(n1048), .B2(mem[790]), .ZN(
        n2584) );
  AOI22_X1 U2166 ( .A1(n1050), .A2(mem[854]), .B1(n1041), .B2(mem[182]), .ZN(
        n2583) );
  NAND4_X1 U2167 ( .A1(n2586), .A2(n2585), .A3(n2584), .A4(n2583), .ZN(n2592)
         );
  AOI22_X1 U2168 ( .A1(n3016), .A2(mem[310]), .B1(n1056), .B2(mem[886]), .ZN(
        n2590) );
  AOI22_X1 U2169 ( .A1(n1745), .A2(mem[630]), .B1(n3010), .B2(mem[566]), .ZN(
        n2589) );
  AOI22_X1 U2170 ( .A1(n2874), .A2(mem[374]), .B1(n1051), .B2(mem[150]), .ZN(
        n2588) );
  AOI22_X1 U2171 ( .A1(n1053), .A2(mem[438]), .B1(n1461), .B2(mem[758]), .ZN(
        n2587) );
  NAND4_X1 U2172 ( .A1(n2590), .A2(n2589), .A3(n2588), .A4(n2587), .ZN(n2591)
         );
  OR4_X1 U2173 ( .A1(n2594), .A2(n2593), .A3(n2592), .A4(n2591), .ZN(
        rdata_c_o[22]) );
  AOI22_X1 U2174 ( .A1(n1033), .A2(mem[415]), .B1(n2578), .B2(mem[671]), .ZN(
        n2598) );
  AOI22_X1 U2175 ( .A1(n1050), .A2(mem[863]), .B1(n2750), .B2(mem[543]), .ZN(
        n2597) );
  AOI22_X1 U2176 ( .A1(n1040), .A2(mem[223]), .B1(n1044), .B2(mem[831]), .ZN(
        n2596) );
  NAND2_X1 U2177 ( .A1(n1042), .A2(mem[255]), .ZN(n2595) );
  NAND4_X1 U2178 ( .A1(n2598), .A2(n2597), .A3(n2596), .A4(n2595), .ZN(n2614)
         );
  AOI22_X1 U2179 ( .A1(n1053), .A2(mem[447]), .B1(n1048), .B2(mem[799]), .ZN(
        n2602) );
  AOI22_X1 U2180 ( .A1(n2668), .A2(mem[639]), .B1(n1043), .B2(mem[127]), .ZN(
        n2601) );
  AOI22_X1 U2181 ( .A1(n1041), .A2(mem[191]), .B1(n3015), .B2(mem[735]), .ZN(
        n2600) );
  AOI22_X1 U2182 ( .A1(n1045), .A2(mem[31]), .B1(n1403), .B2(mem[927]), .ZN(
        n2599) );
  NAND4_X1 U2183 ( .A1(n2602), .A2(n2601), .A3(n2600), .A4(n2599), .ZN(n2613)
         );
  AOI22_X1 U2184 ( .A1(n1054), .A2(mem[351]), .B1(n1052), .B2(mem[703]), .ZN(
        n2606) );
  AOI22_X1 U2185 ( .A1(n2705), .A2(mem[767]), .B1(n1056), .B2(mem[895]), .ZN(
        n2605) );
  AOI22_X1 U2186 ( .A1(n1414), .A2(mem[63]), .B1(n1046), .B2(mem[479]), .ZN(
        n2604) );
  AOI22_X1 U2187 ( .A1(n2874), .A2(mem[383]), .B1(n1051), .B2(mem[159]), .ZN(
        n2603) );
  NAND4_X1 U2188 ( .A1(n2606), .A2(n2605), .A3(n2604), .A4(n2603), .ZN(n2612)
         );
  AOI22_X1 U2189 ( .A1(n2433), .A2(mem[607]), .B1(n1047), .B2(mem[95]), .ZN(
        n2610) );
  AOI22_X1 U2190 ( .A1(n2062), .A2(mem[511]), .B1(n1049), .B2(mem[287]), .ZN(
        n2609) );
  AOI22_X1 U2191 ( .A1(n3016), .A2(mem[319]), .B1(n1039), .B2(mem[959]), .ZN(
        n2608) );
  AOI22_X1 U2192 ( .A1(n1055), .A2(mem[991]), .B1(n3010), .B2(mem[575]), .ZN(
        n2607) );
  NAND4_X1 U2193 ( .A1(n2610), .A2(n2609), .A3(n2608), .A4(n2607), .ZN(n2611)
         );
  OR4_X1 U2194 ( .A1(n2614), .A2(n2613), .A3(n2612), .A4(n2611), .ZN(
        rdata_c_o[31]) );
  AOI22_X1 U2195 ( .A1(mem[703]), .A2(n3161), .B1(n1093), .B2(mem[511]), .ZN(
        n2618) );
  AOI22_X1 U2196 ( .A1(n1015), .A2(mem[607]), .B1(n1029), .B2(mem[127]), .ZN(
        n2617) );
  AOI22_X1 U2197 ( .A1(mem[895]), .A2(n3066), .B1(n1018), .B2(mem[223]), .ZN(
        n2616) );
  NAND2_X1 U2198 ( .A1(n1026), .A2(mem[799]), .ZN(n2615) );
  NAND4_X1 U2199 ( .A1(n2618), .A2(n2617), .A3(n2616), .A4(n2615), .ZN(n2634)
         );
  AOI22_X1 U2200 ( .A1(mem[319]), .A2(n3577), .B1(n995), .B2(mem[479]), .ZN(
        n2622) );
  AOI22_X1 U2201 ( .A1(n1024), .A2(mem[383]), .B1(mem[95]), .B2(n3579), .ZN(
        n2621) );
  AOI22_X1 U2202 ( .A1(n3585), .A2(mem[415]), .B1(mem[927]), .B2(n3594), .ZN(
        n2620) );
  AOI22_X1 U2203 ( .A1(n1081), .A2(mem[735]), .B1(mem[159]), .B2(n1021), .ZN(
        n2619) );
  NAND4_X1 U2204 ( .A1(n2622), .A2(n2621), .A3(n2620), .A4(n2619), .ZN(n2633)
         );
  AOI22_X1 U2205 ( .A1(mem[447]), .A2(n1012), .B1(n1006), .B2(mem[351]), .ZN(
        n2626) );
  AOI22_X1 U2206 ( .A1(mem[63]), .A2(n4730), .B1(n3131), .B2(mem[31]), .ZN(
        n2625) );
  AOI22_X1 U2207 ( .A1(mem[959]), .A2(n3592), .B1(n1087), .B2(mem[767]), .ZN(
        n2624) );
  AOI22_X1 U2208 ( .A1(mem[863]), .A2(n1090), .B1(n3168), .B2(mem[831]), .ZN(
        n2623) );
  NAND4_X1 U2209 ( .A1(n2626), .A2(n2625), .A3(n2624), .A4(n2623), .ZN(n2632)
         );
  AOI22_X1 U2210 ( .A1(mem[639]), .A2(n3162), .B1(n1009), .B2(mem[255]), .ZN(
        n2630) );
  AOI22_X1 U2211 ( .A1(mem[671]), .A2(n3587), .B1(n1084), .B2(mem[287]), .ZN(
        n2629) );
  AOI22_X1 U2212 ( .A1(n3383), .A2(mem[575]), .B1(mem[191]), .B2(n1072), .ZN(
        n2628) );
  AOI22_X1 U2213 ( .A1(n3167), .A2(mem[543]), .B1(mem[991]), .B2(n1073), .ZN(
        n2627) );
  NAND4_X1 U2214 ( .A1(n2630), .A2(n2629), .A3(n2628), .A4(n2627), .ZN(n2631)
         );
  OR4_X1 U2215 ( .A1(n2634), .A2(n2633), .A3(n2632), .A4(n2631), .ZN(
        rdata_a_o[31]) );
  AOI22_X1 U2216 ( .A1(n2798), .A2(mem[95]), .B1(n2954), .B2(mem[383]), .ZN(
        n2638) );
  AOI22_X1 U2217 ( .A1(n2963), .A2(mem[959]), .B1(n2974), .B2(mem[127]), .ZN(
        n2637) );
  AOI22_X1 U2218 ( .A1(n2989), .A2(mem[991]), .B1(n2786), .B2(mem[575]), .ZN(
        n2636) );
  NAND2_X1 U2219 ( .A1(n2775), .A2(mem[63]), .ZN(n2635) );
  NAND4_X1 U2220 ( .A1(n2638), .A2(n2637), .A3(n2636), .A4(n2635), .ZN(n2655)
         );
  AOI22_X1 U2221 ( .A1(n2976), .A2(mem[319]), .B1(n2835), .B2(mem[543]), .ZN(
        n2643) );
  AOI22_X1 U2222 ( .A1(n2764), .A2(mem[767]), .B1(n2955), .B2(mem[831]), .ZN(
        n2642) );
  AOI22_X1 U2223 ( .A1(n2848), .A2(mem[287]), .B1(n2953), .B2(mem[735]), .ZN(
        n2641) );
  AOI22_X1 U2224 ( .A1(n2639), .A2(mem[863]), .B1(n2957), .B2(mem[255]), .ZN(
        n2640) );
  NAND4_X1 U2225 ( .A1(n2643), .A2(n2642), .A3(n2641), .A4(n2640), .ZN(n2654)
         );
  AOI22_X1 U2226 ( .A1(n2992), .A2(mem[895]), .B1(n2833), .B2(mem[479]), .ZN(
        n2647) );
  AOI22_X1 U2227 ( .A1(n2985), .A2(mem[351]), .B1(n2965), .B2(mem[511]), .ZN(
        n2646) );
  AOI22_X1 U2228 ( .A1(n2796), .A2(mem[671]), .B1(n2951), .B2(mem[159]), .ZN(
        n2645) );
  AOI22_X1 U2229 ( .A1(n2770), .A2(mem[639]), .B1(n2975), .B2(mem[799]), .ZN(
        n2644) );
  NAND4_X1 U2230 ( .A1(n2647), .A2(n2646), .A3(n2645), .A4(n2644), .ZN(n2653)
         );
  AOI22_X1 U2231 ( .A1(n2765), .A2(mem[607]), .B1(n2979), .B2(mem[31]), .ZN(
        n2651) );
  AOI22_X1 U2232 ( .A1(n2860), .A2(mem[191]), .B1(n2987), .B2(mem[415]), .ZN(
        n2650) );
  AOI22_X1 U2233 ( .A1(n2850), .A2(mem[703]), .B1(n2832), .B2(mem[447]), .ZN(
        n2649) );
  AOI22_X1 U2234 ( .A1(n2968), .A2(mem[927]), .B1(n2977), .B2(mem[223]), .ZN(
        n2648) );
  NAND4_X1 U2235 ( .A1(n2651), .A2(n2650), .A3(n2649), .A4(n2648), .ZN(n2652)
         );
  OR4_X1 U2236 ( .A1(n2655), .A2(n2654), .A3(n2653), .A4(n2652), .ZN(
        rdata_b_o[31]) );
  AOI22_X1 U2237 ( .A1(n2433), .A2(mem[583]), .B1(n3015), .B2(mem[711]), .ZN(
        n2659) );
  AOI22_X1 U2238 ( .A1(n1033), .A2(mem[391]), .B1(n1049), .B2(mem[263]), .ZN(
        n2658) );
  AOI22_X1 U2239 ( .A1(n1050), .A2(mem[839]), .B1(n3010), .B2(mem[551]), .ZN(
        n2657) );
  NAND2_X1 U2240 ( .A1(n1052), .A2(mem[679]), .ZN(n2656) );
  NAND4_X1 U2241 ( .A1(n2659), .A2(n2658), .A3(n2657), .A4(n2656), .ZN(n2676)
         );
  AOI22_X1 U2242 ( .A1(n1045), .A2(mem[7]), .B1(n1051), .B2(mem[135]), .ZN(
        n2663) );
  AOI22_X1 U2243 ( .A1(n3016), .A2(mem[295]), .B1(n2578), .B2(mem[647]), .ZN(
        n2662) );
  AOI22_X1 U2244 ( .A1(n1054), .A2(mem[327]), .B1(n1461), .B2(mem[743]), .ZN(
        n2661) );
  AOI22_X1 U2245 ( .A1(n1040), .A2(mem[199]), .B1(n1408), .B2(mem[103]), .ZN(
        n2660) );
  NAND4_X1 U2246 ( .A1(n2663), .A2(n2662), .A3(n2661), .A4(n2660), .ZN(n2675)
         );
  AOI22_X1 U2247 ( .A1(n1055), .A2(mem[967]), .B1(n1048), .B2(mem[775]), .ZN(
        n2667) );
  AOI22_X1 U2248 ( .A1(n1047), .A2(mem[71]), .B1(n1044), .B2(mem[807]), .ZN(
        n2666) );
  AOI22_X1 U2249 ( .A1(n1039), .A2(mem[935]), .B1(n1041), .B2(mem[167]), .ZN(
        n2665) );
  AOI22_X1 U2250 ( .A1(n1740), .A2(mem[487]), .B1(n1403), .B2(mem[903]), .ZN(
        n2664) );
  NAND4_X1 U2251 ( .A1(n2667), .A2(n2666), .A3(n2665), .A4(n2664), .ZN(n2674)
         );
  AOI22_X1 U2252 ( .A1(n1414), .A2(mem[39]), .B1(n1424), .B2(mem[359]), .ZN(
        n2672) );
  AOI22_X1 U2253 ( .A1(n2668), .A2(mem[615]), .B1(n1046), .B2(mem[455]), .ZN(
        n2671) );
  AOI22_X1 U2254 ( .A1(n2750), .A2(mem[519]), .B1(n1056), .B2(mem[871]), .ZN(
        n2670) );
  AOI22_X1 U2255 ( .A1(n1042), .A2(mem[231]), .B1(n1053), .B2(mem[423]), .ZN(
        n2669) );
  NAND4_X1 U2256 ( .A1(n2672), .A2(n2671), .A3(n2670), .A4(n2669), .ZN(n2673)
         );
  OR4_X1 U2257 ( .A1(n2676), .A2(n2675), .A3(n2674), .A4(n2673), .ZN(
        rdata_c_o[7]) );
  AOI22_X1 U2258 ( .A1(n2962), .A2(mem[839]), .B1(n2967), .B2(mem[647]), .ZN(
        n2680) );
  AOI22_X1 U2259 ( .A1(n2859), .A2(mem[135]), .B1(n2841), .B2(mem[711]), .ZN(
        n2679) );
  AOI22_X1 U2260 ( .A1(n2798), .A2(mem[71]), .B1(n2955), .B2(mem[807]), .ZN(
        n2678) );
  NAND2_X1 U2261 ( .A1(n2786), .A2(mem[551]), .ZN(n2677) );
  NAND4_X1 U2262 ( .A1(n2680), .A2(n2679), .A3(n2678), .A4(n2677), .ZN(n2696)
         );
  AOI22_X1 U2263 ( .A1(n2985), .A2(mem[327]), .B1(n1228), .B2(mem[167]), .ZN(
        n2684) );
  AOI22_X1 U2264 ( .A1(n2980), .A2(mem[743]), .B1(n2954), .B2(mem[359]), .ZN(
        n2683) );
  AOI22_X1 U2265 ( .A1(n2963), .A2(mem[935]), .B1(n2851), .B2(mem[391]), .ZN(
        n2682) );
  AOI22_X1 U2266 ( .A1(n2974), .A2(mem[103]), .B1(n2976), .B2(mem[295]), .ZN(
        n2681) );
  NAND4_X1 U2267 ( .A1(n2684), .A2(n2683), .A3(n2682), .A4(n2681), .ZN(n2695)
         );
  AOI22_X1 U2268 ( .A1(n2852), .A2(mem[775]), .B1(n2965), .B2(mem[487]), .ZN(
        n2688) );
  AOI22_X1 U2269 ( .A1(n2850), .A2(mem[679]), .B1(n2776), .B2(mem[199]), .ZN(
        n2687) );
  AOI22_X1 U2270 ( .A1(n2833), .A2(mem[455]), .B1(n2989), .B2(mem[967]), .ZN(
        n2686) );
  AOI22_X1 U2271 ( .A1(n2775), .A2(mem[39]), .B1(n2835), .B2(mem[519]), .ZN(
        n2685) );
  NAND4_X1 U2272 ( .A1(n2688), .A2(n2687), .A3(n2686), .A4(n2685), .ZN(n2694)
         );
  AOI22_X1 U2273 ( .A1(n2853), .A2(mem[871]), .B1(n2785), .B2(mem[903]), .ZN(
        n2692) );
  AOI22_X1 U2274 ( .A1(n2986), .A2(mem[583]), .B1(n2957), .B2(mem[231]), .ZN(
        n2691) );
  AOI22_X1 U2275 ( .A1(n2832), .A2(mem[423]), .B1(n2979), .B2(mem[7]), .ZN(
        n2690) );
  AOI22_X1 U2276 ( .A1(n2770), .A2(mem[615]), .B1(n2848), .B2(mem[263]), .ZN(
        n2689) );
  NAND4_X1 U2277 ( .A1(n2692), .A2(n2691), .A3(n2690), .A4(n2689), .ZN(n2693)
         );
  OR4_X1 U2278 ( .A1(n2696), .A2(n2695), .A3(n2694), .A4(n2693), .ZN(
        rdata_b_o[7]) );
  AOI22_X1 U2279 ( .A1(n1053), .A2(mem[431]), .B1(n3010), .B2(mem[559]), .ZN(
        n2700) );
  AOI22_X1 U2280 ( .A1(n1041), .A2(mem[175]), .B1(n1056), .B2(mem[879]), .ZN(
        n2699) );
  AOI22_X1 U2281 ( .A1(n1045), .A2(mem[15]), .B1(n1052), .B2(mem[687]), .ZN(
        n2698) );
  NAND2_X1 U2282 ( .A1(n1408), .A2(mem[111]), .ZN(n2697) );
  NAND4_X1 U2283 ( .A1(n2700), .A2(n2699), .A3(n2698), .A4(n2697), .ZN(n2717)
         );
  AOI22_X1 U2284 ( .A1(n1033), .A2(mem[399]), .B1(n1054), .B2(mem[335]), .ZN(
        n2704) );
  AOI22_X1 U2285 ( .A1(n2062), .A2(mem[495]), .B1(n1055), .B2(mem[975]), .ZN(
        n2703) );
  AOI22_X1 U2286 ( .A1(n2869), .A2(mem[911]), .B1(n1046), .B2(mem[463]), .ZN(
        n2702) );
  AOI22_X1 U2287 ( .A1(n1039), .A2(mem[943]), .B1(n1040), .B2(mem[207]), .ZN(
        n2701) );
  NAND4_X1 U2288 ( .A1(n2704), .A2(n2703), .A3(n2702), .A4(n2701), .ZN(n2716)
         );
  AOI22_X1 U2289 ( .A1(n2705), .A2(mem[751]), .B1(n1044), .B2(mem[815]), .ZN(
        n2709) );
  AOI22_X1 U2290 ( .A1(n3015), .A2(mem[719]), .B1(n2578), .B2(mem[655]), .ZN(
        n2708) );
  AOI22_X1 U2291 ( .A1(n1042), .A2(mem[239]), .B1(n2750), .B2(mem[527]), .ZN(
        n2707) );
  AOI22_X1 U2292 ( .A1(n2433), .A2(mem[591]), .B1(n1049), .B2(mem[271]), .ZN(
        n2706) );
  NAND4_X1 U2293 ( .A1(n2709), .A2(n2708), .A3(n2707), .A4(n2706), .ZN(n2715)
         );
  AOI22_X1 U2294 ( .A1(n1414), .A2(mem[47]), .B1(n1048), .B2(mem[783]), .ZN(
        n2713) );
  AOI22_X1 U2295 ( .A1(n1050), .A2(mem[847]), .B1(n1047), .B2(mem[79]), .ZN(
        n2712) );
  AOI22_X1 U2296 ( .A1(n3016), .A2(mem[303]), .B1(n1424), .B2(mem[367]), .ZN(
        n2711) );
  AOI22_X1 U2297 ( .A1(n2668), .A2(mem[623]), .B1(n1051), .B2(mem[143]), .ZN(
        n2710) );
  NAND4_X1 U2298 ( .A1(n2713), .A2(n2712), .A3(n2711), .A4(n2710), .ZN(n2714)
         );
  OR4_X1 U2299 ( .A1(n2717), .A2(n2716), .A3(n2715), .A4(n2714), .ZN(
        rdata_c_o[15]) );
  AOI22_X1 U2300 ( .A1(n2840), .A2(mem[815]), .B1(n2786), .B2(mem[559]), .ZN(
        n2721) );
  AOI22_X1 U2301 ( .A1(n2989), .A2(mem[975]), .B1(n2985), .B2(mem[335]), .ZN(
        n2720) );
  AOI22_X1 U2302 ( .A1(n2770), .A2(mem[623]), .B1(n2835), .B2(mem[527]), .ZN(
        n2719) );
  NAND2_X1 U2303 ( .A1(n2968), .A2(mem[911]), .ZN(n2718) );
  NAND4_X1 U2304 ( .A1(n2721), .A2(n2720), .A3(n2719), .A4(n2718), .ZN(n2737)
         );
  AOI22_X1 U2305 ( .A1(n2990), .A2(mem[47]), .B1(n1228), .B2(mem[175]), .ZN(
        n2725) );
  AOI22_X1 U2306 ( .A1(n2957), .A2(mem[239]), .B1(n2966), .B2(mem[79]), .ZN(
        n2724) );
  AOI22_X1 U2307 ( .A1(n2963), .A2(mem[943]), .B1(n2841), .B2(mem[719]), .ZN(
        n2723) );
  AOI22_X1 U2308 ( .A1(n2843), .A2(mem[111]), .B1(n2954), .B2(mem[367]), .ZN(
        n2722) );
  NAND4_X1 U2309 ( .A1(n2725), .A2(n2724), .A3(n2723), .A4(n2722), .ZN(n2736)
         );
  AOI22_X1 U2310 ( .A1(n2852), .A2(mem[783]), .B1(n2848), .B2(mem[271]), .ZN(
        n2729) );
  AOI22_X1 U2311 ( .A1(n2833), .A2(mem[463]), .B1(n2776), .B2(mem[207]), .ZN(
        n2728) );
  AOI22_X1 U2312 ( .A1(n2962), .A2(mem[847]), .B1(n2951), .B2(mem[143]), .ZN(
        n2727) );
  AOI22_X1 U2313 ( .A1(n2965), .A2(mem[495]), .B1(n2976), .B2(mem[303]), .ZN(
        n2726) );
  NAND4_X1 U2314 ( .A1(n2729), .A2(n2728), .A3(n2727), .A4(n2726), .ZN(n2735)
         );
  AOI22_X1 U2315 ( .A1(n2850), .A2(mem[687]), .B1(n2765), .B2(mem[591]), .ZN(
        n2733) );
  AOI22_X1 U2316 ( .A1(n2979), .A2(mem[15]), .B1(n2851), .B2(mem[399]), .ZN(
        n2732) );
  AOI22_X1 U2317 ( .A1(n2764), .A2(mem[751]), .B1(n2992), .B2(mem[879]), .ZN(
        n2731) );
  AOI22_X1 U2318 ( .A1(n2796), .A2(mem[655]), .B1(n2964), .B2(mem[431]), .ZN(
        n2730) );
  NAND4_X1 U2319 ( .A1(n2733), .A2(n2732), .A3(n2731), .A4(n2730), .ZN(n2734)
         );
  OR4_X1 U2320 ( .A1(n2737), .A2(n2736), .A3(n2735), .A4(n2734), .ZN(
        rdata_b_o[15]) );
  AOI22_X1 U2321 ( .A1(n1041), .A2(mem[174]), .B1(n2869), .B2(mem[910]), .ZN(
        n2741) );
  AOI22_X1 U2322 ( .A1(n1056), .A2(mem[878]), .B1(n1049), .B2(mem[270]), .ZN(
        n2740) );
  AOI22_X1 U2323 ( .A1(n3016), .A2(mem[302]), .B1(n1424), .B2(mem[366]), .ZN(
        n2739) );
  NAND2_X1 U2324 ( .A1(n1051), .A2(mem[142]), .ZN(n2738) );
  NAND4_X1 U2325 ( .A1(n2741), .A2(n2740), .A3(n2739), .A4(n2738), .ZN(n2758)
         );
  AOI22_X1 U2326 ( .A1(n1042), .A2(mem[238]), .B1(n2705), .B2(mem[750]), .ZN(
        n2745) );
  AOI22_X1 U2327 ( .A1(n3010), .A2(mem[558]), .B1(n1043), .B2(mem[110]), .ZN(
        n2744) );
  AOI22_X1 U2328 ( .A1(n3015), .A2(mem[718]), .B1(n1046), .B2(mem[462]), .ZN(
        n2743) );
  AOI22_X1 U2329 ( .A1(n3001), .A2(mem[46]), .B1(n1402), .B2(mem[942]), .ZN(
        n2742) );
  NAND4_X1 U2330 ( .A1(n2745), .A2(n2744), .A3(n2743), .A4(n2742), .ZN(n2757)
         );
  AOI22_X1 U2331 ( .A1(n1054), .A2(mem[334]), .B1(n1047), .B2(mem[78]), .ZN(
        n2749) );
  AOI22_X1 U2332 ( .A1(n2433), .A2(mem[590]), .B1(n2578), .B2(mem[654]), .ZN(
        n2748) );
  AOI22_X1 U2333 ( .A1(n1045), .A2(mem[14]), .B1(n1053), .B2(mem[430]), .ZN(
        n2747) );
  AOI22_X1 U2334 ( .A1(n1050), .A2(mem[846]), .B1(n1044), .B2(mem[814]), .ZN(
        n2746) );
  NAND4_X1 U2335 ( .A1(n2749), .A2(n2748), .A3(n2747), .A4(n2746), .ZN(n2756)
         );
  AOI22_X1 U2336 ( .A1(n2062), .A2(mem[494]), .B1(n2750), .B2(mem[526]), .ZN(
        n2754) );
  AOI22_X1 U2337 ( .A1(n1055), .A2(mem[974]), .B1(n1052), .B2(mem[686]), .ZN(
        n2753) );
  AOI22_X1 U2338 ( .A1(n1040), .A2(mem[206]), .B1(n1048), .B2(mem[782]), .ZN(
        n2752) );
  AOI22_X1 U2339 ( .A1(n1745), .A2(mem[622]), .B1(n1033), .B2(mem[398]), .ZN(
        n2751) );
  NAND4_X1 U2340 ( .A1(n2754), .A2(n2753), .A3(n2752), .A4(n2751), .ZN(n2755)
         );
  OR4_X1 U2341 ( .A1(n2758), .A2(n2757), .A3(n2756), .A4(n2755), .ZN(
        rdata_c_o[14]) );
  AOI22_X1 U2342 ( .A1(n2963), .A2(mem[942]), .B1(n2966), .B2(mem[78]), .ZN(
        n2763) );
  AOI22_X1 U2343 ( .A1(n2759), .A2(mem[334]), .B1(n2859), .B2(mem[142]), .ZN(
        n2762) );
  AOI22_X1 U2344 ( .A1(n2796), .A2(mem[654]), .B1(n2851), .B2(mem[398]), .ZN(
        n2761) );
  NAND2_X1 U2345 ( .A1(n2850), .A2(mem[686]), .ZN(n2760) );
  NAND4_X1 U2346 ( .A1(n2763), .A2(n2762), .A3(n2761), .A4(n2760), .ZN(n2784)
         );
  AOI22_X1 U2347 ( .A1(n2764), .A2(mem[750]), .B1(n2955), .B2(mem[814]), .ZN(
        n2769) );
  AOI22_X1 U2348 ( .A1(n2853), .A2(mem[878]), .B1(n2965), .B2(mem[494]), .ZN(
        n2768) );
  AOI22_X1 U2349 ( .A1(n2860), .A2(mem[174]), .B1(n2786), .B2(mem[558]), .ZN(
        n2767) );
  AOI22_X1 U2350 ( .A1(n2833), .A2(mem[462]), .B1(n2765), .B2(mem[590]), .ZN(
        n2766) );
  NAND4_X1 U2351 ( .A1(n2769), .A2(n2768), .A3(n2767), .A4(n2766), .ZN(n2783)
         );
  AOI22_X1 U2352 ( .A1(n2832), .A2(mem[430]), .B1(n2954), .B2(mem[366]), .ZN(
        n2774) );
  AOI22_X1 U2353 ( .A1(n2770), .A2(mem[622]), .B1(n2974), .B2(mem[110]), .ZN(
        n2773) );
  AOI22_X1 U2354 ( .A1(n2848), .A2(mem[270]), .B1(n2835), .B2(mem[526]), .ZN(
        n2772) );
  AOI22_X1 U2355 ( .A1(n2976), .A2(mem[302]), .B1(n2979), .B2(mem[14]), .ZN(
        n2771) );
  NAND4_X1 U2356 ( .A1(n2774), .A2(n2773), .A3(n2772), .A4(n2771), .ZN(n2782)
         );
  AOI22_X1 U2357 ( .A1(n2785), .A2(mem[910]), .B1(n2957), .B2(mem[238]), .ZN(
        n2780) );
  AOI22_X1 U2358 ( .A1(n2775), .A2(mem[46]), .B1(n2953), .B2(mem[718]), .ZN(
        n2779) );
  AOI22_X1 U2359 ( .A1(n2962), .A2(mem[846]), .B1(n2989), .B2(mem[974]), .ZN(
        n2778) );
  AOI22_X1 U2360 ( .A1(n2852), .A2(mem[782]), .B1(n2776), .B2(mem[206]), .ZN(
        n2777) );
  NAND4_X1 U2361 ( .A1(n2780), .A2(n2779), .A3(n2778), .A4(n2777), .ZN(n2781)
         );
  OR4_X1 U2362 ( .A1(n2784), .A2(n2783), .A3(n2782), .A4(n2781), .ZN(
        rdata_b_o[14]) );
  AOI22_X1 U2363 ( .A1(n2785), .A2(mem[914]), .B1(n2974), .B2(mem[114]), .ZN(
        n2790) );
  AOI22_X1 U2364 ( .A1(n2952), .A2(mem[466]), .B1(n2851), .B2(mem[402]), .ZN(
        n2789) );
  AOI22_X1 U2365 ( .A1(n2955), .A2(mem[818]), .B1(n2786), .B2(mem[562]), .ZN(
        n2788) );
  NAND2_X1 U2366 ( .A1(n2853), .A2(mem[882]), .ZN(n2787) );
  NAND4_X1 U2367 ( .A1(n2790), .A2(n2789), .A3(n2788), .A4(n2787), .ZN(n2811)
         );
  AOI22_X1 U2368 ( .A1(n2990), .A2(mem[50]), .B1(n2962), .B2(mem[850]), .ZN(
        n2795) );
  AOI22_X1 U2369 ( .A1(n2791), .A2(mem[978]), .B1(n2965), .B2(mem[498]), .ZN(
        n2794) );
  AOI22_X1 U2370 ( .A1(n2951), .A2(mem[146]), .B1(n2976), .B2(mem[306]), .ZN(
        n2793) );
  AOI22_X1 U2371 ( .A1(n2977), .A2(mem[210]), .B1(n1228), .B2(mem[178]), .ZN(
        n2792) );
  NAND4_X1 U2372 ( .A1(n2795), .A2(n2794), .A3(n2793), .A4(n2792), .ZN(n2810)
         );
  AOI22_X1 U2373 ( .A1(n2796), .A2(mem[658]), .B1(n2985), .B2(mem[338]), .ZN(
        n2802) );
  AOI22_X1 U2374 ( .A1(n2797), .A2(mem[946]), .B1(n2956), .B2(mem[626]), .ZN(
        n2801) );
  AOI22_X1 U2375 ( .A1(n2986), .A2(mem[594]), .B1(n2798), .B2(mem[82]), .ZN(
        n2800) );
  AOI22_X1 U2376 ( .A1(n2969), .A2(mem[690]), .B1(n2975), .B2(mem[786]), .ZN(
        n2799) );
  NAND4_X1 U2377 ( .A1(n2802), .A2(n2801), .A3(n2800), .A4(n2799), .ZN(n2809)
         );
  AOI22_X1 U2378 ( .A1(n2842), .A2(mem[370]), .B1(n2953), .B2(mem[722]), .ZN(
        n2807) );
  AOI22_X1 U2379 ( .A1(n2980), .A2(mem[754]), .B1(n2988), .B2(mem[530]), .ZN(
        n2806) );
  AOI22_X1 U2380 ( .A1(n2803), .A2(mem[242]), .B1(n2848), .B2(mem[274]), .ZN(
        n2805) );
  AOI22_X1 U2381 ( .A1(n2832), .A2(mem[434]), .B1(n2834), .B2(mem[18]), .ZN(
        n2804) );
  NAND4_X1 U2382 ( .A1(n2807), .A2(n2806), .A3(n2805), .A4(n2804), .ZN(n2808)
         );
  OR4_X1 U2383 ( .A1(n2811), .A2(n2810), .A3(n2809), .A4(n2808), .ZN(
        rdata_b_o[18]) );
  AOI22_X1 U2384 ( .A1(n1752), .A2(mem[594]), .B1(n3001), .B2(mem[50]), .ZN(
        n2815) );
  AOI22_X1 U2385 ( .A1(n3015), .A2(mem[722]), .B1(n1049), .B2(mem[274]), .ZN(
        n2814) );
  AOI22_X1 U2386 ( .A1(n1044), .A2(mem[818]), .B1(n1056), .B2(mem[882]), .ZN(
        n2813) );
  NAND2_X1 U2387 ( .A1(n2705), .A2(mem[754]), .ZN(n2812) );
  NAND4_X1 U2388 ( .A1(n2815), .A2(n2814), .A3(n2813), .A4(n2812), .ZN(n2831)
         );
  AOI22_X1 U2389 ( .A1(n1039), .A2(mem[946]), .B1(n2869), .B2(mem[914]), .ZN(
        n2819) );
  AOI22_X1 U2390 ( .A1(n1040), .A2(mem[210]), .B1(n1051), .B2(mem[146]), .ZN(
        n2818) );
  AOI22_X1 U2391 ( .A1(n1046), .A2(mem[466]), .B1(n1043), .B2(mem[114]), .ZN(
        n2817) );
  AOI22_X1 U2392 ( .A1(n1055), .A2(mem[978]), .B1(n2067), .B2(mem[658]), .ZN(
        n2816) );
  NAND4_X1 U2393 ( .A1(n2819), .A2(n2818), .A3(n2817), .A4(n2816), .ZN(n2830)
         );
  AOI22_X1 U2394 ( .A1(n1054), .A2(mem[338]), .B1(n1052), .B2(mem[690]), .ZN(
        n2823) );
  AOI22_X1 U2395 ( .A1(n1042), .A2(mem[242]), .B1(n1053), .B2(mem[434]), .ZN(
        n2822) );
  AOI22_X1 U2396 ( .A1(n2668), .A2(mem[626]), .B1(n1394), .B2(mem[562]), .ZN(
        n2821) );
  AOI22_X1 U2397 ( .A1(n1740), .A2(mem[498]), .B1(n1474), .B2(mem[530]), .ZN(
        n2820) );
  NAND4_X1 U2398 ( .A1(n2823), .A2(n2822), .A3(n2821), .A4(n2820), .ZN(n2829)
         );
  AOI22_X1 U2399 ( .A1(n1751), .A2(mem[18]), .B1(n2874), .B2(mem[370]), .ZN(
        n2827) );
  AOI22_X1 U2400 ( .A1(n1033), .A2(mem[402]), .B1(n1430), .B2(mem[178]), .ZN(
        n2826) );
  AOI22_X1 U2401 ( .A1(n3016), .A2(mem[306]), .B1(n1047), .B2(mem[82]), .ZN(
        n2825) );
  AOI22_X1 U2402 ( .A1(n1050), .A2(mem[850]), .B1(n1048), .B2(mem[786]), .ZN(
        n2824) );
  NAND4_X1 U2403 ( .A1(n2827), .A2(n2826), .A3(n2825), .A4(n2824), .ZN(n2828)
         );
  OR4_X1 U2404 ( .A1(n2831), .A2(n2830), .A3(n2829), .A4(n2828), .ZN(
        rdata_c_o[18]) );
  AOI22_X1 U2405 ( .A1(n2968), .A2(mem[917]), .B1(n2832), .B2(mem[437]), .ZN(
        n2839) );
  AOI22_X1 U2406 ( .A1(n2833), .A2(mem[469]), .B1(n2986), .B2(mem[597]), .ZN(
        n2838) );
  AOI22_X1 U2407 ( .A1(n2835), .A2(mem[533]), .B1(n2834), .B2(mem[21]), .ZN(
        n2837) );
  NAND2_X1 U2408 ( .A1(n2989), .A2(mem[981]), .ZN(n2836) );
  NAND4_X1 U2409 ( .A1(n2839), .A2(n2838), .A3(n2837), .A4(n2836), .ZN(n2868)
         );
  AOI22_X1 U2410 ( .A1(n2990), .A2(mem[53]), .B1(n2985), .B2(mem[341]), .ZN(
        n2847) );
  AOI22_X1 U2411 ( .A1(n2980), .A2(mem[757]), .B1(n2840), .B2(mem[821]), .ZN(
        n2846) );
  AOI22_X1 U2412 ( .A1(n2842), .A2(mem[373]), .B1(n2841), .B2(mem[725]), .ZN(
        n2845) );
  AOI22_X1 U2413 ( .A1(n2956), .A2(mem[629]), .B1(n2843), .B2(mem[117]), .ZN(
        n2844) );
  NAND4_X1 U2414 ( .A1(n2847), .A2(n2846), .A3(n2845), .A4(n2844), .ZN(n2867)
         );
  AOI22_X1 U2415 ( .A1(n2977), .A2(mem[213]), .B1(n2848), .B2(mem[277]), .ZN(
        n2857) );
  AOI22_X1 U2416 ( .A1(n2850), .A2(mem[693]), .B1(n2849), .B2(mem[501]), .ZN(
        n2856) );
  AOI22_X1 U2417 ( .A1(n2852), .A2(mem[789]), .B1(n2851), .B2(mem[405]), .ZN(
        n2855) );
  AOI22_X1 U2418 ( .A1(n2853), .A2(mem[885]), .B1(n2957), .B2(mem[245]), .ZN(
        n2854) );
  NAND4_X1 U2419 ( .A1(n2857), .A2(n2856), .A3(n2855), .A4(n2854), .ZN(n2866)
         );
  AOI22_X1 U2420 ( .A1(n2859), .A2(mem[149]), .B1(n2858), .B2(mem[309]), .ZN(
        n2864) );
  AOI22_X1 U2421 ( .A1(n2963), .A2(mem[949]), .B1(n2966), .B2(mem[85]), .ZN(
        n2863) );
  AOI22_X1 U2422 ( .A1(n2962), .A2(mem[853]), .B1(n2967), .B2(mem[661]), .ZN(
        n2862) );
  AOI22_X1 U2423 ( .A1(n2860), .A2(mem[181]), .B1(n2991), .B2(mem[565]), .ZN(
        n2861) );
  NAND4_X1 U2424 ( .A1(n2864), .A2(n2863), .A3(n2862), .A4(n2861), .ZN(n2865)
         );
  OR4_X1 U2425 ( .A1(n2868), .A2(n2867), .A3(n2866), .A4(n2865), .ZN(
        rdata_b_o[21]) );
  AOI22_X1 U2426 ( .A1(n1752), .A2(mem[597]), .B1(n2869), .B2(mem[917]), .ZN(
        n2873) );
  AOI22_X1 U2427 ( .A1(n1040), .A2(mem[213]), .B1(n1049), .B2(mem[277]), .ZN(
        n2872) );
  AOI22_X1 U2428 ( .A1(n1740), .A2(mem[501]), .B1(n3016), .B2(mem[309]), .ZN(
        n2871) );
  NAND2_X1 U2429 ( .A1(n1052), .A2(mem[693]), .ZN(n2870) );
  NAND4_X1 U2430 ( .A1(n2873), .A2(n2872), .A3(n2871), .A4(n2870), .ZN(n2890)
         );
  AOI22_X1 U2431 ( .A1(n1042), .A2(mem[245]), .B1(n2705), .B2(mem[757]), .ZN(
        n2878) );
  AOI22_X1 U2432 ( .A1(n1033), .A2(mem[405]), .B1(n1041), .B2(mem[181]), .ZN(
        n2877) );
  AOI22_X1 U2433 ( .A1(n1055), .A2(mem[981]), .B1(n1043), .B2(mem[117]), .ZN(
        n2876) );
  AOI22_X1 U2434 ( .A1(n2874), .A2(mem[373]), .B1(n2750), .B2(mem[533]), .ZN(
        n2875) );
  NAND4_X1 U2435 ( .A1(n2878), .A2(n2877), .A3(n2876), .A4(n2875), .ZN(n2889)
         );
  AOI22_X1 U2436 ( .A1(n1046), .A2(mem[469]), .B1(n1044), .B2(mem[821]), .ZN(
        n2882) );
  AOI22_X1 U2437 ( .A1(n1050), .A2(mem[853]), .B1(n2578), .B2(mem[661]), .ZN(
        n2881) );
  AOI22_X1 U2438 ( .A1(n1053), .A2(mem[437]), .B1(n1056), .B2(mem[885]), .ZN(
        n2880) );
  AOI22_X1 U2439 ( .A1(n1745), .A2(mem[629]), .B1(n3001), .B2(mem[53]), .ZN(
        n2879) );
  NAND4_X1 U2440 ( .A1(n2882), .A2(n2881), .A3(n2880), .A4(n2879), .ZN(n2888)
         );
  AOI22_X1 U2441 ( .A1(n3015), .A2(mem[725]), .B1(n1051), .B2(mem[149]), .ZN(
        n2886) );
  AOI22_X1 U2442 ( .A1(n1039), .A2(mem[949]), .B1(n3010), .B2(mem[565]), .ZN(
        n2885) );
  AOI22_X1 U2443 ( .A1(n1045), .A2(mem[21]), .B1(n1048), .B2(mem[789]), .ZN(
        n2884) );
  AOI22_X1 U2444 ( .A1(n1054), .A2(mem[341]), .B1(n1047), .B2(mem[85]), .ZN(
        n2883) );
  NAND4_X1 U2445 ( .A1(n2886), .A2(n2885), .A3(n2884), .A4(n2883), .ZN(n2887)
         );
  OR4_X1 U2446 ( .A1(n2890), .A2(n2889), .A3(n2888), .A4(n2887), .ZN(
        rdata_c_o[21]) );
  AOI22_X1 U2447 ( .A1(mem[579]), .A2(n1014), .B1(n994), .B2(mem[451]), .ZN(
        n2894) );
  AOI22_X1 U2448 ( .A1(mem[323]), .A2(n1006), .B1(n1083), .B2(mem[259]), .ZN(
        n2893) );
  AOI22_X1 U2449 ( .A1(mem[707]), .A2(n1080), .B1(n1012), .B2(mem[419]), .ZN(
        n2892) );
  AOI22_X1 U2450 ( .A1(n1010), .A2(mem[227]), .B1(mem[131]), .B2(n1020), .ZN(
        n2891) );
  AOI22_X1 U2451 ( .A1(mem[675]), .A2(n3161), .B1(n3112), .B2(mem[387]), .ZN(
        n2898) );
  AOI22_X1 U2452 ( .A1(mem[611]), .A2(n3162), .B1(n3113), .B2(mem[547]), .ZN(
        n2897) );
  AOI22_X1 U2453 ( .A1(mem[99]), .A2(n1031), .B1(n1019), .B2(mem[195]), .ZN(
        n2896) );
  AOI22_X1 U2454 ( .A1(n3587), .A2(mem[643]), .B1(mem[163]), .B2(n1072), .ZN(
        n2895) );
  AOI22_X1 U2455 ( .A1(mem[355]), .A2(n1024), .B1(n2162), .B2(mem[291]), .ZN(
        n2902) );
  AOI22_X1 U2456 ( .A1(mem[67]), .A2(n3579), .B1(n3131), .B2(mem[3]), .ZN(
        n2901) );
  AOI22_X1 U2457 ( .A1(n1067), .A2(mem[483]), .B1(mem[35]), .B2(n4730), .ZN(
        n2900) );
  NAND2_X1 U2458 ( .A1(n1026), .A2(mem[771]), .ZN(n2899) );
  AOI22_X1 U2459 ( .A1(n3167), .A2(mem[515]), .B1(mem[931]), .B2(n3221), .ZN(
        n2906) );
  AOI22_X1 U2460 ( .A1(mem[963]), .A2(n1073), .B1(n1088), .B2(mem[739]), .ZN(
        n2905) );
  AOI22_X1 U2461 ( .A1(mem[867]), .A2(n3066), .B1(n3168), .B2(mem[803]), .ZN(
        n2904) );
  AOI22_X1 U2462 ( .A1(mem[899]), .A2(n3269), .B1(n1091), .B2(mem[835]), .ZN(
        n2903) );
  NAND4_X1 U2463 ( .A1(n2906), .A2(n2905), .A3(n2904), .A4(n2903), .ZN(n2907)
         );
  AOI22_X1 U2464 ( .A1(mem[577]), .A2(n1015), .B1(n995), .B2(mem[449]), .ZN(
        n2911) );
  AOI22_X1 U2465 ( .A1(mem[321]), .A2(n1006), .B1(n1085), .B2(mem[257]), .ZN(
        n2910) );
  AOI22_X1 U2466 ( .A1(mem[705]), .A2(n1081), .B1(n1013), .B2(mem[417]), .ZN(
        n2909) );
  AOI22_X1 U2467 ( .A1(n1009), .A2(mem[225]), .B1(mem[129]), .B2(n1020), .ZN(
        n2908) );
  AOI22_X1 U2469 ( .A1(mem[673]), .A2(n3161), .B1(n3112), .B2(mem[385]), .ZN(
        n2915) );
  AOI22_X1 U2470 ( .A1(mem[609]), .A2(n3162), .B1(n3113), .B2(mem[545]), .ZN(
        n2914) );
  AOI22_X1 U2471 ( .A1(mem[97]), .A2(n1029), .B1(n1018), .B2(mem[193]), .ZN(
        n2913) );
  AOI22_X1 U2472 ( .A1(n3587), .A2(mem[641]), .B1(mem[161]), .B2(n3517), .ZN(
        n2912) );
  AOI22_X1 U2474 ( .A1(mem[353]), .A2(n1024), .B1(n2162), .B2(mem[289]), .ZN(
        n2919) );
  AOI22_X1 U2475 ( .A1(mem[65]), .A2(n3579), .B1(n3131), .B2(mem[1]), .ZN(
        n2918) );
  AOI22_X1 U2476 ( .A1(n1093), .A2(mem[481]), .B1(mem[33]), .B2(n4729), .ZN(
        n2917) );
  NAND2_X1 U2477 ( .A1(n1027), .A2(mem[769]), .ZN(n2916) );
  AOI22_X1 U2479 ( .A1(n3167), .A2(mem[513]), .B1(mem[929]), .B2(n3592), .ZN(
        n2923) );
  AOI22_X1 U2480 ( .A1(mem[961]), .A2(n1073), .B1(n1087), .B2(mem[737]), .ZN(
        n2922) );
  AOI22_X1 U2481 ( .A1(mem[865]), .A2(n3066), .B1(n3168), .B2(mem[801]), .ZN(
        n2921) );
  AOI22_X1 U2482 ( .A1(mem[897]), .A2(n3269), .B1(n1090), .B2(mem[833]), .ZN(
        n2920) );
  AOI22_X1 U2528 ( .A1(n2952), .A2(mem[473]), .B1(n2951), .B2(mem[153]), .ZN(
        n2961) );
  AOI22_X1 U2529 ( .A1(n2954), .A2(mem[377]), .B1(n2953), .B2(mem[729]), .ZN(
        n2960) );
  AOI22_X1 U2530 ( .A1(n2956), .A2(mem[633]), .B1(n2955), .B2(mem[825]), .ZN(
        n2959) );
  NAND2_X1 U2531 ( .A1(n2957), .A2(mem[249]), .ZN(n2958) );
  NAND4_X1 U2532 ( .A1(n2961), .A2(n2960), .A3(n2959), .A4(n2958), .ZN(n3000)
         );
  AOI22_X1 U2533 ( .A1(n2963), .A2(mem[953]), .B1(n2962), .B2(mem[857]), .ZN(
        n2973) );
  AOI22_X1 U2534 ( .A1(n2965), .A2(mem[505]), .B1(n2964), .B2(mem[441]), .ZN(
        n2972) );
  AOI22_X1 U2535 ( .A1(n2967), .A2(mem[665]), .B1(n2966), .B2(mem[89]), .ZN(
        n2971) );
  AOI22_X1 U2536 ( .A1(n2969), .A2(mem[697]), .B1(n2968), .B2(mem[921]), .ZN(
        n2970) );
  NAND4_X1 U2537 ( .A1(n2973), .A2(n2972), .A3(n2971), .A4(n2970), .ZN(n2999)
         );
  AOI22_X1 U2538 ( .A1(n2975), .A2(mem[793]), .B1(n2974), .B2(mem[121]), .ZN(
        n2984) );
  AOI22_X1 U2539 ( .A1(n2977), .A2(mem[217]), .B1(n2976), .B2(mem[313]), .ZN(
        n2983) );
  AOI22_X1 U2540 ( .A1(n2978), .A2(mem[281]), .B1(n2860), .B2(mem[185]), .ZN(
        n2982) );
  AOI22_X1 U2541 ( .A1(n2980), .A2(mem[761]), .B1(n2979), .B2(mem[25]), .ZN(
        n2981) );
  NAND4_X1 U2542 ( .A1(n2984), .A2(n2983), .A3(n2982), .A4(n2981), .ZN(n2998)
         );
  AOI22_X1 U2543 ( .A1(n2986), .A2(mem[601]), .B1(n2985), .B2(mem[345]), .ZN(
        n2996) );
  AOI22_X1 U2544 ( .A1(n2988), .A2(mem[537]), .B1(n2987), .B2(mem[409]), .ZN(
        n2995) );
  AOI22_X1 U2545 ( .A1(n2990), .A2(mem[57]), .B1(n2989), .B2(mem[985]), .ZN(
        n2994) );
  AOI22_X1 U2546 ( .A1(n2992), .A2(mem[889]), .B1(n2991), .B2(mem[569]), .ZN(
        n2993) );
  NAND4_X1 U2547 ( .A1(n2996), .A2(n2995), .A3(n2994), .A4(n2993), .ZN(n2997)
         );
  OR4_X1 U2548 ( .A1(n3000), .A2(n2999), .A3(n2998), .A4(n2997), .ZN(
        rdata_b_o[25]) );
  AOI22_X1 U2549 ( .A1(n3001), .A2(mem[57]), .B1(n1054), .B2(mem[345]), .ZN(
        n3005) );
  AOI22_X1 U2550 ( .A1(n1040), .A2(mem[217]), .B1(n2578), .B2(mem[665]), .ZN(
        n3004) );
  AOI22_X1 U2551 ( .A1(n1740), .A2(mem[505]), .B1(n1046), .B2(mem[473]), .ZN(
        n3003) );
  NAND2_X1 U2552 ( .A1(n1052), .A2(mem[697]), .ZN(n3002) );
  NAND4_X1 U2553 ( .A1(n3005), .A2(n3004), .A3(n3003), .A4(n3002), .ZN(n3024)
         );
  AOI22_X1 U2554 ( .A1(n1033), .A2(mem[409]), .B1(n1051), .B2(mem[153]), .ZN(
        n3009) );
  AOI22_X1 U2555 ( .A1(n1041), .A2(mem[185]), .B1(n1056), .B2(mem[889]), .ZN(
        n3008) );
  AOI22_X1 U2556 ( .A1(n2668), .A2(mem[633]), .B1(n2874), .B2(mem[377]), .ZN(
        n3007) );
  AOI22_X1 U2557 ( .A1(n1050), .A2(mem[857]), .B1(n1055), .B2(mem[985]), .ZN(
        n3006) );
  NAND4_X1 U2558 ( .A1(n3009), .A2(n3008), .A3(n3007), .A4(n3006), .ZN(n3023)
         );
  AOI22_X1 U2559 ( .A1(n2433), .A2(mem[601]), .B1(n1053), .B2(mem[441]), .ZN(
        n3014) );
  AOI22_X1 U2560 ( .A1(n2869), .A2(mem[921]), .B1(n1461), .B2(mem[761]), .ZN(
        n3013) );
  AOI22_X1 U2561 ( .A1(n1048), .A2(mem[793]), .B1(n3010), .B2(mem[569]), .ZN(
        n3012) );
  AOI22_X1 U2562 ( .A1(n2750), .A2(mem[537]), .B1(n1049), .B2(mem[281]), .ZN(
        n3011) );
  NAND4_X1 U2563 ( .A1(n3014), .A2(n3013), .A3(n3012), .A4(n3011), .ZN(n3022)
         );
  AOI22_X1 U2564 ( .A1(n1045), .A2(mem[25]), .B1(n3015), .B2(mem[729]), .ZN(
        n3020) );
  AOI22_X1 U2565 ( .A1(n3016), .A2(mem[313]), .B1(n1043), .B2(mem[121]), .ZN(
        n3019) );
  AOI22_X1 U2566 ( .A1(n1039), .A2(mem[953]), .B1(n1047), .B2(mem[89]), .ZN(
        n3018) );
  AOI22_X1 U2567 ( .A1(n1042), .A2(mem[249]), .B1(n1044), .B2(mem[825]), .ZN(
        n3017) );
  NAND4_X1 U2568 ( .A1(n3020), .A2(n3019), .A3(n3018), .A4(n3017), .ZN(n3021)
         );
  OR4_X1 U2569 ( .A1(n3024), .A2(n3023), .A3(n3022), .A4(n3021), .ZN(
        rdata_c_o[25]) );
  AOI22_X1 U2570 ( .A1(mem[320]), .A2(n1007), .B1(n1083), .B2(mem[256]), .ZN(
        n3026) );
  AOI22_X1 U2571 ( .A1(mem[704]), .A2(n1080), .B1(n1013), .B2(mem[416]), .ZN(
        n3025) );
  NAND2_X1 U2572 ( .A1(n3026), .A2(n3025), .ZN(n3035) );
  AOI22_X1 U2573 ( .A1(mem[576]), .A2(n1016), .B1(n994), .B2(mem[448]), .ZN(
        n3028) );
  AOI22_X1 U2574 ( .A1(n1010), .A2(mem[224]), .B1(mem[128]), .B2(n1022), .ZN(
        n3027) );
  NAND2_X1 U2575 ( .A1(n3028), .A2(n3027), .ZN(n3034) );
  AOI22_X1 U2576 ( .A1(mem[352]), .A2(n1024), .B1(n2162), .B2(mem[288]), .ZN(
        n3032) );
  AOI22_X1 U2577 ( .A1(n1093), .A2(mem[480]), .B1(mem[32]), .B2(n4730), .ZN(
        n3031) );
  AOI22_X1 U2578 ( .A1(mem[64]), .A2(n3579), .B1(n3131), .B2(mem[0]), .ZN(
        n3030) );
  NAND2_X1 U2579 ( .A1(n1025), .A2(mem[768]), .ZN(n3029) );
  NAND4_X1 U2580 ( .A1(n3032), .A2(n3031), .A3(n3030), .A4(n3029), .ZN(n3033)
         );
  NOR3_X1 U2581 ( .A1(n3035), .A2(n3034), .A3(n3033), .ZN(n3048) );
  AOI22_X1 U2582 ( .A1(mem[672]), .A2(n3161), .B1(n3112), .B2(mem[384]), .ZN(
        n3039) );
  AOI22_X1 U2583 ( .A1(n1019), .A2(mem[192]), .B1(mem[96]), .B2(n1029), .ZN(
        n3038) );
  AOI22_X1 U2584 ( .A1(mem[608]), .A2(n3162), .B1(n3113), .B2(mem[544]), .ZN(
        n3037) );
  AOI22_X1 U2585 ( .A1(n3061), .A2(mem[640]), .B1(mem[160]), .B2(n1072), .ZN(
        n3036) );
  NAND4_X1 U2586 ( .A1(n3039), .A2(n3038), .A3(n3037), .A4(n3036), .ZN(n3046)
         );
  BUF_X1 U2587 ( .A(n3040), .Z(n3433) );
  AOI22_X1 U2588 ( .A1(n3167), .A2(mem[512]), .B1(mem[928]), .B2(n3433), .ZN(
        n3044) );
  AOI22_X1 U2589 ( .A1(mem[960]), .A2(n1073), .B1(n1088), .B2(mem[736]), .ZN(
        n3043) );
  AOI22_X1 U2590 ( .A1(mem[864]), .A2(n3066), .B1(n3168), .B2(mem[800]), .ZN(
        n3042) );
  AOI22_X1 U2591 ( .A1(mem[896]), .A2(n3455), .B1(n1090), .B2(mem[832]), .ZN(
        n3041) );
  NAND4_X1 U2592 ( .A1(n3044), .A2(n3043), .A3(n3042), .A4(n3041), .ZN(n3045)
         );
  NOR2_X1 U2593 ( .A1(n3046), .A2(n3045), .ZN(n3047) );
  NAND2_X1 U2594 ( .A1(n3048), .A2(n3047), .ZN(rdata_a_o[0]) );
  AOI22_X1 U2595 ( .A1(mem[322]), .A2(n1005), .B1(n1083), .B2(mem[258]), .ZN(
        n3050) );
  AOI22_X1 U2596 ( .A1(mem[706]), .A2(n1082), .B1(n1011), .B2(mem[418]), .ZN(
        n3049) );
  NAND2_X1 U2597 ( .A1(n3050), .A2(n3049), .ZN(n3060) );
  AOI22_X1 U2598 ( .A1(mem[578]), .A2(n1015), .B1(n995), .B2(mem[450]), .ZN(
        n3052) );
  AOI22_X1 U2599 ( .A1(n1008), .A2(mem[226]), .B1(mem[130]), .B2(n1021), .ZN(
        n3051) );
  NAND2_X1 U2600 ( .A1(n3052), .A2(n3051), .ZN(n3059) );
  AOI22_X1 U2601 ( .A1(mem[354]), .A2(n1023), .B1(n2162), .B2(mem[290]), .ZN(
        n3057) );
  AOI22_X1 U2602 ( .A1(n1092), .A2(mem[482]), .B1(mem[34]), .B2(n4729), .ZN(
        n3056) );
  AOI22_X1 U2603 ( .A1(mem[66]), .A2(n3579), .B1(n3131), .B2(mem[2]), .ZN(
        n3055) );
  NAND2_X1 U2604 ( .A1(n1027), .A2(mem[770]), .ZN(n3054) );
  NAND4_X1 U2605 ( .A1(n3057), .A2(n3056), .A3(n3055), .A4(n3054), .ZN(n3058)
         );
  NOR3_X1 U2606 ( .A1(n3060), .A2(n3059), .A3(n3058), .ZN(n3074) );
  AOI22_X1 U2607 ( .A1(mem[674]), .A2(n3161), .B1(n3112), .B2(mem[386]), .ZN(
        n3065) );
  AOI22_X1 U2608 ( .A1(n1017), .A2(mem[194]), .B1(mem[98]), .B2(n1029), .ZN(
        n3064) );
  AOI22_X1 U2609 ( .A1(mem[610]), .A2(n3162), .B1(n3113), .B2(mem[546]), .ZN(
        n3063) );
  AOI22_X1 U2610 ( .A1(n3061), .A2(mem[642]), .B1(mem[162]), .B2(n3517), .ZN(
        n3062) );
  NAND4_X1 U2611 ( .A1(n3065), .A2(n3064), .A3(n3063), .A4(n3062), .ZN(n3072)
         );
  AOI22_X1 U2612 ( .A1(n3167), .A2(mem[514]), .B1(mem[930]), .B2(n3592), .ZN(
        n3070) );
  AOI22_X1 U2613 ( .A1(mem[962]), .A2(n1073), .B1(n1086), .B2(mem[738]), .ZN(
        n3069) );
  AOI22_X1 U2614 ( .A1(mem[866]), .A2(n3066), .B1(n3168), .B2(mem[802]), .ZN(
        n3068) );
  AOI22_X1 U2615 ( .A1(mem[898]), .A2(n3455), .B1(n1089), .B2(mem[834]), .ZN(
        n3067) );
  NAND4_X1 U2616 ( .A1(n3070), .A2(n3069), .A3(n3068), .A4(n3067), .ZN(n3071)
         );
  NOR2_X1 U2617 ( .A1(n3072), .A2(n3071), .ZN(n3073) );
  NAND2_X1 U2618 ( .A1(n3074), .A2(n3073), .ZN(rdata_a_o[2]) );
  AOI22_X1 U2619 ( .A1(mem[326]), .A2(n1005), .B1(n1085), .B2(mem[262]), .ZN(
        n3077) );
  AOI22_X1 U2620 ( .A1(mem[710]), .A2(n1082), .B1(n1013), .B2(mem[422]), .ZN(
        n3076) );
  AOI22_X1 U2621 ( .A1(mem[582]), .A2(n1015), .B1(n994), .B2(mem[454]), .ZN(
        n3080) );
  AOI22_X1 U2622 ( .A1(n1008), .A2(mem[230]), .B1(mem[134]), .B2(n1021), .ZN(
        n3079) );
  NAND2_X1 U2623 ( .A1(n3080), .A2(n3079), .ZN(n3086) );
  AOI22_X1 U2624 ( .A1(mem[358]), .A2(n1024), .B1(n3350), .B2(mem[294]), .ZN(
        n3084) );
  AOI22_X1 U2625 ( .A1(n1092), .A2(mem[486]), .B1(mem[38]), .B2(n4729), .ZN(
        n3083) );
  AOI22_X1 U2626 ( .A1(mem[70]), .A2(n3234), .B1(n3131), .B2(mem[6]), .ZN(
        n3082) );
  NAND2_X1 U2627 ( .A1(n1026), .A2(mem[774]), .ZN(n3081) );
  NAND4_X1 U2628 ( .A1(n3084), .A2(n3083), .A3(n3082), .A4(n3081), .ZN(n3085)
         );
  NOR3_X1 U2629 ( .A1(n3087), .A2(n3086), .A3(n3085), .ZN(n3099) );
  AOI22_X1 U2630 ( .A1(mem[678]), .A2(n3161), .B1(n3112), .B2(mem[390]), .ZN(
        n3091) );
  AOI22_X1 U2631 ( .A1(n1017), .A2(mem[198]), .B1(mem[102]), .B2(n4736), .ZN(
        n3090) );
  AOI22_X1 U2632 ( .A1(mem[614]), .A2(n3162), .B1(n3113), .B2(mem[550]), .ZN(
        n3089) );
  AOI22_X1 U2633 ( .A1(n3358), .A2(mem[646]), .B1(mem[166]), .B2(n3517), .ZN(
        n3088) );
  NAND4_X1 U2634 ( .A1(n3091), .A2(n3090), .A3(n3089), .A4(n3088), .ZN(n3098)
         );
  AOI22_X1 U2635 ( .A1(n3167), .A2(mem[518]), .B1(mem[934]), .B2(n3221), .ZN(
        n3096) );
  AOI22_X1 U2636 ( .A1(mem[966]), .A2(n1073), .B1(n1087), .B2(mem[742]), .ZN(
        n3095) );
  AOI22_X1 U2637 ( .A1(mem[870]), .A2(n3363), .B1(n3168), .B2(mem[806]), .ZN(
        n3094) );
  AOI22_X1 U2638 ( .A1(mem[902]), .A2(n3455), .B1(n1090), .B2(mem[838]), .ZN(
        n3093) );
  NAND4_X1 U2639 ( .A1(n3096), .A2(n3095), .A3(n3094), .A4(n3093), .ZN(n3097)
         );
  AOI22_X1 U2640 ( .A1(mem[327]), .A2(n1005), .B1(n1083), .B2(mem[263]), .ZN(
        n3101) );
  AOI22_X1 U2641 ( .A1(mem[711]), .A2(n1080), .B1(n1011), .B2(mem[423]), .ZN(
        n3100) );
  NAND2_X1 U2642 ( .A1(n3101), .A2(n3100), .ZN(n3111) );
  AOI22_X1 U2643 ( .A1(mem[583]), .A2(n1016), .B1(n996), .B2(mem[455]), .ZN(
        n3104) );
  AOI22_X1 U2644 ( .A1(n1009), .A2(mem[231]), .B1(mem[135]), .B2(n1021), .ZN(
        n3103) );
  NAND2_X1 U2645 ( .A1(n3104), .A2(n3103), .ZN(n3110) );
  AOI22_X1 U2646 ( .A1(mem[359]), .A2(n1024), .B1(n3350), .B2(mem[295]), .ZN(
        n3108) );
  AOI22_X1 U2647 ( .A1(n1093), .A2(mem[487]), .B1(mem[39]), .B2(n4729), .ZN(
        n3107) );
  AOI22_X1 U2648 ( .A1(mem[71]), .A2(n3234), .B1(n3131), .B2(mem[7]), .ZN(
        n3106) );
  NAND2_X1 U2649 ( .A1(n1025), .A2(mem[775]), .ZN(n3105) );
  NAND4_X1 U2650 ( .A1(n3108), .A2(n3107), .A3(n3106), .A4(n3105), .ZN(n3109)
         );
  NOR3_X1 U2651 ( .A1(n3111), .A2(n3110), .A3(n3109), .ZN(n3126) );
  AOI22_X1 U2652 ( .A1(mem[679]), .A2(n3161), .B1(n3112), .B2(mem[391]), .ZN(
        n3118) );
  AOI22_X1 U2653 ( .A1(n1019), .A2(mem[199]), .B1(mem[103]), .B2(n1031), .ZN(
        n3117) );
  AOI22_X1 U2654 ( .A1(mem[615]), .A2(n3162), .B1(n3113), .B2(mem[551]), .ZN(
        n3116) );
  AOI22_X1 U2655 ( .A1(n3358), .A2(mem[647]), .B1(mem[167]), .B2(n1072), .ZN(
        n3115) );
  NAND4_X1 U2656 ( .A1(n3118), .A2(n3117), .A3(n3116), .A4(n3115), .ZN(n3124)
         );
  AOI22_X1 U2657 ( .A1(n3167), .A2(mem[519]), .B1(mem[935]), .B2(n3221), .ZN(
        n3122) );
  AOI22_X1 U2658 ( .A1(mem[967]), .A2(n1073), .B1(n1086), .B2(mem[743]), .ZN(
        n3121) );
  AOI22_X1 U2659 ( .A1(mem[871]), .A2(n3363), .B1(n3168), .B2(mem[807]), .ZN(
        n3120) );
  AOI22_X1 U2660 ( .A1(mem[903]), .A2(n3594), .B1(n1089), .B2(mem[839]), .ZN(
        n3119) );
  NAND4_X1 U2661 ( .A1(n3119), .A2(n3121), .A3(n3120), .A4(n3122), .ZN(n3123)
         );
  NOR2_X1 U2662 ( .A1(n3124), .A2(n3123), .ZN(n3125) );
  NAND2_X1 U2663 ( .A1(n3126), .A2(n3125), .ZN(rdata_a_o[7]) );
  AOI22_X1 U2664 ( .A1(mem[328]), .A2(n1005), .B1(n1084), .B2(mem[264]), .ZN(
        n3128) );
  AOI22_X1 U2665 ( .A1(mem[712]), .A2(n1081), .B1(n1011), .B2(mem[424]), .ZN(
        n3127) );
  NAND2_X1 U2666 ( .A1(n3128), .A2(n3127), .ZN(n3138) );
  AOI22_X1 U2667 ( .A1(mem[584]), .A2(n1014), .B1(n994), .B2(mem[456]), .ZN(
        n3130) );
  AOI22_X1 U2668 ( .A1(n1010), .A2(mem[232]), .B1(mem[136]), .B2(n1022), .ZN(
        n3129) );
  NAND2_X1 U2669 ( .A1(n3130), .A2(n3129), .ZN(n3137) );
  AOI22_X1 U2670 ( .A1(mem[360]), .A2(n1023), .B1(n3350), .B2(mem[296]), .ZN(
        n3135) );
  AOI22_X1 U2671 ( .A1(n1067), .A2(mem[488]), .B1(mem[40]), .B2(n4729), .ZN(
        n3134) );
  AOI22_X1 U2672 ( .A1(mem[72]), .A2(n3234), .B1(n3351), .B2(mem[8]), .ZN(
        n3133) );
  NAND2_X1 U2673 ( .A1(n1027), .A2(mem[776]), .ZN(n3132) );
  NAND4_X1 U2674 ( .A1(n3135), .A2(n3134), .A3(n3133), .A4(n3132), .ZN(n3136)
         );
  NOR3_X1 U2675 ( .A1(n3136), .A2(n3137), .A3(n3138), .ZN(n3150) );
  AOI22_X1 U2676 ( .A1(mem[680]), .A2(n3161), .B1(n3382), .B2(mem[392]), .ZN(
        n3142) );
  AOI22_X1 U2677 ( .A1(n1018), .A2(mem[200]), .B1(mem[104]), .B2(n1029), .ZN(
        n3141) );
  AOI22_X1 U2678 ( .A1(mem[616]), .A2(n3162), .B1(n3383), .B2(mem[552]), .ZN(
        n3140) );
  AOI22_X1 U2679 ( .A1(n3358), .A2(mem[648]), .B1(mem[168]), .B2(n1072), .ZN(
        n3139) );
  NAND4_X1 U2680 ( .A1(n3142), .A2(n3141), .A3(n3140), .A4(n3139), .ZN(n3148)
         );
  AOI22_X1 U2681 ( .A1(n3167), .A2(mem[520]), .B1(mem[936]), .B2(n3221), .ZN(
        n3146) );
  AOI22_X1 U2682 ( .A1(mem[968]), .A2(n1073), .B1(n1087), .B2(mem[744]), .ZN(
        n3145) );
  AOI22_X1 U2683 ( .A1(mem[872]), .A2(n3363), .B1(n3168), .B2(mem[808]), .ZN(
        n3144) );
  AOI22_X1 U2684 ( .A1(mem[904]), .A2(n3455), .B1(n1090), .B2(mem[840]), .ZN(
        n3143) );
  NAND4_X1 U2685 ( .A1(n3146), .A2(n3145), .A3(n3144), .A4(n3143), .ZN(n3147)
         );
  NOR2_X1 U2686 ( .A1(n3148), .A2(n3147), .ZN(n3149) );
  NAND2_X1 U2687 ( .A1(n3150), .A2(n3149), .ZN(rdata_a_o[8]) );
  AOI22_X1 U2688 ( .A1(mem[329]), .A2(n1005), .B1(n1085), .B2(mem[265]), .ZN(
        n3152) );
  AOI22_X1 U2689 ( .A1(mem[713]), .A2(n1082), .B1(n1013), .B2(mem[425]), .ZN(
        n3151) );
  NAND2_X1 U2690 ( .A1(n3152), .A2(n3151), .ZN(n3160) );
  AOI22_X1 U2691 ( .A1(mem[585]), .A2(n1014), .B1(n995), .B2(mem[457]), .ZN(
        n3154) );
  AOI22_X1 U2692 ( .A1(n1010), .A2(mem[233]), .B1(mem[137]), .B2(n1022), .ZN(
        n3153) );
  NAND2_X1 U2693 ( .A1(n3154), .A2(n3153), .ZN(n3159) );
  AOI22_X1 U2694 ( .A1(mem[361]), .A2(n1024), .B1(n3350), .B2(mem[297]), .ZN(
        n3158) );
  AOI22_X1 U2695 ( .A1(n1067), .A2(mem[489]), .B1(mem[41]), .B2(n4730), .ZN(
        n3157) );
  AOI22_X1 U2696 ( .A1(mem[73]), .A2(n3234), .B1(n3351), .B2(mem[9]), .ZN(
        n3156) );
  NAND2_X1 U2697 ( .A1(n1027), .A2(mem[777]), .ZN(n3155) );
  AOI22_X1 U2698 ( .A1(mem[681]), .A2(n3161), .B1(n3382), .B2(mem[393]), .ZN(
        n3166) );
  AOI22_X1 U2699 ( .A1(n1018), .A2(mem[201]), .B1(mem[105]), .B2(n4736), .ZN(
        n3165) );
  AOI22_X1 U2700 ( .A1(mem[617]), .A2(n3162), .B1(n3383), .B2(mem[553]), .ZN(
        n3164) );
  AOI22_X1 U2701 ( .A1(n3358), .A2(mem[649]), .B1(mem[169]), .B2(n1072), .ZN(
        n3163) );
  NAND4_X1 U2702 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n3174)
         );
  AOI22_X1 U2703 ( .A1(n3167), .A2(mem[521]), .B1(mem[937]), .B2(n3221), .ZN(
        n3172) );
  AOI22_X1 U2704 ( .A1(mem[969]), .A2(n1073), .B1(n1086), .B2(mem[745]), .ZN(
        n3171) );
  AOI22_X1 U2705 ( .A1(mem[873]), .A2(n3363), .B1(n3168), .B2(mem[809]), .ZN(
        n3170) );
  AOI22_X1 U2706 ( .A1(mem[905]), .A2(n3594), .B1(n1089), .B2(mem[841]), .ZN(
        n3169) );
  NAND4_X1 U2707 ( .A1(n3172), .A2(n3171), .A3(n3170), .A4(n3169), .ZN(n3173)
         );
  NOR2_X1 U2708 ( .A1(n3174), .A2(n3173), .ZN(n3175) );
  AOI22_X1 U2709 ( .A1(mem[330]), .A2(n1007), .B1(n1085), .B2(mem[266]), .ZN(
        n3178) );
  AOI22_X1 U2710 ( .A1(mem[714]), .A2(n1080), .B1(n1012), .B2(mem[426]), .ZN(
        n3177) );
  NAND2_X1 U2711 ( .A1(n3178), .A2(n3177), .ZN(n3187) );
  AOI22_X1 U2712 ( .A1(mem[586]), .A2(n1015), .B1(n996), .B2(mem[458]), .ZN(
        n3180) );
  AOI22_X1 U2713 ( .A1(n1008), .A2(mem[234]), .B1(mem[138]), .B2(n1022), .ZN(
        n3179) );
  NAND2_X1 U2714 ( .A1(n3180), .A2(n3179), .ZN(n3186) );
  AOI22_X1 U2715 ( .A1(mem[362]), .A2(n1023), .B1(n3350), .B2(mem[298]), .ZN(
        n3184) );
  AOI22_X1 U2716 ( .A1(n1093), .A2(mem[490]), .B1(mem[42]), .B2(n4730), .ZN(
        n3183) );
  AOI22_X1 U2717 ( .A1(mem[74]), .A2(n3234), .B1(n3351), .B2(mem[10]), .ZN(
        n3182) );
  NAND2_X1 U2718 ( .A1(n1025), .A2(mem[778]), .ZN(n3181) );
  NAND4_X1 U2719 ( .A1(n3184), .A2(n3183), .A3(n3182), .A4(n3181), .ZN(n3185)
         );
  NOR3_X1 U2720 ( .A1(n3187), .A2(n3186), .A3(n3185), .ZN(n3204) );
  AOI22_X1 U2721 ( .A1(mem[682]), .A2(n1070), .B1(n3382), .B2(mem[394]), .ZN(
        n3193) );
  AOI22_X1 U2722 ( .A1(n1019), .A2(mem[202]), .B1(mem[106]), .B2(n1029), .ZN(
        n3192) );
  AOI22_X1 U2723 ( .A1(mem[618]), .A2(n1071), .B1(n3383), .B2(mem[554]), .ZN(
        n3191) );
  AOI22_X1 U2724 ( .A1(n3358), .A2(mem[650]), .B1(mem[170]), .B2(n1072), .ZN(
        n3190) );
  NAND4_X1 U2725 ( .A1(n3193), .A2(n3192), .A3(n3191), .A4(n3190), .ZN(n3202)
         );
  AOI22_X1 U2726 ( .A1(n1068), .A2(mem[522]), .B1(mem[938]), .B2(n3221), .ZN(
        n3200) );
  AOI22_X1 U2727 ( .A1(mem[970]), .A2(n1073), .B1(n1088), .B2(mem[746]), .ZN(
        n3199) );
  AOI22_X1 U2728 ( .A1(mem[874]), .A2(n3363), .B1(n1069), .B2(mem[810]), .ZN(
        n3198) );
  AOI22_X1 U2729 ( .A1(mem[906]), .A2(n3594), .B1(n1091), .B2(mem[842]), .ZN(
        n3197) );
  NAND4_X1 U2730 ( .A1(n3200), .A2(n3199), .A3(n3198), .A4(n3197), .ZN(n3201)
         );
  NOR2_X1 U2731 ( .A1(n3202), .A2(n3201), .ZN(n3203) );
  NAND2_X1 U2732 ( .A1(n3204), .A2(n3203), .ZN(rdata_a_o[10]) );
  AOI22_X1 U2733 ( .A1(mem[331]), .A2(n1007), .B1(n1083), .B2(mem[267]), .ZN(
        n3206) );
  AOI22_X1 U2734 ( .A1(mem[715]), .A2(n1080), .B1(n1012), .B2(mem[427]), .ZN(
        n3205) );
  AOI22_X1 U2735 ( .A1(mem[587]), .A2(n1014), .B1(n994), .B2(mem[459]), .ZN(
        n3209) );
  AOI22_X1 U2736 ( .A1(n1008), .A2(mem[235]), .B1(mem[139]), .B2(n1020), .ZN(
        n3208) );
  NAND2_X1 U2737 ( .A1(n3209), .A2(n3208), .ZN(n3216) );
  AOI22_X1 U2738 ( .A1(mem[363]), .A2(n1023), .B1(n3350), .B2(mem[299]), .ZN(
        n3214) );
  AOI22_X1 U2739 ( .A1(n1093), .A2(mem[491]), .B1(mem[43]), .B2(n4729), .ZN(
        n3213) );
  AOI22_X1 U2740 ( .A1(mem[75]), .A2(n3234), .B1(n3351), .B2(mem[11]), .ZN(
        n3212) );
  NAND2_X1 U2741 ( .A1(n1026), .A2(mem[779]), .ZN(n3211) );
  NAND4_X1 U2742 ( .A1(n3214), .A2(n3213), .A3(n3212), .A4(n3211), .ZN(n3215)
         );
  AOI22_X1 U2743 ( .A1(mem[683]), .A2(n1070), .B1(n3382), .B2(mem[395]), .ZN(
        n3220) );
  AOI22_X1 U2744 ( .A1(n1019), .A2(mem[203]), .B1(mem[107]), .B2(n1029), .ZN(
        n3219) );
  AOI22_X1 U2745 ( .A1(mem[619]), .A2(n1071), .B1(n3383), .B2(mem[555]), .ZN(
        n3218) );
  AOI22_X1 U2746 ( .A1(n3358), .A2(mem[651]), .B1(mem[171]), .B2(n1072), .ZN(
        n3217) );
  NAND4_X1 U2747 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .ZN(n3228)
         );
  AOI22_X1 U2748 ( .A1(n1068), .A2(mem[523]), .B1(mem[939]), .B2(n3221), .ZN(
        n3226) );
  AOI22_X1 U2749 ( .A1(mem[971]), .A2(n1073), .B1(n1088), .B2(mem[747]), .ZN(
        n3225) );
  AOI22_X1 U2750 ( .A1(mem[875]), .A2(n3363), .B1(n1069), .B2(mem[811]), .ZN(
        n3224) );
  AOI22_X1 U2751 ( .A1(mem[907]), .A2(n3269), .B1(n1091), .B2(mem[843]), .ZN(
        n3223) );
  NAND4_X1 U2752 ( .A1(n3226), .A2(n3225), .A3(n3224), .A4(n3223), .ZN(n3227)
         );
  NOR2_X1 U2753 ( .A1(n3228), .A2(n3227), .ZN(n3229) );
  AOI22_X1 U2754 ( .A1(mem[332]), .A2(n1006), .B1(n1083), .B2(mem[268]), .ZN(
        n3231) );
  AOI22_X1 U2755 ( .A1(mem[716]), .A2(n1081), .B1(n1013), .B2(mem[428]), .ZN(
        n3230) );
  NAND2_X1 U2756 ( .A1(n3231), .A2(n3230), .ZN(n3241) );
  AOI22_X1 U2757 ( .A1(mem[588]), .A2(n1015), .B1(n994), .B2(mem[460]), .ZN(
        n3233) );
  AOI22_X1 U2758 ( .A1(n1009), .A2(mem[236]), .B1(mem[140]), .B2(n1021), .ZN(
        n3232) );
  NAND2_X1 U2759 ( .A1(n3233), .A2(n3232), .ZN(n3240) );
  AOI22_X1 U2760 ( .A1(mem[364]), .A2(n1024), .B1(n3350), .B2(mem[300]), .ZN(
        n3238) );
  AOI22_X1 U2761 ( .A1(n1067), .A2(mem[492]), .B1(mem[44]), .B2(n4729), .ZN(
        n3237) );
  AOI22_X1 U2762 ( .A1(mem[76]), .A2(n3234), .B1(n3351), .B2(mem[12]), .ZN(
        n3236) );
  NAND2_X1 U2763 ( .A1(n1025), .A2(mem[780]), .ZN(n3235) );
  NAND4_X1 U2764 ( .A1(n3238), .A2(n3237), .A3(n3236), .A4(n3235), .ZN(n3239)
         );
  NOR3_X1 U2765 ( .A1(n3241), .A2(n3240), .A3(n3239), .ZN(n3253) );
  AOI22_X1 U2766 ( .A1(mem[684]), .A2(n1070), .B1(n3382), .B2(mem[396]), .ZN(
        n3245) );
  AOI22_X1 U2767 ( .A1(n1018), .A2(mem[204]), .B1(mem[108]), .B2(n4736), .ZN(
        n3244) );
  AOI22_X1 U2768 ( .A1(mem[620]), .A2(n1071), .B1(n3383), .B2(mem[556]), .ZN(
        n3243) );
  AOI22_X1 U2769 ( .A1(n3358), .A2(mem[652]), .B1(mem[172]), .B2(n1072), .ZN(
        n3242) );
  NAND4_X1 U2770 ( .A1(n3245), .A2(n3244), .A3(n3243), .A4(n3242), .ZN(n3251)
         );
  AOI22_X1 U2771 ( .A1(n1068), .A2(mem[524]), .B1(mem[940]), .B2(n3433), .ZN(
        n3249) );
  AOI22_X1 U2772 ( .A1(mem[972]), .A2(n1073), .B1(n1088), .B2(mem[748]), .ZN(
        n3248) );
  AOI22_X1 U2773 ( .A1(mem[876]), .A2(n3363), .B1(n1069), .B2(mem[812]), .ZN(
        n3247) );
  AOI22_X1 U2774 ( .A1(mem[908]), .A2(n3594), .B1(n1091), .B2(mem[844]), .ZN(
        n3246) );
  NAND4_X1 U2775 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3250)
         );
  NOR2_X1 U2776 ( .A1(n3251), .A2(n3250), .ZN(n3252) );
  NAND2_X1 U2777 ( .A1(n3253), .A2(n3252), .ZN(rdata_a_o[12]) );
  AOI22_X1 U2778 ( .A1(mem[333]), .A2(n1005), .B1(n1084), .B2(mem[269]), .ZN(
        n3255) );
  AOI22_X1 U2779 ( .A1(mem[717]), .A2(n1082), .B1(n1012), .B2(mem[429]), .ZN(
        n3254) );
  NAND2_X1 U2780 ( .A1(n3255), .A2(n3254), .ZN(n3264) );
  AOI22_X1 U2781 ( .A1(mem[589]), .A2(n1016), .B1(n996), .B2(mem[461]), .ZN(
        n3257) );
  AOI22_X1 U2782 ( .A1(n1008), .A2(mem[237]), .B1(mem[141]), .B2(n1020), .ZN(
        n3256) );
  NAND2_X1 U2783 ( .A1(n3257), .A2(n3256), .ZN(n3263) );
  AOI22_X1 U2784 ( .A1(mem[365]), .A2(n1023), .B1(n3350), .B2(mem[301]), .ZN(
        n3261) );
  AOI22_X1 U2785 ( .A1(n1067), .A2(mem[493]), .B1(mem[45]), .B2(n4730), .ZN(
        n3260) );
  AOI22_X1 U2786 ( .A1(mem[77]), .A2(n3512), .B1(n3351), .B2(mem[13]), .ZN(
        n3259) );
  NAND2_X1 U2787 ( .A1(n1027), .A2(mem[781]), .ZN(n3258) );
  NAND4_X1 U2788 ( .A1(n3261), .A2(n3260), .A3(n3259), .A4(n3258), .ZN(n3262)
         );
  NOR3_X1 U2789 ( .A1(n3264), .A2(n3263), .A3(n3262), .ZN(n3277) );
  AOI22_X1 U2790 ( .A1(mem[685]), .A2(n1070), .B1(n3382), .B2(mem[397]), .ZN(
        n3268) );
  AOI22_X1 U2791 ( .A1(n1017), .A2(mem[205]), .B1(mem[109]), .B2(n1029), .ZN(
        n3267) );
  AOI22_X1 U2792 ( .A1(mem[621]), .A2(n1071), .B1(n3383), .B2(mem[557]), .ZN(
        n3266) );
  AOI22_X1 U2793 ( .A1(n3358), .A2(mem[653]), .B1(mem[173]), .B2(n1072), .ZN(
        n3265) );
  NAND4_X1 U2794 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3275)
         );
  AOI22_X1 U2795 ( .A1(n1068), .A2(mem[525]), .B1(mem[941]), .B2(n3433), .ZN(
        n3273) );
  AOI22_X1 U2796 ( .A1(mem[973]), .A2(n1073), .B1(n1087), .B2(mem[749]), .ZN(
        n3272) );
  AOI22_X1 U2797 ( .A1(mem[877]), .A2(n3363), .B1(n1069), .B2(mem[813]), .ZN(
        n3271) );
  AOI22_X1 U2798 ( .A1(mem[909]), .A2(n3455), .B1(n1090), .B2(mem[845]), .ZN(
        n3270) );
  NAND4_X1 U2799 ( .A1(n3273), .A2(n3272), .A3(n3271), .A4(n3270), .ZN(n3274)
         );
  NOR2_X1 U2800 ( .A1(n3275), .A2(n3274), .ZN(n3276) );
  NAND2_X1 U2801 ( .A1(n3277), .A2(n3276), .ZN(rdata_a_o[13]) );
  AOI22_X1 U2802 ( .A1(mem[334]), .A2(n1006), .B1(n1083), .B2(mem[270]), .ZN(
        n3279) );
  AOI22_X1 U2803 ( .A1(mem[718]), .A2(n1082), .B1(n1012), .B2(mem[430]), .ZN(
        n3278) );
  NAND2_X1 U2804 ( .A1(n3279), .A2(n3278), .ZN(n3288) );
  AOI22_X1 U2805 ( .A1(mem[590]), .A2(n1016), .B1(n996), .B2(mem[462]), .ZN(
        n3281) );
  AOI22_X1 U2806 ( .A1(n1009), .A2(mem[238]), .B1(mem[142]), .B2(n1021), .ZN(
        n3280) );
  NAND2_X1 U2807 ( .A1(n3281), .A2(n3280), .ZN(n3287) );
  AOI22_X1 U2808 ( .A1(mem[366]), .A2(n1023), .B1(n3350), .B2(mem[302]), .ZN(
        n3285) );
  AOI22_X1 U2809 ( .A1(n1092), .A2(mem[494]), .B1(mem[46]), .B2(n4730), .ZN(
        n3284) );
  AOI22_X1 U2810 ( .A1(mem[78]), .A2(n3512), .B1(n3351), .B2(mem[14]), .ZN(
        n3283) );
  NAND2_X1 U2811 ( .A1(n1027), .A2(mem[782]), .ZN(n3282) );
  NAND4_X1 U2812 ( .A1(n3285), .A2(n3284), .A3(n3283), .A4(n3282), .ZN(n3286)
         );
  NOR3_X1 U2813 ( .A1(n3288), .A2(n3287), .A3(n3286), .ZN(n3300) );
  AOI22_X1 U2814 ( .A1(mem[686]), .A2(n1070), .B1(n3382), .B2(mem[398]), .ZN(
        n3292) );
  AOI22_X1 U2815 ( .A1(n1018), .A2(mem[206]), .B1(mem[110]), .B2(n1029), .ZN(
        n3291) );
  AOI22_X1 U2816 ( .A1(mem[622]), .A2(n1071), .B1(n3383), .B2(mem[558]), .ZN(
        n3290) );
  AOI22_X1 U2817 ( .A1(n3358), .A2(mem[654]), .B1(mem[174]), .B2(n1072), .ZN(
        n3289) );
  NAND4_X1 U2818 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3298)
         );
  AOI22_X1 U2819 ( .A1(n1068), .A2(mem[526]), .B1(mem[942]), .B2(n3433), .ZN(
        n3296) );
  AOI22_X1 U2820 ( .A1(mem[974]), .A2(n3564), .B1(n1086), .B2(mem[750]), .ZN(
        n3295) );
  AOI22_X1 U2821 ( .A1(mem[878]), .A2(n3363), .B1(n1069), .B2(mem[814]), .ZN(
        n3294) );
  AOI22_X1 U2822 ( .A1(mem[910]), .A2(n3455), .B1(n1089), .B2(mem[846]), .ZN(
        n3293) );
  NAND4_X1 U2823 ( .A1(n3296), .A2(n3295), .A3(n3294), .A4(n3293), .ZN(n3297)
         );
  NOR2_X1 U2824 ( .A1(n3298), .A2(n3297), .ZN(n3299) );
  NAND2_X1 U2825 ( .A1(n3300), .A2(n3299), .ZN(rdata_a_o[14]) );
  AOI22_X1 U2826 ( .A1(mem[335]), .A2(n1007), .B1(n1085), .B2(mem[271]), .ZN(
        n3302) );
  AOI22_X1 U2827 ( .A1(mem[719]), .A2(n1081), .B1(n1011), .B2(mem[431]), .ZN(
        n3301) );
  NAND2_X1 U2828 ( .A1(n3302), .A2(n3301), .ZN(n3311) );
  AOI22_X1 U2829 ( .A1(mem[591]), .A2(n1014), .B1(n995), .B2(mem[463]), .ZN(
        n3304) );
  AOI22_X1 U2830 ( .A1(n1010), .A2(mem[239]), .B1(mem[143]), .B2(n1020), .ZN(
        n3303) );
  NAND2_X1 U2831 ( .A1(n3304), .A2(n3303), .ZN(n3310) );
  AOI22_X1 U2832 ( .A1(mem[367]), .A2(n1023), .B1(n3350), .B2(mem[303]), .ZN(
        n3308) );
  AOI22_X1 U2833 ( .A1(n1067), .A2(mem[495]), .B1(mem[47]), .B2(n4730), .ZN(
        n3307) );
  AOI22_X1 U2834 ( .A1(mem[79]), .A2(n3512), .B1(n3351), .B2(mem[15]), .ZN(
        n3306) );
  NAND2_X1 U2835 ( .A1(n1026), .A2(mem[783]), .ZN(n3305) );
  NAND4_X1 U2836 ( .A1(n3308), .A2(n3307), .A3(n3306), .A4(n3305), .ZN(n3309)
         );
  NOR3_X1 U2837 ( .A1(n3311), .A2(n3310), .A3(n3309), .ZN(n3323) );
  AOI22_X1 U2838 ( .A1(mem[687]), .A2(n1070), .B1(n3382), .B2(mem[399]), .ZN(
        n3315) );
  AOI22_X1 U2839 ( .A1(n1017), .A2(mem[207]), .B1(mem[111]), .B2(n4736), .ZN(
        n3314) );
  AOI22_X1 U2840 ( .A1(mem[623]), .A2(n1071), .B1(n3383), .B2(mem[559]), .ZN(
        n3313) );
  AOI22_X1 U2841 ( .A1(n3358), .A2(mem[655]), .B1(mem[175]), .B2(n1072), .ZN(
        n3312) );
  NAND4_X1 U2842 ( .A1(n3315), .A2(n3314), .A3(n3313), .A4(n3312), .ZN(n3321)
         );
  AOI22_X1 U2843 ( .A1(n1068), .A2(mem[527]), .B1(mem[943]), .B2(n3433), .ZN(
        n3319) );
  AOI22_X1 U2844 ( .A1(mem[975]), .A2(n3564), .B1(n1088), .B2(mem[751]), .ZN(
        n3318) );
  AOI22_X1 U2845 ( .A1(mem[879]), .A2(n3363), .B1(n1069), .B2(mem[815]), .ZN(
        n3317) );
  AOI22_X1 U2846 ( .A1(mem[911]), .A2(n3455), .B1(n1091), .B2(mem[847]), .ZN(
        n3316) );
  NAND4_X1 U2847 ( .A1(n3319), .A2(n3318), .A3(n3317), .A4(n3316), .ZN(n3320)
         );
  NOR2_X1 U2848 ( .A1(n3321), .A2(n3320), .ZN(n3322) );
  NAND2_X1 U2849 ( .A1(n3323), .A2(n3322), .ZN(rdata_a_o[15]) );
  AOI22_X1 U2850 ( .A1(mem[592]), .A2(n1015), .B1(n996), .B2(mem[464]), .ZN(
        n3327) );
  AOI22_X1 U2851 ( .A1(mem[336]), .A2(n1005), .B1(n1085), .B2(mem[272]), .ZN(
        n3326) );
  AOI22_X1 U2852 ( .A1(mem[720]), .A2(n1081), .B1(n1012), .B2(mem[432]), .ZN(
        n3325) );
  AOI22_X1 U2853 ( .A1(n1009), .A2(mem[240]), .B1(mem[144]), .B2(n1021), .ZN(
        n3324) );
  NAND4_X1 U2854 ( .A1(n3327), .A2(n3326), .A3(n3325), .A4(n3324), .ZN(n3333)
         );
  AOI22_X1 U2855 ( .A1(mem[368]), .A2(n1024), .B1(n3350), .B2(mem[304]), .ZN(
        n3331) );
  AOI22_X1 U2856 ( .A1(n1067), .A2(mem[496]), .B1(mem[48]), .B2(n4729), .ZN(
        n3330) );
  AOI22_X1 U2857 ( .A1(mem[80]), .A2(n3512), .B1(n3351), .B2(mem[16]), .ZN(
        n3329) );
  NAND2_X1 U2858 ( .A1(n1025), .A2(mem[784]), .ZN(n3328) );
  NAND4_X1 U2859 ( .A1(n3331), .A2(n3330), .A3(n3329), .A4(n3328), .ZN(n3332)
         );
  NOR2_X1 U2860 ( .A1(n3333), .A2(n3332), .ZN(n3345) );
  AOI22_X1 U2861 ( .A1(mem[688]), .A2(n1070), .B1(n3382), .B2(mem[400]), .ZN(
        n3337) );
  AOI22_X1 U2862 ( .A1(n1018), .A2(mem[208]), .B1(mem[112]), .B2(n1031), .ZN(
        n3336) );
  AOI22_X1 U2863 ( .A1(mem[624]), .A2(n1071), .B1(n3383), .B2(mem[560]), .ZN(
        n3335) );
  AOI22_X1 U2864 ( .A1(n3358), .A2(mem[656]), .B1(mem[176]), .B2(n3517), .ZN(
        n3334) );
  NAND4_X1 U2865 ( .A1(n3337), .A2(n3336), .A3(n3335), .A4(n3334), .ZN(n3343)
         );
  AOI22_X1 U2866 ( .A1(n1068), .A2(mem[528]), .B1(mem[944]), .B2(n3433), .ZN(
        n3341) );
  AOI22_X1 U2867 ( .A1(mem[976]), .A2(n3564), .B1(n1086), .B2(mem[752]), .ZN(
        n3340) );
  AOI22_X1 U2868 ( .A1(mem[880]), .A2(n3363), .B1(n1069), .B2(mem[816]), .ZN(
        n3339) );
  AOI22_X1 U2869 ( .A1(mem[912]), .A2(n3455), .B1(n1089), .B2(mem[848]), .ZN(
        n3338) );
  NAND4_X1 U2870 ( .A1(n3341), .A2(n3340), .A3(n3339), .A4(n3338), .ZN(n3342)
         );
  NOR2_X1 U2871 ( .A1(n3343), .A2(n3342), .ZN(n3344) );
  NAND2_X1 U2872 ( .A1(n3345), .A2(n3344), .ZN(rdata_a_o[16]) );
  AOI22_X1 U2873 ( .A1(mem[593]), .A2(n1014), .B1(n995), .B2(mem[465]), .ZN(
        n3349) );
  AOI22_X1 U2874 ( .A1(mem[337]), .A2(n1007), .B1(n1084), .B2(mem[273]), .ZN(
        n3348) );
  AOI22_X1 U2875 ( .A1(mem[721]), .A2(n1081), .B1(n1011), .B2(mem[433]), .ZN(
        n3347) );
  AOI22_X1 U2876 ( .A1(n1008), .A2(mem[241]), .B1(mem[145]), .B2(n1020), .ZN(
        n3346) );
  NAND4_X1 U2877 ( .A1(n3349), .A2(n3348), .A3(n3347), .A4(n3346), .ZN(n3357)
         );
  AOI22_X1 U2878 ( .A1(mem[369]), .A2(n1023), .B1(n3350), .B2(mem[305]), .ZN(
        n3355) );
  AOI22_X1 U2879 ( .A1(n1092), .A2(mem[497]), .B1(mem[49]), .B2(n4729), .ZN(
        n3354) );
  AOI22_X1 U2880 ( .A1(mem[81]), .A2(n3512), .B1(n3351), .B2(mem[17]), .ZN(
        n3353) );
  NAND2_X1 U2881 ( .A1(n1026), .A2(mem[785]), .ZN(n3352) );
  NAND4_X1 U2882 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3356)
         );
  NOR2_X1 U2883 ( .A1(n3357), .A2(n3356), .ZN(n3371) );
  AOI22_X1 U2884 ( .A1(mem[689]), .A2(n1070), .B1(n3382), .B2(mem[401]), .ZN(
        n3362) );
  AOI22_X1 U2885 ( .A1(n1017), .A2(mem[209]), .B1(mem[113]), .B2(n4736), .ZN(
        n3361) );
  AOI22_X1 U2886 ( .A1(mem[625]), .A2(n1071), .B1(n3383), .B2(mem[561]), .ZN(
        n3360) );
  AOI22_X1 U2887 ( .A1(n3358), .A2(mem[657]), .B1(mem[177]), .B2(n3517), .ZN(
        n3359) );
  NAND4_X1 U2888 ( .A1(n3362), .A2(n3361), .A3(n3360), .A4(n3359), .ZN(n3369)
         );
  AOI22_X1 U2889 ( .A1(n1068), .A2(mem[529]), .B1(mem[945]), .B2(n3433), .ZN(
        n3367) );
  AOI22_X1 U2890 ( .A1(mem[977]), .A2(n3564), .B1(n1087), .B2(mem[753]), .ZN(
        n3366) );
  AOI22_X1 U2891 ( .A1(mem[881]), .A2(n3363), .B1(n1069), .B2(mem[817]), .ZN(
        n3365) );
  AOI22_X1 U2892 ( .A1(mem[913]), .A2(n3594), .B1(n1091), .B2(mem[849]), .ZN(
        n3364) );
  NAND4_X1 U2893 ( .A1(n3367), .A2(n3366), .A3(n3365), .A4(n3364), .ZN(n3368)
         );
  NOR2_X1 U2894 ( .A1(n3369), .A2(n3368), .ZN(n3370) );
  NAND2_X1 U2895 ( .A1(n3371), .A2(n3370), .ZN(rdata_a_o[17]) );
  AOI22_X1 U2896 ( .A1(mem[594]), .A2(n1014), .B1(n995), .B2(mem[466]), .ZN(
        n3375) );
  AOI22_X1 U2897 ( .A1(mem[338]), .A2(n1006), .B1(n1084), .B2(mem[274]), .ZN(
        n3374) );
  AOI22_X1 U2898 ( .A1(mem[722]), .A2(n1080), .B1(n1013), .B2(mem[434]), .ZN(
        n3373) );
  AOI22_X1 U2899 ( .A1(n1010), .A2(mem[242]), .B1(mem[146]), .B2(n1022), .ZN(
        n3372) );
  NAND4_X1 U2900 ( .A1(n3375), .A2(n3374), .A3(n3373), .A4(n3372), .ZN(n3381)
         );
  AOI22_X1 U2901 ( .A1(mem[370]), .A2(n2161), .B1(n3577), .B2(mem[306]), .ZN(
        n3379) );
  AOI22_X1 U2902 ( .A1(n1067), .A2(mem[498]), .B1(mem[50]), .B2(n4730), .ZN(
        n3378) );
  AOI22_X1 U2903 ( .A1(mem[82]), .A2(n3512), .B1(n3578), .B2(mem[18]), .ZN(
        n3377) );
  NAND2_X1 U2904 ( .A1(n1026), .A2(mem[786]), .ZN(n3376) );
  NAND4_X1 U2905 ( .A1(n3379), .A2(n3378), .A3(n3377), .A4(n3376), .ZN(n3380)
         );
  NOR2_X1 U2906 ( .A1(n3381), .A2(n3380), .ZN(n3395) );
  AOI22_X1 U2907 ( .A1(mem[690]), .A2(n1070), .B1(n3382), .B2(mem[402]), .ZN(
        n3387) );
  AOI22_X1 U2908 ( .A1(n1019), .A2(mem[210]), .B1(mem[114]), .B2(n4736), .ZN(
        n3386) );
  AOI22_X1 U2909 ( .A1(mem[626]), .A2(n1071), .B1(n3383), .B2(mem[562]), .ZN(
        n3385) );
  AOI22_X1 U2910 ( .A1(n3587), .A2(mem[658]), .B1(mem[178]), .B2(n3517), .ZN(
        n3384) );
  NAND4_X1 U2911 ( .A1(n3387), .A2(n3386), .A3(n3385), .A4(n3384), .ZN(n3393)
         );
  AOI22_X1 U2912 ( .A1(n1068), .A2(mem[530]), .B1(mem[946]), .B2(n3433), .ZN(
        n3391) );
  AOI22_X1 U2913 ( .A1(mem[978]), .A2(n3564), .B1(n1087), .B2(mem[754]), .ZN(
        n3390) );
  AOI22_X1 U2914 ( .A1(mem[882]), .A2(n3593), .B1(n1069), .B2(mem[818]), .ZN(
        n3389) );
  AOI22_X1 U2915 ( .A1(mem[914]), .A2(n3594), .B1(n1090), .B2(mem[850]), .ZN(
        n3388) );
  NAND4_X1 U2916 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(n3392)
         );
  NOR2_X1 U2917 ( .A1(n3393), .A2(n3392), .ZN(n3394) );
  NAND2_X1 U2918 ( .A1(n3395), .A2(n3394), .ZN(rdata_a_o[18]) );
  AOI22_X1 U2919 ( .A1(mem[595]), .A2(n1016), .B1(n996), .B2(mem[467]), .ZN(
        n3399) );
  AOI22_X1 U2920 ( .A1(mem[339]), .A2(n1006), .B1(n1085), .B2(mem[275]), .ZN(
        n3398) );
  AOI22_X1 U2921 ( .A1(mem[723]), .A2(n1080), .B1(n1011), .B2(mem[435]), .ZN(
        n3397) );
  AOI22_X1 U2922 ( .A1(n1008), .A2(mem[243]), .B1(mem[147]), .B2(n1020), .ZN(
        n3396) );
  NAND4_X1 U2923 ( .A1(n3399), .A2(n3398), .A3(n3397), .A4(n3396), .ZN(n3405)
         );
  AOI22_X1 U2924 ( .A1(mem[371]), .A2(n1024), .B1(n3577), .B2(mem[307]), .ZN(
        n3403) );
  AOI22_X1 U2925 ( .A1(n1093), .A2(mem[499]), .B1(mem[51]), .B2(n4730), .ZN(
        n3402) );
  AOI22_X1 U2926 ( .A1(mem[83]), .A2(n3512), .B1(n3578), .B2(mem[19]), .ZN(
        n3401) );
  NAND2_X1 U2927 ( .A1(n1026), .A2(mem[787]), .ZN(n3400) );
  NAND4_X1 U2928 ( .A1(n3403), .A2(n3402), .A3(n3401), .A4(n3400), .ZN(n3404)
         );
  NOR2_X1 U2929 ( .A1(n3405), .A2(n3404), .ZN(n3417) );
  AOI22_X1 U2930 ( .A1(mem[691]), .A2(n1070), .B1(n3585), .B2(mem[403]), .ZN(
        n3409) );
  AOI22_X1 U2931 ( .A1(n1018), .A2(mem[211]), .B1(mem[115]), .B2(n1031), .ZN(
        n3408) );
  AOI22_X1 U2932 ( .A1(mem[627]), .A2(n1071), .B1(n3586), .B2(mem[563]), .ZN(
        n3407) );
  AOI22_X1 U2933 ( .A1(n3587), .A2(mem[659]), .B1(mem[179]), .B2(n3517), .ZN(
        n3406) );
  NAND4_X1 U2934 ( .A1(n3409), .A2(n3408), .A3(n3407), .A4(n3406), .ZN(n3415)
         );
  AOI22_X1 U2935 ( .A1(n1068), .A2(mem[531]), .B1(mem[947]), .B2(n3433), .ZN(
        n3413) );
  AOI22_X1 U2936 ( .A1(mem[979]), .A2(n3564), .B1(n1086), .B2(mem[755]), .ZN(
        n3412) );
  AOI22_X1 U2937 ( .A1(mem[883]), .A2(n3593), .B1(n1069), .B2(mem[819]), .ZN(
        n3411) );
  AOI22_X1 U2938 ( .A1(mem[915]), .A2(n3594), .B1(n1089), .B2(mem[851]), .ZN(
        n3410) );
  NAND2_X1 U2939 ( .A1(n3417), .A2(n3416), .ZN(rdata_a_o[19]) );
  AOI22_X1 U2940 ( .A1(mem[596]), .A2(n1014), .B1(n994), .B2(mem[468]), .ZN(
        n3421) );
  AOI22_X1 U2941 ( .A1(mem[340]), .A2(n1005), .B1(n1083), .B2(mem[276]), .ZN(
        n3420) );
  AOI22_X1 U2942 ( .A1(mem[724]), .A2(n1080), .B1(n1011), .B2(mem[436]), .ZN(
        n3419) );
  AOI22_X1 U2943 ( .A1(n1008), .A2(mem[244]), .B1(mem[148]), .B2(n1020), .ZN(
        n3418) );
  NAND4_X1 U2944 ( .A1(n3421), .A2(n3420), .A3(n3419), .A4(n3418), .ZN(n3428)
         );
  AOI22_X1 U2945 ( .A1(mem[372]), .A2(n1024), .B1(n3577), .B2(mem[308]), .ZN(
        n3426) );
  AOI22_X1 U2946 ( .A1(n1092), .A2(mem[500]), .B1(mem[52]), .B2(n4730), .ZN(
        n3425) );
  AOI22_X1 U2947 ( .A1(mem[84]), .A2(n3512), .B1(n3578), .B2(mem[20]), .ZN(
        n3424) );
  NAND2_X1 U2948 ( .A1(n1027), .A2(mem[788]), .ZN(n3423) );
  NAND4_X1 U2949 ( .A1(n3426), .A2(n3425), .A3(n3424), .A4(n3423), .ZN(n3427)
         );
  NOR2_X1 U2950 ( .A1(n3428), .A2(n3427), .ZN(n3441) );
  AOI22_X1 U2951 ( .A1(mem[692]), .A2(n1070), .B1(n3585), .B2(mem[404]), .ZN(
        n3432) );
  AOI22_X1 U2952 ( .A1(n1017), .A2(mem[212]), .B1(mem[116]), .B2(n1029), .ZN(
        n3431) );
  AOI22_X1 U2953 ( .A1(mem[628]), .A2(n1071), .B1(n3586), .B2(mem[564]), .ZN(
        n3430) );
  AOI22_X1 U2954 ( .A1(n3587), .A2(mem[660]), .B1(mem[180]), .B2(n3517), .ZN(
        n3429) );
  NAND4_X1 U2955 ( .A1(n3432), .A2(n3431), .A3(n3430), .A4(n3429), .ZN(n3439)
         );
  AOI22_X1 U2956 ( .A1(n1068), .A2(mem[532]), .B1(mem[948]), .B2(n3433), .ZN(
        n3437) );
  AOI22_X1 U2957 ( .A1(mem[980]), .A2(n3564), .B1(n1086), .B2(mem[756]), .ZN(
        n3436) );
  AOI22_X1 U2958 ( .A1(mem[884]), .A2(n3593), .B1(n1069), .B2(mem[820]), .ZN(
        n3435) );
  AOI22_X1 U2959 ( .A1(mem[916]), .A2(n3455), .B1(n1090), .B2(mem[852]), .ZN(
        n3434) );
  NAND4_X1 U2960 ( .A1(n3437), .A2(n3436), .A3(n3435), .A4(n3434), .ZN(n3438)
         );
  NOR2_X1 U2961 ( .A1(n3439), .A2(n3438), .ZN(n3440) );
  NAND2_X1 U2962 ( .A1(n3441), .A2(n3440), .ZN(rdata_a_o[20]) );
  AOI22_X1 U2963 ( .A1(mem[597]), .A2(n1016), .B1(n996), .B2(mem[469]), .ZN(
        n3445) );
  AOI22_X1 U2964 ( .A1(mem[341]), .A2(n1007), .B1(n1085), .B2(mem[277]), .ZN(
        n3444) );
  AOI22_X1 U2965 ( .A1(mem[725]), .A2(n1082), .B1(n1011), .B2(mem[437]), .ZN(
        n3443) );
  AOI22_X1 U2966 ( .A1(n1010), .A2(mem[245]), .B1(mem[149]), .B2(n1022), .ZN(
        n3442) );
  AOI22_X1 U2967 ( .A1(mem[373]), .A2(n1023), .B1(n3577), .B2(mem[309]), .ZN(
        n3449) );
  AOI22_X1 U2968 ( .A1(n1093), .A2(mem[501]), .B1(mem[53]), .B2(n4730), .ZN(
        n3448) );
  AOI22_X1 U2969 ( .A1(mem[85]), .A2(n3579), .B1(n3578), .B2(mem[21]), .ZN(
        n3447) );
  NAND2_X1 U2970 ( .A1(n1025), .A2(mem[789]), .ZN(n3446) );
  NAND4_X1 U2971 ( .A1(n3449), .A2(n3448), .A3(n3447), .A4(n3446), .ZN(n3450)
         );
  AOI22_X1 U2972 ( .A1(mem[693]), .A2(n1070), .B1(n3585), .B2(mem[405]), .ZN(
        n3454) );
  AOI22_X1 U2973 ( .A1(n1018), .A2(mem[213]), .B1(mem[117]), .B2(n1029), .ZN(
        n3453) );
  AOI22_X1 U2974 ( .A1(mem[629]), .A2(n1071), .B1(n3586), .B2(mem[565]), .ZN(
        n3452) );
  AOI22_X1 U2975 ( .A1(n3587), .A2(mem[661]), .B1(mem[181]), .B2(n3517), .ZN(
        n3451) );
  NAND4_X1 U2976 ( .A1(n3454), .A2(n3453), .A3(n3452), .A4(n3451), .ZN(n3461)
         );
  AOI22_X1 U2977 ( .A1(n1068), .A2(mem[533]), .B1(mem[949]), .B2(n3592), .ZN(
        n3459) );
  AOI22_X1 U2978 ( .A1(mem[981]), .A2(n3564), .B1(n1088), .B2(mem[757]), .ZN(
        n3458) );
  AOI22_X1 U2979 ( .A1(mem[885]), .A2(n3593), .B1(n1069), .B2(mem[821]), .ZN(
        n3457) );
  AOI22_X1 U2980 ( .A1(mem[917]), .A2(n3594), .B1(n1089), .B2(mem[853]), .ZN(
        n3456) );
  NAND4_X1 U2981 ( .A1(n3459), .A2(n3458), .A3(n3457), .A4(n3456), .ZN(n3460)
         );
  NOR2_X1 U2982 ( .A1(n3461), .A2(n3460), .ZN(n3462) );
  NAND2_X1 U2983 ( .A1(n3463), .A2(n3462), .ZN(rdata_a_o[21]) );
  AOI22_X1 U2984 ( .A1(mem[598]), .A2(n1015), .B1(n995), .B2(mem[470]), .ZN(
        n3467) );
  AOI22_X1 U2985 ( .A1(mem[342]), .A2(n1006), .B1(n1083), .B2(mem[278]), .ZN(
        n3466) );
  AOI22_X1 U2986 ( .A1(mem[726]), .A2(n1082), .B1(n1012), .B2(mem[438]), .ZN(
        n3465) );
  AOI22_X1 U2987 ( .A1(n1009), .A2(mem[246]), .B1(mem[150]), .B2(n1021), .ZN(
        n3464) );
  NAND4_X1 U2988 ( .A1(n3467), .A2(n3466), .A3(n3465), .A4(n3464), .ZN(n3473)
         );
  AOI22_X1 U2989 ( .A1(mem[374]), .A2(n1023), .B1(n3577), .B2(mem[310]), .ZN(
        n3471) );
  AOI22_X1 U2990 ( .A1(n1093), .A2(mem[502]), .B1(mem[54]), .B2(n4729), .ZN(
        n3470) );
  AOI22_X1 U2991 ( .A1(mem[86]), .A2(n3579), .B1(n3578), .B2(mem[22]), .ZN(
        n3469) );
  NAND2_X1 U2992 ( .A1(n1027), .A2(mem[790]), .ZN(n3468) );
  NAND4_X1 U2993 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n3472)
         );
  NOR2_X1 U2994 ( .A1(n3473), .A2(n3472), .ZN(n3485) );
  AOI22_X1 U2995 ( .A1(mem[694]), .A2(n1070), .B1(n3585), .B2(mem[406]), .ZN(
        n3477) );
  AOI22_X1 U2996 ( .A1(n1017), .A2(mem[214]), .B1(mem[118]), .B2(n4736), .ZN(
        n3476) );
  AOI22_X1 U2997 ( .A1(mem[630]), .A2(n1071), .B1(n3586), .B2(mem[566]), .ZN(
        n3475) );
  AOI22_X1 U2998 ( .A1(n3587), .A2(mem[662]), .B1(mem[182]), .B2(n3517), .ZN(
        n3474) );
  NAND4_X1 U2999 ( .A1(n3477), .A2(n3476), .A3(n3475), .A4(n3474), .ZN(n3483)
         );
  AOI22_X1 U3000 ( .A1(n1068), .A2(mem[534]), .B1(mem[950]), .B2(n3592), .ZN(
        n3481) );
  AOI22_X1 U3001 ( .A1(mem[982]), .A2(n1073), .B1(n1086), .B2(mem[758]), .ZN(
        n3480) );
  AOI22_X1 U3002 ( .A1(mem[886]), .A2(n3593), .B1(n1069), .B2(mem[822]), .ZN(
        n3479) );
  AOI22_X1 U3003 ( .A1(mem[918]), .A2(n3455), .B1(n1091), .B2(mem[854]), .ZN(
        n3478) );
  NAND4_X1 U3004 ( .A1(n3481), .A2(n3480), .A3(n3479), .A4(n3478), .ZN(n3482)
         );
  NOR2_X1 U3005 ( .A1(n3483), .A2(n3482), .ZN(n3484) );
  NAND2_X1 U3006 ( .A1(n3485), .A2(n3484), .ZN(rdata_a_o[22]) );
  AOI22_X1 U3007 ( .A1(mem[599]), .A2(n1015), .B1(n996), .B2(mem[471]), .ZN(
        n3489) );
  AOI22_X1 U3008 ( .A1(mem[343]), .A2(n1006), .B1(n1083), .B2(mem[279]), .ZN(
        n3488) );
  AOI22_X1 U3009 ( .A1(mem[727]), .A2(n1082), .B1(n1012), .B2(mem[439]), .ZN(
        n3487) );
  AOI22_X1 U3010 ( .A1(n1010), .A2(mem[247]), .B1(mem[151]), .B2(n1022), .ZN(
        n3486) );
  NAND4_X1 U3011 ( .A1(n3489), .A2(n3488), .A3(n3487), .A4(n3486), .ZN(n3495)
         );
  AOI22_X1 U3012 ( .A1(mem[375]), .A2(n2161), .B1(n3577), .B2(mem[311]), .ZN(
        n3493) );
  AOI22_X1 U3013 ( .A1(n1092), .A2(mem[503]), .B1(mem[55]), .B2(n4730), .ZN(
        n3492) );
  AOI22_X1 U3014 ( .A1(mem[87]), .A2(n3579), .B1(n3578), .B2(mem[23]), .ZN(
        n3491) );
  NAND2_X1 U3015 ( .A1(n1027), .A2(mem[791]), .ZN(n3490) );
  NAND4_X1 U3016 ( .A1(n3493), .A2(n3492), .A3(n3491), .A4(n3490), .ZN(n3494)
         );
  NOR2_X1 U3017 ( .A1(n3495), .A2(n3494), .ZN(n3507) );
  AOI22_X1 U3018 ( .A1(mem[695]), .A2(n1070), .B1(n3585), .B2(mem[407]), .ZN(
        n3499) );
  AOI22_X1 U3019 ( .A1(n1017), .A2(mem[215]), .B1(mem[119]), .B2(n4736), .ZN(
        n3498) );
  AOI22_X1 U3020 ( .A1(mem[631]), .A2(n1071), .B1(n3586), .B2(mem[567]), .ZN(
        n3497) );
  AOI22_X1 U3021 ( .A1(n3587), .A2(mem[663]), .B1(mem[183]), .B2(n3517), .ZN(
        n3496) );
  NAND4_X1 U3022 ( .A1(n3499), .A2(n3498), .A3(n3497), .A4(n3496), .ZN(n3505)
         );
  AOI22_X1 U3023 ( .A1(n1068), .A2(mem[535]), .B1(mem[951]), .B2(n3592), .ZN(
        n3503) );
  AOI22_X1 U3024 ( .A1(mem[983]), .A2(n3564), .B1(n1087), .B2(mem[759]), .ZN(
        n3502) );
  AOI22_X1 U3025 ( .A1(mem[887]), .A2(n3593), .B1(n1069), .B2(mem[823]), .ZN(
        n3501) );
  AOI22_X1 U3026 ( .A1(mem[919]), .A2(n3455), .B1(n1090), .B2(mem[855]), .ZN(
        n3500) );
  NAND4_X1 U3027 ( .A1(n3503), .A2(n3502), .A3(n3501), .A4(n3500), .ZN(n3504)
         );
  NOR2_X1 U3028 ( .A1(n3505), .A2(n3504), .ZN(n3506) );
  NAND2_X1 U3029 ( .A1(n3507), .A2(n3506), .ZN(rdata_a_o[23]) );
  AOI22_X1 U3030 ( .A1(mem[600]), .A2(n1014), .B1(n996), .B2(mem[472]), .ZN(
        n3511) );
  AOI22_X1 U3031 ( .A1(mem[344]), .A2(n1005), .B1(n1085), .B2(mem[280]), .ZN(
        n3510) );
  AOI22_X1 U3032 ( .A1(mem[728]), .A2(n1081), .B1(n1011), .B2(mem[440]), .ZN(
        n3509) );
  AOI22_X1 U3033 ( .A1(n1008), .A2(mem[248]), .B1(mem[152]), .B2(n1020), .ZN(
        n3508) );
  AND4_X1 U3034 ( .A1(n3511), .A2(n3510), .A3(n3509), .A4(n3508), .ZN(n3529)
         );
  AOI22_X1 U3035 ( .A1(mem[376]), .A2(n1023), .B1(n3577), .B2(mem[312]), .ZN(
        n3516) );
  AOI22_X1 U3036 ( .A1(mem[88]), .A2(n3512), .B1(n3578), .B2(mem[24]), .ZN(
        n3515) );
  AOI22_X1 U3037 ( .A1(n1067), .A2(mem[504]), .B1(mem[56]), .B2(n4729), .ZN(
        n3514) );
  NAND2_X1 U3038 ( .A1(n1025), .A2(mem[792]), .ZN(n3513) );
  AND4_X1 U3039 ( .A1(n3516), .A2(n3515), .A3(n3514), .A4(n3513), .ZN(n3528)
         );
  AOI22_X1 U3040 ( .A1(mem[696]), .A2(n1070), .B1(n3585), .B2(mem[408]), .ZN(
        n3521) );
  AOI22_X1 U3041 ( .A1(n1019), .A2(mem[216]), .B1(mem[120]), .B2(n4736), .ZN(
        n3520) );
  AOI22_X1 U3042 ( .A1(mem[632]), .A2(n1071), .B1(n3586), .B2(mem[568]), .ZN(
        n3519) );
  AOI22_X1 U3043 ( .A1(n3587), .A2(mem[664]), .B1(mem[184]), .B2(n3517), .ZN(
        n3518) );
  AND4_X1 U3044 ( .A1(n3521), .A2(n3520), .A3(n3519), .A4(n3518), .ZN(n3527)
         );
  AOI22_X1 U3045 ( .A1(n1068), .A2(mem[536]), .B1(mem[952]), .B2(n3592), .ZN(
        n3525) );
  AOI22_X1 U3046 ( .A1(mem[984]), .A2(n1073), .B1(n1088), .B2(mem[760]), .ZN(
        n3524) );
  AOI22_X1 U3047 ( .A1(mem[888]), .A2(n3593), .B1(n1069), .B2(mem[824]), .ZN(
        n3523) );
  AOI22_X1 U3048 ( .A1(mem[920]), .A2(n3455), .B1(n1089), .B2(mem[856]), .ZN(
        n3522) );
  AND4_X1 U3049 ( .A1(n3525), .A2(n3524), .A3(n3523), .A4(n3522), .ZN(n3526)
         );
  NAND4_X1 U3050 ( .A1(n3529), .A2(n3528), .A3(n3527), .A4(n3526), .ZN(
        rdata_a_o[24]) );
  AOI22_X1 U3051 ( .A1(mem[345]), .A2(n1005), .B1(n1083), .B2(mem[281]), .ZN(
        n3531) );
  AOI22_X1 U3052 ( .A1(mem[729]), .A2(n1080), .B1(n1011), .B2(mem[441]), .ZN(
        n3530) );
  AND2_X1 U3053 ( .A1(n3531), .A2(n3530), .ZN(n3551) );
  AOI22_X1 U3054 ( .A1(mem[601]), .A2(n1016), .B1(n996), .B2(mem[473]), .ZN(
        n3533) );
  AOI22_X1 U3055 ( .A1(n1010), .A2(mem[249]), .B1(mem[153]), .B2(n1022), .ZN(
        n3532) );
  AND2_X1 U3056 ( .A1(n3533), .A2(n3532), .ZN(n3550) );
  AOI22_X1 U3057 ( .A1(mem[697]), .A2(n1070), .B1(n3585), .B2(mem[409]), .ZN(
        n3537) );
  AOI22_X1 U3058 ( .A1(n1019), .A2(mem[217]), .B1(mem[121]), .B2(n4736), .ZN(
        n3536) );
  AOI22_X1 U3059 ( .A1(mem[633]), .A2(n1071), .B1(n3586), .B2(mem[569]), .ZN(
        n3535) );
  AOI22_X1 U3060 ( .A1(n3587), .A2(mem[665]), .B1(mem[185]), .B2(n1072), .ZN(
        n3534) );
  NAND4_X1 U3061 ( .A1(n3537), .A2(n3536), .A3(n3535), .A4(n3534), .ZN(n3543)
         );
  AOI22_X1 U3062 ( .A1(n1068), .A2(mem[537]), .B1(mem[953]), .B2(n3592), .ZN(
        n3541) );
  AOI22_X1 U3063 ( .A1(mem[985]), .A2(n3564), .B1(n1087), .B2(mem[761]), .ZN(
        n3540) );
  AOI22_X1 U3064 ( .A1(mem[889]), .A2(n3593), .B1(n1069), .B2(mem[825]), .ZN(
        n3539) );
  AOI22_X1 U3065 ( .A1(mem[921]), .A2(n3269), .B1(n1091), .B2(mem[857]), .ZN(
        n3538) );
  NAND4_X1 U3066 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), .ZN(n3542)
         );
  NOR2_X1 U3067 ( .A1(n3543), .A2(n3542), .ZN(n3549) );
  AOI22_X1 U3068 ( .A1(mem[377]), .A2(n1023), .B1(n3577), .B2(mem[313]), .ZN(
        n3547) );
  AOI22_X1 U3069 ( .A1(mem[89]), .A2(n3579), .B1(n3578), .B2(mem[25]), .ZN(
        n3546) );
  AOI22_X1 U3070 ( .A1(n1067), .A2(mem[505]), .B1(mem[57]), .B2(n4730), .ZN(
        n3545) );
  NAND2_X1 U3071 ( .A1(n1026), .A2(mem[793]), .ZN(n3544) );
  AND4_X1 U3072 ( .A1(n3547), .A2(n3546), .A3(n3545), .A4(n3544), .ZN(n3548)
         );
  NAND4_X1 U3073 ( .A1(n3551), .A2(n3550), .A3(n3549), .A4(n3548), .ZN(
        rdata_a_o[25]) );
  AOI22_X1 U3074 ( .A1(mem[602]), .A2(n1014), .B1(n995), .B2(mem[474]), .ZN(
        n3555) );
  AOI22_X1 U3075 ( .A1(mem[346]), .A2(n1005), .B1(n1085), .B2(mem[282]), .ZN(
        n3554) );
  AOI22_X1 U3076 ( .A1(mem[730]), .A2(n1080), .B1(n1013), .B2(mem[442]), .ZN(
        n3553) );
  AOI22_X1 U3077 ( .A1(n1008), .A2(mem[250]), .B1(mem[154]), .B2(n1020), .ZN(
        n3552) );
  AND4_X1 U3078 ( .A1(n3555), .A2(n3554), .A3(n3553), .A4(n3552), .ZN(n3572)
         );
  AOI22_X1 U3079 ( .A1(mem[378]), .A2(n1023), .B1(n3577), .B2(mem[314]), .ZN(
        n3559) );
  AOI22_X1 U3080 ( .A1(mem[90]), .A2(n3579), .B1(n3578), .B2(mem[26]), .ZN(
        n3558) );
  AOI22_X1 U3081 ( .A1(n1067), .A2(mem[506]), .B1(mem[58]), .B2(n4730), .ZN(
        n3557) );
  NAND2_X1 U3082 ( .A1(n1025), .A2(mem[794]), .ZN(n3556) );
  AND4_X1 U3083 ( .A1(n3559), .A2(n3558), .A3(n3557), .A4(n3556), .ZN(n3571)
         );
  AOI22_X1 U3084 ( .A1(mem[698]), .A2(n1070), .B1(n3585), .B2(mem[410]), .ZN(
        n3563) );
  AOI22_X1 U3085 ( .A1(n1019), .A2(mem[218]), .B1(mem[122]), .B2(n1029), .ZN(
        n3562) );
  AOI22_X1 U3086 ( .A1(mem[634]), .A2(n1071), .B1(n3586), .B2(mem[570]), .ZN(
        n3561) );
  AOI22_X1 U3087 ( .A1(n3587), .A2(mem[666]), .B1(mem[186]), .B2(n1072), .ZN(
        n3560) );
  AND4_X1 U3088 ( .A1(n3563), .A2(n3562), .A3(n3561), .A4(n3560), .ZN(n3570)
         );
  AOI22_X1 U3089 ( .A1(n1068), .A2(mem[538]), .B1(mem[954]), .B2(n3592), .ZN(
        n3568) );
  AOI22_X1 U3090 ( .A1(mem[986]), .A2(n3564), .B1(n1088), .B2(mem[762]), .ZN(
        n3567) );
  AOI22_X1 U3091 ( .A1(mem[890]), .A2(n3593), .B1(n1069), .B2(mem[826]), .ZN(
        n3566) );
  AOI22_X1 U3092 ( .A1(mem[922]), .A2(n3594), .B1(n1089), .B2(mem[858]), .ZN(
        n3565) );
  AND4_X1 U3093 ( .A1(n3568), .A2(n3567), .A3(n3566), .A4(n3565), .ZN(n3569)
         );
  NAND4_X1 U3094 ( .A1(n3572), .A2(n3571), .A3(n3570), .A4(n3569), .ZN(
        rdata_a_o[26]) );
  AOI22_X1 U3095 ( .A1(mem[603]), .A2(n1015), .B1(n995), .B2(mem[475]), .ZN(
        n3576) );
  AOI22_X1 U3096 ( .A1(mem[347]), .A2(n1006), .B1(n1084), .B2(mem[283]), .ZN(
        n3575) );
  AOI22_X1 U3097 ( .A1(mem[731]), .A2(n1081), .B1(n1012), .B2(mem[443]), .ZN(
        n3574) );
  AOI22_X1 U3098 ( .A1(n1009), .A2(mem[251]), .B1(mem[155]), .B2(n1021), .ZN(
        n3573) );
  AND4_X1 U3099 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3602)
         );
  AOI22_X1 U3100 ( .A1(mem[379]), .A2(n1024), .B1(n3577), .B2(mem[315]), .ZN(
        n3584) );
  AOI22_X1 U3101 ( .A1(mem[91]), .A2(n3579), .B1(n3578), .B2(mem[27]), .ZN(
        n3583) );
  AOI22_X1 U3102 ( .A1(n1093), .A2(mem[507]), .B1(mem[59]), .B2(n4729), .ZN(
        n3582) );
  NAND2_X1 U3103 ( .A1(n1026), .A2(mem[795]), .ZN(n3581) );
  AND4_X1 U3104 ( .A1(n3584), .A2(n3583), .A3(n3582), .A4(n3581), .ZN(n3601)
         );
  AOI22_X1 U3105 ( .A1(mem[699]), .A2(n1070), .B1(n3585), .B2(mem[411]), .ZN(
        n3591) );
  AOI22_X1 U3106 ( .A1(n1019), .A2(mem[219]), .B1(mem[123]), .B2(n1029), .ZN(
        n3590) );
  AOI22_X1 U3107 ( .A1(mem[635]), .A2(n1071), .B1(n3586), .B2(mem[571]), .ZN(
        n3589) );
  AOI22_X1 U3108 ( .A1(n3587), .A2(mem[667]), .B1(mem[187]), .B2(n1072), .ZN(
        n3588) );
  AND4_X1 U3109 ( .A1(n3591), .A2(n3590), .A3(n3589), .A4(n3588), .ZN(n3600)
         );
  AOI22_X1 U3110 ( .A1(n1068), .A2(mem[539]), .B1(mem[955]), .B2(n3592), .ZN(
        n3598) );
  AOI22_X1 U3111 ( .A1(mem[987]), .A2(n1073), .B1(n1088), .B2(mem[763]), .ZN(
        n3597) );
  AOI22_X1 U3112 ( .A1(mem[891]), .A2(n3593), .B1(n1069), .B2(mem[827]), .ZN(
        n3596) );
  AOI22_X1 U3113 ( .A1(mem[923]), .A2(n3269), .B1(n1089), .B2(mem[859]), .ZN(
        n3595) );
  AND4_X1 U3114 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3599)
         );
  NAND4_X1 U3115 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(
        rdata_a_o[27]) );
  BUF_X1 U3125 ( .A(wdata_a_i[7]), .Z(n4486) );
  INV_X1 U3141 ( .A(wdata_b_i[14]), .ZN(n4436) );
  INV_X1 U3144 ( .A(wdata_b_i[15]), .ZN(n4439) );
  INV_X1 U3147 ( .A(wdata_b_i[16]), .ZN(n4441) );
  INV_X1 U3150 ( .A(wdata_b_i[17]), .ZN(n4037) );
  INV_X1 U3156 ( .A(wdata_b_i[19]), .ZN(n4040) );
  INV_X1 U3159 ( .A(wdata_b_i[20]), .ZN(n4447) );
  INV_X1 U3162 ( .A(wdata_b_i[22]), .ZN(n4043) );
  INV_X1 U3174 ( .A(wdata_b_i[26]), .ZN(n4458) );
  INV_X1 U3177 ( .A(wdata_b_i[27]), .ZN(n4461) );
  INV_X1 U3185 ( .A(wdata_b_i[30]), .ZN(n4470) );
  NOR2_X1 U3415 ( .A1(n3769), .A2(n3768), .ZN(n3846) );
  NAND2_X1 U3417 ( .A1(n3771), .A2(n3847), .ZN(n3772) );
  NAND2_X1 U3542 ( .A1(n3848), .A2(n3847), .ZN(n3849) );
  SDFFR_X1 mem_reg_1__31_ ( .D(n8404), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[31]) );
  SDFFR_X1 mem_reg_1__30_ ( .D(n8405), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[30]) );
  SDFFR_X1 mem_reg_1__29_ ( .D(n8406), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[29]) );
  SDFFR_X1 mem_reg_1__26_ ( .D(n8409), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[26]) );
  SDFFR_X1 mem_reg_1__23_ ( .D(n8412), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[23]) );
  SDFFR_X1 mem_reg_1__18_ ( .D(n8417), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[18]) );
  SDFFR_X1 mem_reg_1__16_ ( .D(n8419), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[16]) );
  SDFFR_X1 mem_reg_1__14_ ( .D(n8421), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[14]) );
  SDFFR_X1 mem_reg_1__13_ ( .D(n8422), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[13]) );
  SDFFR_X1 mem_reg_1__12_ ( .D(n8423), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[12]) );
  SDFFR_X1 mem_reg_1__11_ ( .D(n8424), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[11]) );
  SDFFR_X1 mem_reg_1__10_ ( .D(n8425), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[10]) );
  SDFFR_X1 mem_reg_1__9_ ( .D(n8426), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[9]) );
  SDFFR_X1 mem_reg_1__8_ ( .D(n8427), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[8]) );
  SDFFR_X1 mem_reg_1__7_ ( .D(n8428), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[7]) );
  SDFFR_X1 mem_reg_1__6_ ( .D(n8429), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[6]) );
  SDFFR_X1 mem_reg_1__5_ ( .D(n8430), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[5]) );
  SDFFR_X1 mem_reg_1__4_ ( .D(n8431), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[4]) );
  SDFFR_X1 mem_reg_1__3_ ( .D(n8432), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[3]) );
  SDFFR_X1 mem_reg_1__2_ ( .D(n8433), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[2]) );
  SDFFR_X1 mem_reg_1__1_ ( .D(n8434), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[1]) );
  SDFFR_X1 mem_reg_2__31_ ( .D(n8788), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[63]) );
  SDFFR_X1 mem_reg_2__30_ ( .D(n8789), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[62]) );
  SDFFR_X1 mem_reg_2__29_ ( .D(n8790), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[61]) );
  SDFFR_X1 mem_reg_2__26_ ( .D(n8793), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[58]) );
  SDFFR_X1 mem_reg_2__23_ ( .D(n8796), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[55]) );
  SDFFR_X1 mem_reg_2__18_ ( .D(n8801), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[50]) );
  SDFFR_X1 mem_reg_2__16_ ( .D(n8803), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[48]) );
  SDFFR_X1 mem_reg_2__15_ ( .D(n8804), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[47]) );
  SDFFR_X1 mem_reg_2__14_ ( .D(n8805), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[46]) );
  SDFFR_X1 mem_reg_2__13_ ( .D(n8806), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[45]) );
  SDFFR_X1 mem_reg_2__12_ ( .D(n8807), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[44]) );
  SDFFR_X1 mem_reg_2__11_ ( .D(n8808), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[43]) );
  SDFFR_X1 mem_reg_2__10_ ( .D(n8809), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[42]) );
  SDFFR_X1 mem_reg_2__9_ ( .D(n8810), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[41]) );
  SDFFR_X1 mem_reg_2__8_ ( .D(n8811), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[40]) );
  SDFFR_X1 mem_reg_2__7_ ( .D(n8812), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[39]) );
  SDFFR_X1 mem_reg_2__6_ ( .D(n8813), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[38]) );
  SDFFR_X1 mem_reg_2__4_ ( .D(n8815), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[36]) );
  SDFFR_X1 mem_reg_2__3_ ( .D(n8816), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[35]) );
  SDFFR_X1 mem_reg_2__2_ ( .D(n8817), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[34]) );
  SDFFR_X1 mem_reg_2__1_ ( .D(n8818), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[33]) );
  SDFFR_X1 mem_reg_3__31_ ( .D(n8915), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[95]) );
  SDFFR_X1 mem_reg_3__30_ ( .D(n8916), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[94]) );
  SDFFR_X1 mem_reg_3__29_ ( .D(n8917), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[93]) );
  SDFFR_X1 mem_reg_3__26_ ( .D(n8920), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[90]) );
  SDFFR_X1 mem_reg_3__24_ ( .D(n8922), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[88]) );
  SDFFR_X1 mem_reg_3__23_ ( .D(n8924), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[87]) );
  SDFFR_X1 mem_reg_3__18_ ( .D(n8929), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[82]) );
  SDFFR_X1 mem_reg_3__16_ ( .D(n8931), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[80]) );
  SDFFR_X1 mem_reg_3__14_ ( .D(n8933), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[78]) );
  SDFFR_X1 mem_reg_3__13_ ( .D(n8934), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[77]) );
  SDFFR_X1 mem_reg_3__12_ ( .D(n8935), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[76]) );
  SDFFR_X1 mem_reg_3__11_ ( .D(n8936), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[75]) );
  SDFFR_X1 mem_reg_3__10_ ( .D(n8937), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[74]) );
  SDFFR_X1 mem_reg_3__9_ ( .D(n8938), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[73]) );
  SDFFR_X1 mem_reg_3__8_ ( .D(n8939), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[72]) );
  SDFFR_X1 mem_reg_3__7_ ( .D(n8940), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[71]) );
  SDFFR_X1 mem_reg_3__6_ ( .D(n8941), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[70]) );
  SDFFR_X1 mem_reg_3__5_ ( .D(n8942), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[69]) );
  SDFFR_X1 mem_reg_3__4_ ( .D(n8943), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[68]) );
  SDFFR_X1 mem_reg_3__3_ ( .D(n8944), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[67]) );
  SDFFR_X1 mem_reg_3__2_ ( .D(n8945), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[66]) );
  SDFFR_X1 mem_reg_3__1_ ( .D(n8946), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[65]) );
  SDFFR_X1 mem_reg_4__31_ ( .D(n8951), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[127]) );
  SDFFR_X1 mem_reg_4__30_ ( .D(n8952), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[126]) );
  SDFFR_X1 mem_reg_4__29_ ( .D(n8953), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[125]) );
  SDFFR_X1 mem_reg_4__28_ ( .D(n8954), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[124]) );
  SDFFR_X1 mem_reg_4__27_ ( .D(n8955), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[123]) );
  SDFFR_X1 mem_reg_4__26_ ( .D(n8956), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[122]) );
  SDFFR_X1 mem_reg_4__25_ ( .D(n8957), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[121]) );
  SDFFR_X1 mem_reg_4__24_ ( .D(n8958), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[120]) );
  SDFFR_X1 mem_reg_4__23_ ( .D(n8959), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[119]) );
  SDFFR_X1 mem_reg_4__18_ ( .D(n8964), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[114]) );
  SDFFR_X1 mem_reg_4__16_ ( .D(n8966), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[112]) );
  SDFFR_X1 mem_reg_4__15_ ( .D(n8967), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[111]) );
  SDFFR_X1 mem_reg_4__14_ ( .D(n8968), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[110]) );
  SDFFR_X1 mem_reg_4__13_ ( .D(n8969), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[109]) );
  SDFFR_X1 mem_reg_4__12_ ( .D(n8970), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[108]) );
  SDFFR_X1 mem_reg_4__11_ ( .D(n8971), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[107]) );
  SDFFR_X1 mem_reg_4__10_ ( .D(n8972), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[106]) );
  SDFFR_X1 mem_reg_4__9_ ( .D(n8973), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[105]) );
  SDFFR_X1 mem_reg_4__8_ ( .D(n8974), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[104]) );
  SDFFR_X1 mem_reg_4__7_ ( .D(n8975), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[103]) );
  SDFFR_X1 mem_reg_4__6_ ( .D(n8976), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[102]) );
  SDFFR_X1 mem_reg_4__4_ ( .D(n8978), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[100]) );
  SDFFR_X1 mem_reg_4__3_ ( .D(n8979), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[99]) );
  SDFFR_X1 mem_reg_4__2_ ( .D(n8980), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[98]) );
  SDFFR_X1 mem_reg_4__1_ ( .D(n8981), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[97]) );
  SDFFR_X1 mem_reg_5__31_ ( .D(n8986), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[159]) );
  SDFFR_X1 mem_reg_5__30_ ( .D(n8987), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[158]) );
  SDFFR_X1 mem_reg_5__29_ ( .D(n8988), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[157]) );
  SDFFR_X1 mem_reg_5__26_ ( .D(n8991), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[154]) );
  SDFFR_X1 mem_reg_5__24_ ( .D(n8993), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[152]) );
  SDFFR_X1 mem_reg_5__18_ ( .D(n8999), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[146]) );
  SDFFR_X1 mem_reg_5__16_ ( .D(n9001), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[144]) );
  SDFFR_X1 mem_reg_5__15_ ( .D(n9002), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[143]) );
  SDFFR_X1 mem_reg_5__14_ ( .D(n9003), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[142]) );
  SDFFR_X1 mem_reg_5__13_ ( .D(n9004), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[141]) );
  SDFFR_X1 mem_reg_5__12_ ( .D(n9005), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[140]) );
  SDFFR_X1 mem_reg_5__11_ ( .D(n9006), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[139]) );
  SDFFR_X1 mem_reg_5__10_ ( .D(n9007), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[138]) );
  SDFFR_X1 mem_reg_5__9_ ( .D(n9008), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[137]) );
  SDFFR_X1 mem_reg_5__8_ ( .D(n9009), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[136]) );
  SDFFR_X1 mem_reg_5__7_ ( .D(n9010), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[135]) );
  SDFFR_X1 mem_reg_5__6_ ( .D(n9011), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[134]) );
  SDFFR_X1 mem_reg_5__5_ ( .D(n9012), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[133]) );
  SDFFR_X1 mem_reg_5__4_ ( .D(n9013), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[132]) );
  SDFFR_X1 mem_reg_5__3_ ( .D(n9014), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[131]) );
  SDFFR_X1 mem_reg_5__2_ ( .D(n9015), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[130]) );
  SDFFR_X1 mem_reg_5__1_ ( .D(n9016), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[129]) );
  SDFFR_X1 mem_reg_6__31_ ( .D(n9021), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[191]) );
  SDFFR_X1 mem_reg_6__30_ ( .D(n9022), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[190]) );
  SDFFR_X1 mem_reg_6__29_ ( .D(n9023), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[189]) );
  SDFFR_X1 mem_reg_6__28_ ( .D(n9024), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[188]) );
  SDFFR_X1 mem_reg_6__27_ ( .D(n9025), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[187]) );
  SDFFR_X1 mem_reg_6__26_ ( .D(n9026), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[186]) );
  SDFFR_X1 mem_reg_6__25_ ( .D(n9027), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[185]) );
  SDFFR_X1 mem_reg_6__24_ ( .D(n9028), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[184]) );
  SDFFR_X1 mem_reg_6__23_ ( .D(n9029), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[183]) );
  SDFFR_X1 mem_reg_6__21_ ( .D(n9031), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[181]) );
  SDFFR_X1 mem_reg_6__18_ ( .D(n9035), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[178]) );
  SDFFR_X1 mem_reg_6__16_ ( .D(n9037), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[176]) );
  SDFFR_X1 mem_reg_6__15_ ( .D(n9038), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[175]) );
  SDFFR_X1 mem_reg_6__14_ ( .D(n9039), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[174]) );
  SDFFR_X1 mem_reg_6__13_ ( .D(n9040), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[173]) );
  SDFFR_X1 mem_reg_6__12_ ( .D(n9041), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[172]) );
  SDFFR_X1 mem_reg_6__11_ ( .D(n9042), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[171]) );
  SDFFR_X1 mem_reg_6__10_ ( .D(n9043), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[170]) );
  SDFFR_X1 mem_reg_6__9_ ( .D(n9044), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[169]) );
  SDFFR_X1 mem_reg_6__8_ ( .D(n9045), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[168]) );
  SDFFR_X1 mem_reg_6__7_ ( .D(n9046), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[167]) );
  SDFFR_X1 mem_reg_6__6_ ( .D(n9047), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[166]) );
  SDFFR_X1 mem_reg_6__5_ ( .D(n9048), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[165]) );
  SDFFR_X1 mem_reg_6__4_ ( .D(n9049), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[164]) );
  SDFFR_X1 mem_reg_6__3_ ( .D(n9050), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[163]) );
  SDFFR_X1 mem_reg_6__2_ ( .D(n9051), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[162]) );
  SDFFR_X1 mem_reg_6__1_ ( .D(n9052), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[161]) );
  SDFFR_X1 mem_reg_7__31_ ( .D(n9057), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[223]) );
  SDFFR_X1 mem_reg_7__30_ ( .D(n9058), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[222]) );
  SDFFR_X1 mem_reg_7__29_ ( .D(n9059), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[221]) );
  SDFFR_X1 mem_reg_7__27_ ( .D(n9061), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[219]) );
  SDFFR_X1 mem_reg_7__26_ ( .D(n9062), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[218]) );
  SDFFR_X1 mem_reg_7__24_ ( .D(n9065), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[216]) );
  SDFFR_X1 mem_reg_7__23_ ( .D(n9066), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[215]) );
  SDFFR_X1 mem_reg_7__22_ ( .D(n9067), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[214]) );
  SDFFR_X1 mem_reg_7__21_ ( .D(n9069), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[213]) );
  SDFFR_X1 mem_reg_7__20_ ( .D(n9071), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[212]) );
  SDFFR_X1 mem_reg_7__19_ ( .D(n9073), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[211]) );
  SDFFR_X1 mem_reg_7__18_ ( .D(n9075), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[210]) );
  SDFFR_X1 mem_reg_7__17_ ( .D(n9077), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[209]) );
  SDFFR_X1 mem_reg_7__16_ ( .D(n9079), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[208]) );
  SDFFR_X1 mem_reg_7__15_ ( .D(n9080), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[207]) );
  SDFFR_X1 mem_reg_7__14_ ( .D(n9082), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[206]) );
  SDFFR_X1 mem_reg_7__13_ ( .D(n9083), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[205]) );
  SDFFR_X1 mem_reg_7__12_ ( .D(n9084), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[204]) );
  SDFFR_X1 mem_reg_7__11_ ( .D(n9086), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[203]) );
  SDFFR_X1 mem_reg_7__10_ ( .D(n9088), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[202]) );
  SDFFR_X1 mem_reg_7__9_ ( .D(n9090), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[201]) );
  SDFFR_X1 mem_reg_7__8_ ( .D(n9092), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[200]) );
  SDFFR_X1 mem_reg_7__7_ ( .D(n9093), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[199]) );
  SDFFR_X1 mem_reg_7__6_ ( .D(n9094), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[198]) );
  SDFFR_X1 mem_reg_7__5_ ( .D(n9095), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[197]) );
  SDFFR_X1 mem_reg_7__4_ ( .D(n9097), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[196]) );
  SDFFR_X1 mem_reg_7__3_ ( .D(n9099), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[195]) );
  SDFFR_X1 mem_reg_7__2_ ( .D(n9101), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[194]) );
  SDFFR_X1 mem_reg_7__1_ ( .D(n9103), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[193]) );
  SDFFR_X1 mem_reg_7__0_ ( .D(n9105), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[192]) );
  SDFFR_X1 mem_reg_8__29_ ( .D(n9111), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[253]) );
  SDFFR_X1 mem_reg_8__28_ ( .D(n9112), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[252]) );
  SDFFR_X1 mem_reg_8__27_ ( .D(n9113), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[251]) );
  SDFFR_X1 mem_reg_8__26_ ( .D(n9114), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[250]) );
  SDFFR_X1 mem_reg_8__25_ ( .D(n9115), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[249]) );
  SDFFR_X1 mem_reg_8__24_ ( .D(n9116), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[248]) );
  SDFFR_X1 mem_reg_8__16_ ( .D(n9124), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[240]) );
  SDFFR_X1 mem_reg_8__14_ ( .D(n9126), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[238]) );
  SDFFR_X1 mem_reg_8__13_ ( .D(n9127), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[237]) );
  SDFFR_X1 mem_reg_8__12_ ( .D(n9128), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[236]) );
  SDFFR_X1 mem_reg_8__11_ ( .D(n9129), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[235]) );
  SDFFR_X1 mem_reg_8__9_ ( .D(n9131), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[233]) );
  SDFFR_X1 mem_reg_8__8_ ( .D(n9132), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[232]) );
  SDFFR_X1 mem_reg_8__6_ ( .D(n9134), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[230]) );
  SDFFR_X1 mem_reg_8__4_ ( .D(n9136), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[228]) );
  SDFFR_X1 mem_reg_8__3_ ( .D(n9137), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[227]) );
  SDFFR_X1 mem_reg_8__2_ ( .D(n9138), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[226]) );
  SDFFR_X1 mem_reg_8__1_ ( .D(n9139), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[225]) );
  SDFFR_X1 mem_reg_9__31_ ( .D(n9144), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[287]) );
  SDFFR_X1 mem_reg_9__30_ ( .D(n9145), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[286]) );
  SDFFR_X1 mem_reg_9__29_ ( .D(n9147), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[285]) );
  SDFFR_X1 mem_reg_9__28_ ( .D(n9148), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[284]) );
  SDFFR_X1 mem_reg_9__27_ ( .D(n9149), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[283]) );
  SDFFR_X1 mem_reg_9__26_ ( .D(n9151), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[282]) );
  SDFFR_X1 mem_reg_9__25_ ( .D(n9153), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[281]) );
  SDFFR_X1 mem_reg_9__24_ ( .D(n9154), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[280]) );
  SDFFR_X1 mem_reg_9__23_ ( .D(n9156), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[279]) );
  SDFFR_X1 mem_reg_9__22_ ( .D(n9158), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[278]) );
  SDFFR_X1 mem_reg_9__21_ ( .D(n9160), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[277]) );
  SDFFR_X1 mem_reg_9__20_ ( .D(n9161), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[276]) );
  SDFFR_X1 mem_reg_9__19_ ( .D(n9163), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[275]) );
  SDFFR_X1 mem_reg_9__18_ ( .D(n9165), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[274]) );
  SDFFR_X1 mem_reg_9__17_ ( .D(n9167), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[273]) );
  SDFFR_X1 mem_reg_9__16_ ( .D(n9169), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[272]) );
  SDFFR_X1 mem_reg_9__15_ ( .D(n9170), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[271]) );
  SDFFR_X1 mem_reg_9__14_ ( .D(n9171), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[270]) );
  SDFFR_X1 mem_reg_9__13_ ( .D(n9173), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[269]) );
  SDFFR_X1 mem_reg_9__12_ ( .D(n9175), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[268]) );
  SDFFR_X1 mem_reg_9__11_ ( .D(n9176), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[267]) );
  SDFFR_X1 mem_reg_9__10_ ( .D(n9177), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[266]) );
  SDFFR_X1 mem_reg_9__9_ ( .D(n9179), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[265]) );
  SDFFR_X1 mem_reg_9__8_ ( .D(n9180), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[264]) );
  SDFFR_X1 mem_reg_9__7_ ( .D(n9181), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[263]) );
  SDFFR_X1 mem_reg_9__6_ ( .D(n9183), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[262]) );
  SDFFR_X1 mem_reg_9__5_ ( .D(n9185), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[261]) );
  SDFFR_X1 mem_reg_9__4_ ( .D(n9187), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[260]) );
  SDFFR_X1 mem_reg_9__3_ ( .D(n9188), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[259]) );
  SDFFR_X1 mem_reg_9__2_ ( .D(n9190), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[258]) );
  SDFFR_X1 mem_reg_9__1_ ( .D(n9192), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[257]) );
  SDFFR_X1 mem_reg_9__0_ ( .D(n9194), .SI(1'b0), .SE(1'b0), .CK(n9196), .RN(
        rst_n), .Q(mem[256]) );
  SDFFR_X1 mem_reg_10__29_ ( .D(n8055), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[317]) );
  SDFFR_X1 mem_reg_10__28_ ( .D(n8056), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[316]) );
  SDFFR_X1 mem_reg_10__27_ ( .D(n8057), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[315]) );
  SDFFR_X1 mem_reg_10__26_ ( .D(n8058), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[314]) );
  SDFFR_X1 mem_reg_10__25_ ( .D(n8059), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[313]) );
  SDFFR_X1 mem_reg_10__24_ ( .D(n8060), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[312]) );
  SDFFR_X1 mem_reg_10__16_ ( .D(n8068), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[304]) );
  SDFFR_X1 mem_reg_10__14_ ( .D(n8070), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[302]) );
  SDFFR_X1 mem_reg_10__13_ ( .D(n8071), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[301]) );
  SDFFR_X1 mem_reg_10__12_ ( .D(n8072), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[300]) );
  SDFFR_X1 mem_reg_10__11_ ( .D(n8073), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[299]) );
  SDFFR_X1 mem_reg_10__9_ ( .D(n8075), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[297]) );
  SDFFR_X1 mem_reg_10__8_ ( .D(n8076), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[296]) );
  SDFFR_X1 mem_reg_10__6_ ( .D(n8078), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[294]) );
  SDFFR_X1 mem_reg_10__5_ ( .D(n8079), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[293]) );
  SDFFR_X1 mem_reg_10__4_ ( .D(n8080), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[292]) );
  SDFFR_X1 mem_reg_10__3_ ( .D(n8081), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[291]) );
  SDFFR_X1 mem_reg_10__2_ ( .D(n8082), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[290]) );
  SDFFR_X1 mem_reg_10__1_ ( .D(n8083), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[289]) );
  SDFFR_X1 mem_reg_11__29_ ( .D(n8090), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[349]) );
  SDFFR_X1 mem_reg_11__16_ ( .D(n8103), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[336]) );
  SDFFR_X1 mem_reg_11__14_ ( .D(n8105), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[334]) );
  SDFFR_X1 mem_reg_11__13_ ( .D(n8106), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[333]) );
  SDFFR_X1 mem_reg_11__12_ ( .D(n8107), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[332]) );
  SDFFR_X1 mem_reg_11__11_ ( .D(n8108), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[331]) );
  SDFFR_X1 mem_reg_11__10_ ( .D(n8109), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[330]) );
  SDFFR_X1 mem_reg_11__9_ ( .D(n8110), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[329]) );
  SDFFR_X1 mem_reg_11__8_ ( .D(n8111), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[328]) );
  SDFFR_X1 mem_reg_11__7_ ( .D(n8112), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[327]) );
  SDFFR_X1 mem_reg_11__6_ ( .D(n8113), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[326]) );
  SDFFR_X1 mem_reg_11__4_ ( .D(n8115), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[324]) );
  SDFFR_X1 mem_reg_11__3_ ( .D(n8116), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[323]) );
  SDFFR_X1 mem_reg_11__2_ ( .D(n8117), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[322]) );
  SDFFR_X1 mem_reg_11__1_ ( .D(n8118), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[321]) );
  SDFFR_X1 mem_reg_12__29_ ( .D(n8125), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[381]) );
  SDFFR_X1 mem_reg_12__28_ ( .D(n8126), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[380]) );
  SDFFR_X1 mem_reg_12__27_ ( .D(n8127), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[379]) );
  SDFFR_X1 mem_reg_12__26_ ( .D(n8128), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[378]) );
  SDFFR_X1 mem_reg_12__25_ ( .D(n8129), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[377]) );
  SDFFR_X1 mem_reg_12__24_ ( .D(n8130), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[376]) );
  SDFFR_X1 mem_reg_12__16_ ( .D(n8138), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[368]) );
  SDFFR_X1 mem_reg_12__14_ ( .D(n8140), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[366]) );
  SDFFR_X1 mem_reg_12__13_ ( .D(n8141), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[365]) );
  SDFFR_X1 mem_reg_12__12_ ( .D(n8142), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[364]) );
  SDFFR_X1 mem_reg_12__11_ ( .D(n8143), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[363]) );
  SDFFR_X1 mem_reg_12__9_ ( .D(n8145), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[361]) );
  SDFFR_X1 mem_reg_12__8_ ( .D(n8146), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[360]) );
  SDFFR_X1 mem_reg_12__7_ ( .D(n8147), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[359]) );
  SDFFR_X1 mem_reg_12__6_ ( .D(n8148), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[358]) );
  SDFFR_X1 mem_reg_12__5_ ( .D(n8149), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[357]) );
  SDFFR_X1 mem_reg_12__4_ ( .D(n8150), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[356]) );
  SDFFR_X1 mem_reg_12__3_ ( .D(n8151), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[355]) );
  SDFFR_X1 mem_reg_12__2_ ( .D(n8152), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[354]) );
  SDFFR_X1 mem_reg_12__1_ ( .D(n8153), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[353]) );
  SDFFR_X1 mem_reg_12__0_ ( .D(n8154), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[352]) );
  SDFFR_X1 mem_reg_13__31_ ( .D(n8158), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[415]) );
  SDFFR_X1 mem_reg_13__16_ ( .D(n8173), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[400]) );
  SDFFR_X1 mem_reg_13__14_ ( .D(n8175), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[398]) );
  SDFFR_X1 mem_reg_13__13_ ( .D(n8176), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[397]) );
  SDFFR_X1 mem_reg_13__12_ ( .D(n8177), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[396]) );
  SDFFR_X1 mem_reg_13__11_ ( .D(n8178), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[395]) );
  SDFFR_X1 mem_reg_13__10_ ( .D(n8179), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[394]) );
  SDFFR_X1 mem_reg_13__9_ ( .D(n8180), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[393]) );
  SDFFR_X1 mem_reg_13__8_ ( .D(n8181), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[392]) );
  SDFFR_X1 mem_reg_13__7_ ( .D(n8182), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[391]) );
  SDFFR_X1 mem_reg_13__6_ ( .D(n8183), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[390]) );
  SDFFR_X1 mem_reg_13__5_ ( .D(n8184), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[389]) );
  SDFFR_X1 mem_reg_13__4_ ( .D(n8185), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[388]) );
  SDFFR_X1 mem_reg_13__3_ ( .D(n8186), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[387]) );
  SDFFR_X1 mem_reg_13__2_ ( .D(n8187), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[386]) );
  SDFFR_X1 mem_reg_13__1_ ( .D(n8188), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[385]) );
  SDFFR_X1 mem_reg_13__0_ ( .D(n8189), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[384]) );
  SDFFR_X1 mem_reg_14__29_ ( .D(n8195), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[445]) );
  SDFFR_X1 mem_reg_14__28_ ( .D(n8196), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[444]) );
  SDFFR_X1 mem_reg_14__27_ ( .D(n8197), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[443]) );
  SDFFR_X1 mem_reg_14__26_ ( .D(n8198), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[442]) );
  SDFFR_X1 mem_reg_14__25_ ( .D(n8199), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[441]) );
  SDFFR_X1 mem_reg_14__24_ ( .D(n8200), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[440]) );
  SDFFR_X1 mem_reg_14__16_ ( .D(n8208), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[432]) );
  SDFFR_X1 mem_reg_14__14_ ( .D(n8210), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[430]) );
  SDFFR_X1 mem_reg_14__13_ ( .D(n8211), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[429]) );
  SDFFR_X1 mem_reg_14__12_ ( .D(n8212), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[428]) );
  SDFFR_X1 mem_reg_14__11_ ( .D(n8213), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[427]) );
  SDFFR_X1 mem_reg_14__9_ ( .D(n8215), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[425]) );
  SDFFR_X1 mem_reg_14__8_ ( .D(n8216), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[424]) );
  SDFFR_X1 mem_reg_14__6_ ( .D(n8218), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[422]) );
  SDFFR_X1 mem_reg_14__4_ ( .D(n8220), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[420]) );
  SDFFR_X1 mem_reg_14__3_ ( .D(n8221), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[419]) );
  SDFFR_X1 mem_reg_14__2_ ( .D(n8222), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[418]) );
  SDFFR_X1 mem_reg_14__1_ ( .D(n8223), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[417]) );
  SDFFR_X1 mem_reg_14__0_ ( .D(n8224), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[416]) );
  SDFFR_X1 mem_reg_15__31_ ( .D(n8228), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[479]) );
  SDFFR_X1 mem_reg_15__30_ ( .D(n8229), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[478]) );
  SDFFR_X1 mem_reg_15__29_ ( .D(n8230), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[477]) );
  SDFFR_X1 mem_reg_15__28_ ( .D(n8231), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[476]) );
  SDFFR_X1 mem_reg_15__27_ ( .D(n8232), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[475]) );
  SDFFR_X1 mem_reg_15__26_ ( .D(n8233), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[474]) );
  SDFFR_X1 mem_reg_15__25_ ( .D(n8234), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[473]) );
  SDFFR_X1 mem_reg_15__24_ ( .D(n8235), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[472]) );
  SDFFR_X1 mem_reg_15__22_ ( .D(n8237), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[470]) );
  SDFFR_X1 mem_reg_15__18_ ( .D(n8241), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[466]) );
  SDFFR_X1 mem_reg_15__16_ ( .D(n8243), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[464]) );
  SDFFR_X1 mem_reg_15__15_ ( .D(n8244), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[463]) );
  SDFFR_X1 mem_reg_15__14_ ( .D(n8245), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[462]) );
  SDFFR_X1 mem_reg_15__13_ ( .D(n8246), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[461]) );
  SDFFR_X1 mem_reg_15__12_ ( .D(n8247), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[460]) );
  SDFFR_X1 mem_reg_15__11_ ( .D(n8248), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[459]) );
  SDFFR_X1 mem_reg_15__10_ ( .D(n8249), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[458]) );
  SDFFR_X1 mem_reg_15__9_ ( .D(n8250), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[457]) );
  SDFFR_X1 mem_reg_15__8_ ( .D(n8251), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[456]) );
  SDFFR_X1 mem_reg_15__7_ ( .D(n8252), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[455]) );
  SDFFR_X1 mem_reg_15__6_ ( .D(n8253), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[454]) );
  SDFFR_X1 mem_reg_15__5_ ( .D(n8254), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[453]) );
  SDFFR_X1 mem_reg_15__4_ ( .D(n8255), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[452]) );
  SDFFR_X1 mem_reg_15__3_ ( .D(n8256), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[451]) );
  SDFFR_X1 mem_reg_15__2_ ( .D(n8257), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[450]) );
  SDFFR_X1 mem_reg_15__1_ ( .D(n8258), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[449]) );
  SDFFR_X1 mem_reg_15__0_ ( .D(n8259), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[448]) );
  SDFFR_X1 mem_reg_16__29_ ( .D(n8265), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[509]) );
  SDFFR_X1 mem_reg_16__28_ ( .D(n8266), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[508]) );
  SDFFR_X1 mem_reg_16__27_ ( .D(n8267), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[507]) );
  SDFFR_X1 mem_reg_16__26_ ( .D(n8268), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[506]) );
  SDFFR_X1 mem_reg_16__25_ ( .D(n8269), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[505]) );
  SDFFR_X1 mem_reg_16__24_ ( .D(n8270), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[504]) );
  SDFFR_X1 mem_reg_16__16_ ( .D(n8278), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[496]) );
  SDFFR_X1 mem_reg_16__14_ ( .D(n8280), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[494]) );
  SDFFR_X1 mem_reg_16__13_ ( .D(n8281), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[493]) );
  SDFFR_X1 mem_reg_16__12_ ( .D(n8282), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[492]) );
  SDFFR_X1 mem_reg_16__11_ ( .D(n8283), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[491]) );
  SDFFR_X1 mem_reg_16__9_ ( .D(n8285), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[489]) );
  SDFFR_X1 mem_reg_16__8_ ( .D(n8286), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[488]) );
  SDFFR_X1 mem_reg_16__6_ ( .D(n8288), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[486]) );
  SDFFR_X1 mem_reg_16__5_ ( .D(n8289), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[485]) );
  SDFFR_X1 mem_reg_16__4_ ( .D(n8290), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[484]) );
  SDFFR_X1 mem_reg_16__3_ ( .D(n8291), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[483]) );
  SDFFR_X1 mem_reg_16__2_ ( .D(n8292), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[482]) );
  SDFFR_X1 mem_reg_16__1_ ( .D(n8293), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[481]) );
  SDFFR_X1 mem_reg_16__0_ ( .D(n8294), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[480]) );
  SDFFR_X1 mem_reg_17__29_ ( .D(n8300), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[541]) );
  SDFFR_X1 mem_reg_17__28_ ( .D(n8301), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[540]) );
  SDFFR_X1 mem_reg_17__27_ ( .D(n8302), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[539]) );
  SDFFR_X1 mem_reg_17__26_ ( .D(n8303), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[538]) );
  SDFFR_X1 mem_reg_17__25_ ( .D(n8304), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[537]) );
  SDFFR_X1 mem_reg_17__24_ ( .D(n8305), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[536]) );
  SDFFR_X1 mem_reg_17__16_ ( .D(n8313), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[528]) );
  SDFFR_X1 mem_reg_17__14_ ( .D(n8315), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[526]) );
  SDFFR_X1 mem_reg_17__13_ ( .D(n8316), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[525]) );
  SDFFR_X1 mem_reg_17__12_ ( .D(n8317), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[524]) );
  SDFFR_X1 mem_reg_17__11_ ( .D(n8318), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[523]) );
  SDFFR_X1 mem_reg_17__9_ ( .D(n8320), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[521]) );
  SDFFR_X1 mem_reg_17__8_ ( .D(n8321), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[520]) );
  SDFFR_X1 mem_reg_17__7_ ( .D(n8322), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[519]) );
  SDFFR_X1 mem_reg_17__6_ ( .D(n8323), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[518]) );
  SDFFR_X1 mem_reg_17__5_ ( .D(n8324), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[517]) );
  SDFFR_X1 mem_reg_17__4_ ( .D(n8325), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[516]) );
  SDFFR_X1 mem_reg_17__3_ ( .D(n8326), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[515]) );
  SDFFR_X1 mem_reg_17__2_ ( .D(n8327), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[514]) );
  SDFFR_X1 mem_reg_17__1_ ( .D(n8328), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[513]) );
  SDFFR_X1 mem_reg_17__0_ ( .D(n8329), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[512]) );
  SDFFR_X1 mem_reg_18__29_ ( .D(n8335), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[573]) );
  SDFFR_X1 mem_reg_18__28_ ( .D(n8336), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[572]) );
  SDFFR_X1 mem_reg_18__27_ ( .D(n8337), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[571]) );
  SDFFR_X1 mem_reg_18__26_ ( .D(n8338), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[570]) );
  SDFFR_X1 mem_reg_18__25_ ( .D(n8339), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[569]) );
  SDFFR_X1 mem_reg_18__24_ ( .D(n8340), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[568]) );
  SDFFR_X1 mem_reg_18__16_ ( .D(n8348), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[560]) );
  SDFFR_X1 mem_reg_18__14_ ( .D(n8351), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[558]) );
  SDFFR_X1 mem_reg_18__13_ ( .D(n8352), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[557]) );
  SDFFR_X1 mem_reg_18__12_ ( .D(n8353), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[556]) );
  SDFFR_X1 mem_reg_18__11_ ( .D(n8354), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[555]) );
  SDFFR_X1 mem_reg_18__9_ ( .D(n8356), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[553]) );
  SDFFR_X1 mem_reg_18__8_ ( .D(n8357), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[552]) );
  SDFFR_X1 mem_reg_18__6_ ( .D(n8359), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[550]) );
  SDFFR_X1 mem_reg_18__4_ ( .D(n8361), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[548]) );
  SDFFR_X1 mem_reg_18__3_ ( .D(n8362), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[547]) );
  SDFFR_X1 mem_reg_18__2_ ( .D(n8363), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[546]) );
  SDFFR_X1 mem_reg_18__1_ ( .D(n8364), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[545]) );
  SDFFR_X1 mem_reg_18__0_ ( .D(n8365), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[544]) );
  SDFFR_X1 mem_reg_19__29_ ( .D(n8371), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[605]) );
  SDFFR_X1 mem_reg_19__28_ ( .D(n8372), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[604]) );
  SDFFR_X1 mem_reg_19__27_ ( .D(n8373), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[603]) );
  SDFFR_X1 mem_reg_19__26_ ( .D(n8374), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[602]) );
  SDFFR_X1 mem_reg_19__25_ ( .D(n8375), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[601]) );
  SDFFR_X1 mem_reg_19__24_ ( .D(n8376), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[600]) );
  SDFFR_X1 mem_reg_19__16_ ( .D(n8384), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[592]) );
  SDFFR_X1 mem_reg_19__14_ ( .D(n8386), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[590]) );
  SDFFR_X1 mem_reg_19__13_ ( .D(n8387), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[589]) );
  SDFFR_X1 mem_reg_19__12_ ( .D(n8388), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[588]) );
  SDFFR_X1 mem_reg_19__11_ ( .D(n8389), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[587]) );
  SDFFR_X1 mem_reg_19__9_ ( .D(n8391), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[585]) );
  SDFFR_X1 mem_reg_19__8_ ( .D(n8392), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[584]) );
  SDFFR_X1 mem_reg_19__7_ ( .D(n8393), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[583]) );
  SDFFR_X1 mem_reg_19__6_ ( .D(n8394), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[582]) );
  SDFFR_X1 mem_reg_19__5_ ( .D(n8395), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[581]) );
  SDFFR_X1 mem_reg_19__4_ ( .D(n8396), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[580]) );
  SDFFR_X1 mem_reg_19__3_ ( .D(n8397), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[579]) );
  SDFFR_X1 mem_reg_19__2_ ( .D(n8398), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[578]) );
  SDFFR_X1 mem_reg_19__1_ ( .D(n8399), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[577]) );
  SDFFR_X1 mem_reg_19__0_ ( .D(n8400), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[576]) );
  SDFFR_X1 mem_reg_20__29_ ( .D(n8441), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[637]) );
  SDFFR_X1 mem_reg_20__28_ ( .D(n8442), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[636]) );
  SDFFR_X1 mem_reg_20__27_ ( .D(n8443), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[635]) );
  SDFFR_X1 mem_reg_20__26_ ( .D(n8444), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[634]) );
  SDFFR_X1 mem_reg_20__25_ ( .D(n8445), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[633]) );
  SDFFR_X1 mem_reg_20__24_ ( .D(n8446), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[632]) );
  SDFFR_X1 mem_reg_20__16_ ( .D(n8454), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[624]) );
  SDFFR_X1 mem_reg_20__14_ ( .D(n8456), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[622]) );
  SDFFR_X1 mem_reg_20__13_ ( .D(n8457), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[621]) );
  SDFFR_X1 mem_reg_20__12_ ( .D(n8458), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[620]) );
  SDFFR_X1 mem_reg_20__11_ ( .D(n8459), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[619]) );
  SDFFR_X1 mem_reg_20__9_ ( .D(n8461), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[617]) );
  SDFFR_X1 mem_reg_20__8_ ( .D(n8462), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[616]) );
  SDFFR_X1 mem_reg_20__6_ ( .D(n8464), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[614]) );
  SDFFR_X1 mem_reg_20__5_ ( .D(n8465), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[613]) );
  SDFFR_X1 mem_reg_20__4_ ( .D(n8466), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[612]) );
  SDFFR_X1 mem_reg_20__3_ ( .D(n8467), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[611]) );
  SDFFR_X1 mem_reg_20__2_ ( .D(n8468), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[610]) );
  SDFFR_X1 mem_reg_20__1_ ( .D(n8469), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[609]) );
  SDFFR_X1 mem_reg_20__0_ ( .D(n8470), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[608]) );
  SDFFR_X1 mem_reg_21__29_ ( .D(n8476), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[669]) );
  SDFFR_X1 mem_reg_21__28_ ( .D(n8477), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[668]) );
  SDFFR_X1 mem_reg_21__27_ ( .D(n8478), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[667]) );
  SDFFR_X1 mem_reg_21__26_ ( .D(n8479), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[666]) );
  SDFFR_X1 mem_reg_21__25_ ( .D(n8480), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[665]) );
  SDFFR_X1 mem_reg_21__24_ ( .D(n8481), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[664]) );
  SDFFR_X1 mem_reg_21__16_ ( .D(n8489), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[656]) );
  SDFFR_X1 mem_reg_21__14_ ( .D(n8491), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[654]) );
  SDFFR_X1 mem_reg_21__13_ ( .D(n8492), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[653]) );
  SDFFR_X1 mem_reg_21__12_ ( .D(n8493), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[652]) );
  SDFFR_X1 mem_reg_21__9_ ( .D(n8496), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[649]) );
  SDFFR_X1 mem_reg_21__8_ ( .D(n8497), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[648]) );
  SDFFR_X1 mem_reg_21__7_ ( .D(n8498), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[647]) );
  SDFFR_X1 mem_reg_21__6_ ( .D(n8499), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[646]) );
  SDFFR_X1 mem_reg_21__5_ ( .D(n8500), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[645]) );
  SDFFR_X1 mem_reg_21__4_ ( .D(n8501), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[644]) );
  SDFFR_X1 mem_reg_21__3_ ( .D(n8502), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[643]) );
  SDFFR_X1 mem_reg_21__2_ ( .D(n8503), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[642]) );
  SDFFR_X1 mem_reg_21__1_ ( .D(n8504), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[641]) );
  SDFFR_X1 mem_reg_21__0_ ( .D(n8505), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[640]) );
  SDFFR_X1 mem_reg_22__29_ ( .D(n8511), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[701]) );
  SDFFR_X1 mem_reg_22__28_ ( .D(n8512), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[700]) );
  SDFFR_X1 mem_reg_22__27_ ( .D(n8513), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[699]) );
  SDFFR_X1 mem_reg_22__26_ ( .D(n8514), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[698]) );
  SDFFR_X1 mem_reg_22__25_ ( .D(n8515), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[697]) );
  SDFFR_X1 mem_reg_22__24_ ( .D(n8516), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[696]) );
  SDFFR_X1 mem_reg_22__16_ ( .D(n8524), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[688]) );
  SDFFR_X1 mem_reg_22__14_ ( .D(n8526), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[686]) );
  SDFFR_X1 mem_reg_22__13_ ( .D(n8527), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[685]) );
  SDFFR_X1 mem_reg_22__12_ ( .D(n8528), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[684]) );
  SDFFR_X1 mem_reg_22__11_ ( .D(n8529), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[683]) );
  SDFFR_X1 mem_reg_22__9_ ( .D(n8531), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[681]) );
  SDFFR_X1 mem_reg_22__8_ ( .D(n8532), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[680]) );
  SDFFR_X1 mem_reg_22__7_ ( .D(n8533), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[679]) );
  SDFFR_X1 mem_reg_22__6_ ( .D(n8534), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[678]) );
  SDFFR_X1 mem_reg_22__5_ ( .D(n8535), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[677]) );
  SDFFR_X1 mem_reg_22__4_ ( .D(n8536), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[676]) );
  SDFFR_X1 mem_reg_22__3_ ( .D(n8537), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[675]) );
  SDFFR_X1 mem_reg_22__2_ ( .D(n8538), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[674]) );
  SDFFR_X1 mem_reg_22__1_ ( .D(n8539), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[673]) );
  SDFFR_X1 mem_reg_22__0_ ( .D(n8540), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[672]) );
  SDFFR_X1 mem_reg_23__29_ ( .D(n8546), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[733]) );
  SDFFR_X1 mem_reg_23__28_ ( .D(n8547), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[732]) );
  SDFFR_X1 mem_reg_23__27_ ( .D(n8548), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[731]) );
  SDFFR_X1 mem_reg_23__26_ ( .D(n8549), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[730]) );
  SDFFR_X1 mem_reg_23__25_ ( .D(n8550), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[729]) );
  SDFFR_X1 mem_reg_23__24_ ( .D(n8551), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[728]) );
  SDFFR_X1 mem_reg_23__16_ ( .D(n8559), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[720]) );
  SDFFR_X1 mem_reg_23__14_ ( .D(n8561), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[718]) );
  SDFFR_X1 mem_reg_23__13_ ( .D(n8562), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[717]) );
  SDFFR_X1 mem_reg_23__12_ ( .D(n8563), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[716]) );
  SDFFR_X1 mem_reg_23__11_ ( .D(n8564), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[715]) );
  SDFFR_X1 mem_reg_23__9_ ( .D(n8566), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[713]) );
  SDFFR_X1 mem_reg_23__8_ ( .D(n8567), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[712]) );
  SDFFR_X1 mem_reg_23__7_ ( .D(n8568), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[711]) );
  SDFFR_X1 mem_reg_23__6_ ( .D(n8569), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[710]) );
  SDFFR_X1 mem_reg_23__5_ ( .D(n8570), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[709]) );
  SDFFR_X1 mem_reg_23__4_ ( .D(n8571), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[708]) );
  SDFFR_X1 mem_reg_23__3_ ( .D(n8572), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[707]) );
  SDFFR_X1 mem_reg_23__2_ ( .D(n8573), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[706]) );
  SDFFR_X1 mem_reg_23__1_ ( .D(n8574), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[705]) );
  SDFFR_X1 mem_reg_23__0_ ( .D(n8575), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[704]) );
  SDFFR_X1 mem_reg_24__29_ ( .D(n8581), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[765]) );
  SDFFR_X1 mem_reg_24__19_ ( .D(n8591), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[755]) );
  SDFFR_X1 mem_reg_24__17_ ( .D(n8593), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[753]) );
  SDFFR_X1 mem_reg_24__16_ ( .D(n8594), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[752]) );
  SDFFR_X1 mem_reg_24__15_ ( .D(n8595), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[751]) );
  SDFFR_X1 mem_reg_24__13_ ( .D(n8597), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[749]) );
  SDFFR_X1 mem_reg_24__12_ ( .D(n8598), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[748]) );
  SDFFR_X1 mem_reg_24__11_ ( .D(n8599), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[747]) );
  SDFFR_X1 mem_reg_24__10_ ( .D(n8600), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[746]) );
  SDFFR_X1 mem_reg_24__9_ ( .D(n8601), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[745]) );
  SDFFR_X1 mem_reg_24__8_ ( .D(n8602), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[744]) );
  SDFFR_X1 mem_reg_24__6_ ( .D(n8604), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[742]) );
  SDFFR_X1 mem_reg_24__5_ ( .D(n8605), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[741]) );
  SDFFR_X1 mem_reg_24__4_ ( .D(n8606), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[740]) );
  SDFFR_X1 mem_reg_24__3_ ( .D(n8607), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[739]) );
  SDFFR_X1 mem_reg_24__2_ ( .D(n8608), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[738]) );
  SDFFR_X1 mem_reg_24__1_ ( .D(n8609), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[737]) );
  SDFFR_X1 mem_reg_24__0_ ( .D(n8610), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[736]) );
  SDFFR_X1 mem_reg_25__29_ ( .D(n8616), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[797]) );
  SDFFR_X1 mem_reg_25__16_ ( .D(n8628), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[784]) );
  SDFFR_X1 mem_reg_25__13_ ( .D(n8631), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[781]) );
  SDFFR_X1 mem_reg_25__12_ ( .D(n8632), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[780]) );
  SDFFR_X1 mem_reg_25__11_ ( .D(n8633), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[779]) );
  SDFFR_X1 mem_reg_25__10_ ( .D(n8634), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[778]) );
  SDFFR_X1 mem_reg_25__9_ ( .D(n8635), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[777]) );
  SDFFR_X1 mem_reg_25__8_ ( .D(n8636), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[776]) );
  SDFFR_X1 mem_reg_25__7_ ( .D(n8637), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[775]) );
  SDFFR_X1 mem_reg_25__6_ ( .D(n8638), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[774]) );
  SDFFR_X1 mem_reg_25__5_ ( .D(n8639), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[773]) );
  SDFFR_X1 mem_reg_25__4_ ( .D(n8640), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[772]) );
  SDFFR_X1 mem_reg_25__3_ ( .D(n8641), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[771]) );
  SDFFR_X1 mem_reg_25__2_ ( .D(n8642), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[770]) );
  SDFFR_X1 mem_reg_25__1_ ( .D(n8643), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[769]) );
  SDFFR_X1 mem_reg_25__0_ ( .D(n8644), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[768]) );
  SDFFR_X1 mem_reg_26__29_ ( .D(n8650), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[829]) );
  SDFFR_X1 mem_reg_26__16_ ( .D(n8663), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[816]) );
  SDFFR_X1 mem_reg_26__15_ ( .D(n8664), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[815]) );
  SDFFR_X1 mem_reg_26__13_ ( .D(n8666), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[813]) );
  SDFFR_X1 mem_reg_26__12_ ( .D(n8667), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[812]) );
  SDFFR_X1 mem_reg_26__11_ ( .D(n8668), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[811]) );
  SDFFR_X1 mem_reg_26__10_ ( .D(n8669), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[810]) );
  SDFFR_X1 mem_reg_26__9_ ( .D(n8670), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[809]) );
  SDFFR_X1 mem_reg_26__8_ ( .D(n8671), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[808]) );
  SDFFR_X1 mem_reg_26__6_ ( .D(n8673), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[806]) );
  SDFFR_X1 mem_reg_26__5_ ( .D(n8674), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[805]) );
  SDFFR_X1 mem_reg_26__4_ ( .D(n8675), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[804]) );
  SDFFR_X1 mem_reg_26__3_ ( .D(n8676), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[803]) );
  SDFFR_X1 mem_reg_26__2_ ( .D(n8677), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[802]) );
  SDFFR_X1 mem_reg_26__1_ ( .D(n8678), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[801]) );
  SDFFR_X1 mem_reg_26__0_ ( .D(n8679), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[800]) );
  SDFFR_X1 mem_reg_27__29_ ( .D(n8685), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[861]) );
  SDFFR_X1 mem_reg_27__28_ ( .D(n8686), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[860]) );
  SDFFR_X1 mem_reg_27__27_ ( .D(n8687), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[859]) );
  SDFFR_X1 mem_reg_27__26_ ( .D(n8688), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[858]) );
  SDFFR_X1 mem_reg_27__25_ ( .D(n8689), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[857]) );
  SDFFR_X1 mem_reg_27__24_ ( .D(n8690), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[856]) );
  SDFFR_X1 mem_reg_27__16_ ( .D(n8698), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[848]) );
  SDFFR_X1 mem_reg_27__14_ ( .D(n8700), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[846]) );
  SDFFR_X1 mem_reg_27__13_ ( .D(n8701), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[845]) );
  SDFFR_X1 mem_reg_27__12_ ( .D(n8702), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[844]) );
  SDFFR_X1 mem_reg_27__11_ ( .D(n8703), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[843]) );
  SDFFR_X1 mem_reg_27__9_ ( .D(n8705), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[841]) );
  SDFFR_X1 mem_reg_27__8_ ( .D(n8706), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[840]) );
  SDFFR_X1 mem_reg_27__7_ ( .D(n8707), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[839]) );
  SDFFR_X1 mem_reg_27__6_ ( .D(n8708), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[838]) );
  SDFFR_X1 mem_reg_27__5_ ( .D(n8709), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[837]) );
  SDFFR_X1 mem_reg_27__4_ ( .D(n8710), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[836]) );
  SDFFR_X1 mem_reg_27__3_ ( .D(n8711), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[835]) );
  SDFFR_X1 mem_reg_27__2_ ( .D(n8712), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[834]) );
  SDFFR_X1 mem_reg_27__1_ ( .D(n8713), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[833]) );
  SDFFR_X1 mem_reg_27__0_ ( .D(n8714), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[832]) );
  SDFFR_X1 mem_reg_28__29_ ( .D(n8720), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[893]) );
  SDFFR_X1 mem_reg_28__22_ ( .D(n8727), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[886]) );
  SDFFR_X1 mem_reg_28__16_ ( .D(n8733), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[880]) );
  SDFFR_X1 mem_reg_28__13_ ( .D(n8736), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[877]) );
  SDFFR_X1 mem_reg_28__12_ ( .D(n8737), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[876]) );
  SDFFR_X1 mem_reg_28__11_ ( .D(n8738), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[875]) );
  SDFFR_X1 mem_reg_28__10_ ( .D(n8739), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[874]) );
  SDFFR_X1 mem_reg_28__9_ ( .D(n8740), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[873]) );
  SDFFR_X1 mem_reg_28__8_ ( .D(n8741), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[872]) );
  SDFFR_X1 mem_reg_28__7_ ( .D(n8742), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[871]) );
  SDFFR_X1 mem_reg_28__6_ ( .D(n8743), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[870]) );
  SDFFR_X1 mem_reg_28__5_ ( .D(n8744), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[869]) );
  SDFFR_X1 mem_reg_28__4_ ( .D(n8745), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[868]) );
  SDFFR_X1 mem_reg_28__3_ ( .D(n8746), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[867]) );
  SDFFR_X1 mem_reg_28__2_ ( .D(n8747), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[866]) );
  SDFFR_X1 mem_reg_28__1_ ( .D(n8748), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[865]) );
  SDFFR_X1 mem_reg_28__0_ ( .D(n8749), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[864]) );
  SDFFR_X1 mem_reg_29__29_ ( .D(n8755), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[925]) );
  SDFFR_X1 mem_reg_29__28_ ( .D(n8756), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[924]) );
  SDFFR_X1 mem_reg_29__27_ ( .D(n8757), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[923]) );
  SDFFR_X1 mem_reg_29__26_ ( .D(n8758), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[922]) );
  SDFFR_X1 mem_reg_29__25_ ( .D(n8759), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[921]) );
  SDFFR_X1 mem_reg_29__24_ ( .D(n8760), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[920]) );
  SDFFR_X1 mem_reg_29__16_ ( .D(n8768), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[912]) );
  SDFFR_X1 mem_reg_29__14_ ( .D(n8770), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[910]) );
  SDFFR_X1 mem_reg_29__13_ ( .D(n8771), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[909]) );
  SDFFR_X1 mem_reg_29__12_ ( .D(n8772), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[908]) );
  SDFFR_X1 mem_reg_29__11_ ( .D(n8773), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[907]) );
  SDFFR_X1 mem_reg_29__9_ ( .D(n8775), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[905]) );
  SDFFR_X1 mem_reg_29__8_ ( .D(n8776), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[904]) );
  SDFFR_X1 mem_reg_29__7_ ( .D(n8777), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[903]) );
  SDFFR_X1 mem_reg_29__6_ ( .D(n8778), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[902]) );
  SDFFR_X1 mem_reg_29__5_ ( .D(n8779), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[901]) );
  SDFFR_X1 mem_reg_29__4_ ( .D(n8780), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[900]) );
  SDFFR_X1 mem_reg_29__3_ ( .D(n8781), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[899]) );
  SDFFR_X1 mem_reg_29__2_ ( .D(n8782), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[898]) );
  SDFFR_X1 mem_reg_29__1_ ( .D(n8783), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[897]) );
  SDFFR_X1 mem_reg_29__0_ ( .D(n8784), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[896]) );
  SDFFR_X1 mem_reg_30__29_ ( .D(n8825), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[957]) );
  SDFFR_X1 mem_reg_30__16_ ( .D(n8838), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[944]) );
  SDFFR_X1 mem_reg_30__13_ ( .D(n8841), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[941]) );
  SDFFR_X1 mem_reg_30__12_ ( .D(n8842), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[940]) );
  SDFFR_X1 mem_reg_30__11_ ( .D(n8843), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[939]) );
  SDFFR_X1 mem_reg_30__10_ ( .D(n8844), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[938]) );
  SDFFR_X1 mem_reg_30__9_ ( .D(n8845), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[937]) );
  SDFFR_X1 mem_reg_30__8_ ( .D(n8846), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[936]) );
  SDFFR_X1 mem_reg_30__7_ ( .D(n8847), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[935]) );
  SDFFR_X1 mem_reg_30__6_ ( .D(n8849), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[934]) );
  SDFFR_X1 mem_reg_30__5_ ( .D(n8850), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[933]) );
  SDFFR_X1 mem_reg_30__4_ ( .D(n8851), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[932]) );
  SDFFR_X1 mem_reg_30__3_ ( .D(n8852), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[931]) );
  SDFFR_X1 mem_reg_30__2_ ( .D(n8853), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[930]) );
  SDFFR_X1 mem_reg_30__1_ ( .D(n8854), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[929]) );
  SDFFR_X1 mem_reg_30__0_ ( .D(n8855), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[928]) );
  SDFFR_X1 mem_reg_31__31_ ( .D(n8859), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[991]) );
  SDFFR_X1 mem_reg_31__30_ ( .D(n8860), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[990]) );
  SDFFR_X1 mem_reg_31__29_ ( .D(n8862), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[989]) );
  SDFFR_X1 mem_reg_31__28_ ( .D(n8863), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[988]) );
  SDFFR_X1 mem_reg_31__27_ ( .D(n8864), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[987]) );
  SDFFR_X1 mem_reg_31__26_ ( .D(n8866), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[986]) );
  SDFFR_X1 mem_reg_31__25_ ( .D(n8868), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[985]) );
  SDFFR_X1 mem_reg_31__23_ ( .D(n8870), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[983]) );
  SDFFR_X1 mem_reg_31__22_ ( .D(n8872), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[982]) );
  SDFFR_X1 mem_reg_31__20_ ( .D(n8874), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[980]) );
  SDFFR_X1 mem_reg_31__19_ ( .D(n8876), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[979]) );
  SDFFR_X1 mem_reg_31__18_ ( .D(n8878), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[978]) );
  SDFFR_X1 mem_reg_31__17_ ( .D(n8880), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[977]) );
  SDFFR_X1 mem_reg_31__16_ ( .D(n8882), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[976]) );
  SDFFR_X1 mem_reg_31__15_ ( .D(n8884), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[975]) );
  SDFFR_X1 mem_reg_31__14_ ( .D(n8886), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[974]) );
  SDFFR_X1 mem_reg_31__13_ ( .D(n8888), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[973]) );
  SDFFR_X1 mem_reg_31__12_ ( .D(n8889), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[972]) );
  SDFFR_X1 mem_reg_31__11_ ( .D(n8891), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[971]) );
  SDFFR_X1 mem_reg_31__10_ ( .D(n8893), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[970]) );
  SDFFR_X1 mem_reg_31__9_ ( .D(n8895), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[969]) );
  SDFFR_X1 mem_reg_31__8_ ( .D(n8897), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[968]) );
  SDFFR_X1 mem_reg_31__7_ ( .D(n8899), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[967]) );
  SDFFR_X1 mem_reg_31__6_ ( .D(n8900), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[966]) );
  SDFFR_X1 mem_reg_31__5_ ( .D(n8901), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[965]) );
  SDFFR_X1 mem_reg_31__4_ ( .D(n8903), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[964]) );
  SDFFR_X1 mem_reg_31__3_ ( .D(n8905), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[963]) );
  SDFFR_X1 mem_reg_31__2_ ( .D(n8907), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[962]) );
  SDFFR_X1 mem_reg_31__1_ ( .D(n8909), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[961]) );
  SDFFR_X1 mem_reg_31__0_ ( .D(n8911), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[960]) );
  OR4_X2 U1696 ( .A1(n2194), .A2(n2193), .A3(n2192), .A4(n2191), .ZN(
        rdata_a_o[4]) );
  SDFFR_X2 mem_reg_1__28_ ( .D(n8407), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[28]) );
  SDFFR_X2 mem_reg_1__25_ ( .D(n8410), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[25]) );
  SDFFR_X2 mem_reg_1__24_ ( .D(n8411), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[24]) );
  SDFFR_X2 mem_reg_1__22_ ( .D(n8413), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[22]) );
  SDFFR_X2 mem_reg_1__21_ ( .D(n8414), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[21]) );
  SDFFR_X2 mem_reg_1__19_ ( .D(n8416), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[19]) );
  SDFFR_X2 mem_reg_1__17_ ( .D(n8418), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[17]) );
  SDFFR_X2 mem_reg_1__15_ ( .D(n8420), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[15]) );
  SDFFR_X2 mem_reg_1__0_ ( .D(n8435), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[0]) );
  SDFFR_X2 mem_reg_2__28_ ( .D(n8791), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[60]) );
  SDFFR_X2 mem_reg_2__25_ ( .D(n8794), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[57]) );
  SDFFR_X2 mem_reg_2__24_ ( .D(n8795), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[56]) );
  SDFFR_X2 mem_reg_2__22_ ( .D(n8797), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[54]) );
  SDFFR_X2 mem_reg_2__21_ ( .D(n8798), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[53]) );
  SDFFR_X2 mem_reg_2__19_ ( .D(n8800), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[51]) );
  SDFFR_X2 mem_reg_2__17_ ( .D(n8802), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[49]) );
  SDFFR_X2 mem_reg_2__0_ ( .D(n8819), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[32]) );
  SDFFR_X2 mem_reg_3__28_ ( .D(n8918), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[92]) );
  SDFFR_X2 mem_reg_3__25_ ( .D(n8921), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[89]) );
  SDFFR_X2 mem_reg_3__22_ ( .D(n8925), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[86]) );
  SDFFR_X2 mem_reg_3__21_ ( .D(n8926), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[85]) );
  SDFFR_X2 mem_reg_3__19_ ( .D(n8928), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[83]) );
  SDFFR_X2 mem_reg_3__17_ ( .D(n8930), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[81]) );
  SDFFR_X2 mem_reg_3__15_ ( .D(n8932), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[79]) );
  SDFFR_X2 mem_reg_3__0_ ( .D(n8947), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[64]) );
  SDFFR_X2 mem_reg_4__22_ ( .D(n8960), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[118]) );
  SDFFR_X2 mem_reg_4__21_ ( .D(n8961), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[117]) );
  SDFFR_X2 mem_reg_4__19_ ( .D(n8963), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[115]) );
  SDFFR_X2 mem_reg_4__17_ ( .D(n8965), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[113]) );
  SDFFR_X2 mem_reg_4__0_ ( .D(n8982), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[96]) );
  SDFFR_X2 mem_reg_5__28_ ( .D(n8989), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[156]) );
  SDFFR_X2 mem_reg_5__25_ ( .D(n8992), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[153]) );
  SDFFR_X2 mem_reg_5__22_ ( .D(n8995), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[150]) );
  SDFFR_X2 mem_reg_5__21_ ( .D(n8996), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[149]) );
  SDFFR_X2 mem_reg_5__19_ ( .D(n8998), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[147]) );
  SDFFR_X2 mem_reg_5__17_ ( .D(n9000), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[145]) );
  SDFFR_X2 mem_reg_5__0_ ( .D(n9017), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[128]) );
  SDFFR_X2 mem_reg_6__22_ ( .D(n9030), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[182]) );
  SDFFR_X2 mem_reg_6__19_ ( .D(n9034), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[179]) );
  SDFFR_X2 mem_reg_6__17_ ( .D(n9036), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[177]) );
  SDFFR_X2 mem_reg_6__0_ ( .D(n9053), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[160]) );
  SDFFR_X2 mem_reg_8__31_ ( .D(n9109), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[255]) );
  SDFFR_X2 mem_reg_8__30_ ( .D(n9110), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[254]) );
  SDFFR_X2 mem_reg_8__23_ ( .D(n9117), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[247]) );
  SDFFR_X2 mem_reg_8__22_ ( .D(n9118), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[246]) );
  SDFFR_X2 mem_reg_8__21_ ( .D(n9119), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[245]) );
  SDFFR_X2 mem_reg_8__20_ ( .D(n9120), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[244]) );
  SDFFR_X2 mem_reg_8__19_ ( .D(n9121), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[243]) );
  SDFFR_X2 mem_reg_8__18_ ( .D(n9122), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[242]) );
  SDFFR_X2 mem_reg_8__17_ ( .D(n9123), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[241]) );
  SDFFR_X2 mem_reg_8__15_ ( .D(n9125), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[239]) );
  SDFFR_X2 mem_reg_8__10_ ( .D(n9130), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[234]) );
  SDFFR_X2 mem_reg_8__0_ ( .D(n9140), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[224]) );
  SDFFR_X2 mem_reg_10__31_ ( .D(n8053), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[319]) );
  SDFFR_X2 mem_reg_10__30_ ( .D(n8054), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[318]) );
  SDFFR_X2 mem_reg_10__23_ ( .D(n8061), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[311]) );
  SDFFR_X2 mem_reg_10__22_ ( .D(n8062), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[310]) );
  SDFFR_X2 mem_reg_10__21_ ( .D(n8063), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[309]) );
  SDFFR_X2 mem_reg_10__20_ ( .D(n8064), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[308]) );
  SDFFR_X2 mem_reg_10__19_ ( .D(n8065), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[307]) );
  SDFFR_X2 mem_reg_10__18_ ( .D(n8066), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[306]) );
  SDFFR_X2 mem_reg_10__17_ ( .D(n8067), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[305]) );
  SDFFR_X2 mem_reg_10__15_ ( .D(n8069), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[303]) );
  SDFFR_X2 mem_reg_10__10_ ( .D(n8074), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[298]) );
  SDFFR_X2 mem_reg_10__0_ ( .D(n8084), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[288]) );
  SDFFR_X2 mem_reg_11__31_ ( .D(n8088), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[351]) );
  SDFFR_X2 mem_reg_11__30_ ( .D(n8089), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[350]) );
  SDFFR_X2 mem_reg_11__28_ ( .D(n8091), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[348]) );
  SDFFR_X2 mem_reg_11__27_ ( .D(n8092), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[347]) );
  SDFFR_X2 mem_reg_11__26_ ( .D(n8093), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[346]) );
  SDFFR_X2 mem_reg_11__25_ ( .D(n8094), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[345]) );
  SDFFR_X2 mem_reg_11__24_ ( .D(n8095), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[344]) );
  SDFFR_X2 mem_reg_11__23_ ( .D(n8096), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[343]) );
  SDFFR_X2 mem_reg_11__22_ ( .D(n8097), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[342]) );
  SDFFR_X2 mem_reg_11__21_ ( .D(n8098), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[341]) );
  SDFFR_X2 mem_reg_11__20_ ( .D(n8099), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[340]) );
  SDFFR_X2 mem_reg_11__19_ ( .D(n8100), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[339]) );
  SDFFR_X2 mem_reg_11__18_ ( .D(n8101), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[338]) );
  SDFFR_X2 mem_reg_11__17_ ( .D(n8102), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[337]) );
  SDFFR_X2 mem_reg_11__15_ ( .D(n8104), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[335]) );
  SDFFR_X2 mem_reg_11__0_ ( .D(n8119), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[320]) );
  SDFFR_X2 mem_reg_7__28_ ( .D(n9060), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[220]) );
  SDFFR_X2 mem_reg_7__25_ ( .D(n9064), .SI(1'b0), .SE(1'b0), .CK(n9106), .RN(
        rst_n), .Q(mem[217]) );
  SDFFR_X2 mem_reg_12__31_ ( .D(n8123), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[383]) );
  SDFFR_X2 mem_reg_12__30_ ( .D(n8124), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[382]) );
  SDFFR_X2 mem_reg_12__23_ ( .D(n8131), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[375]) );
  SDFFR_X2 mem_reg_12__22_ ( .D(n8132), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[374]) );
  SDFFR_X2 mem_reg_12__21_ ( .D(n8133), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[373]) );
  SDFFR_X2 mem_reg_12__20_ ( .D(n8134), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[372]) );
  SDFFR_X2 mem_reg_12__19_ ( .D(n8135), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[371]) );
  SDFFR_X2 mem_reg_12__18_ ( .D(n8136), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[370]) );
  SDFFR_X2 mem_reg_12__17_ ( .D(n8137), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[369]) );
  SDFFR_X2 mem_reg_12__15_ ( .D(n8139), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[367]) );
  SDFFR_X2 mem_reg_12__10_ ( .D(n8144), .SI(1'b0), .SE(1'b0), .CK(n8155), .RN(
        rst_n), .Q(mem[362]) );
  SDFFR_X2 mem_reg_13__30_ ( .D(n8159), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[414]) );
  SDFFR_X2 mem_reg_13__29_ ( .D(n8160), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[413]) );
  SDFFR_X2 mem_reg_13__28_ ( .D(n8161), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[412]) );
  SDFFR_X2 mem_reg_13__27_ ( .D(n8162), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[411]) );
  SDFFR_X2 mem_reg_13__26_ ( .D(n8163), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[410]) );
  SDFFR_X2 mem_reg_13__25_ ( .D(n8164), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[409]) );
  SDFFR_X2 mem_reg_13__24_ ( .D(n8165), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[408]) );
  SDFFR_X2 mem_reg_13__23_ ( .D(n8166), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[407]) );
  SDFFR_X2 mem_reg_13__22_ ( .D(n8167), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[406]) );
  SDFFR_X2 mem_reg_13__21_ ( .D(n8168), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[405]) );
  SDFFR_X2 mem_reg_13__20_ ( .D(n8169), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[404]) );
  SDFFR_X2 mem_reg_13__19_ ( .D(n8170), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[403]) );
  SDFFR_X2 mem_reg_13__18_ ( .D(n8171), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[402]) );
  SDFFR_X2 mem_reg_13__17_ ( .D(n8172), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[401]) );
  SDFFR_X2 mem_reg_13__15_ ( .D(n8174), .SI(1'b0), .SE(1'b0), .CK(n8190), .RN(
        rst_n), .Q(mem[399]) );
  SDFFR_X2 mem_reg_14__31_ ( .D(n8193), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[447]) );
  SDFFR_X2 mem_reg_14__30_ ( .D(n8194), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[446]) );
  SDFFR_X2 mem_reg_14__23_ ( .D(n8201), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[439]) );
  SDFFR_X2 mem_reg_14__22_ ( .D(n8202), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[438]) );
  SDFFR_X2 mem_reg_14__21_ ( .D(n8203), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[437]) );
  SDFFR_X2 mem_reg_14__20_ ( .D(n8204), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[436]) );
  SDFFR_X2 mem_reg_14__19_ ( .D(n8205), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[435]) );
  SDFFR_X2 mem_reg_14__18_ ( .D(n8206), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[434]) );
  SDFFR_X2 mem_reg_14__17_ ( .D(n8207), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[433]) );
  SDFFR_X2 mem_reg_14__15_ ( .D(n8209), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[431]) );
  SDFFR_X2 mem_reg_14__10_ ( .D(n8214), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[426]) );
  SDFFR_X2 mem_reg_16__31_ ( .D(n8263), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[511]) );
  SDFFR_X2 mem_reg_16__30_ ( .D(n8264), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[510]) );
  SDFFR_X2 mem_reg_16__23_ ( .D(n8271), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[503]) );
  SDFFR_X2 mem_reg_16__22_ ( .D(n8272), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[502]) );
  SDFFR_X2 mem_reg_16__21_ ( .D(n8273), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[501]) );
  SDFFR_X2 mem_reg_16__20_ ( .D(n8274), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[500]) );
  SDFFR_X2 mem_reg_16__19_ ( .D(n8275), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[499]) );
  SDFFR_X2 mem_reg_16__18_ ( .D(n8276), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[498]) );
  SDFFR_X2 mem_reg_16__17_ ( .D(n8277), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[497]) );
  SDFFR_X2 mem_reg_16__15_ ( .D(n8279), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[495]) );
  SDFFR_X2 mem_reg_16__10_ ( .D(n8284), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[490]) );
  SDFFR_X2 mem_reg_17__31_ ( .D(n8298), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[543]) );
  SDFFR_X2 mem_reg_17__30_ ( .D(n8299), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[542]) );
  SDFFR_X2 mem_reg_17__23_ ( .D(n8306), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[535]) );
  SDFFR_X2 mem_reg_17__22_ ( .D(n8307), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[534]) );
  SDFFR_X2 mem_reg_17__20_ ( .D(n8309), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[532]) );
  SDFFR_X2 mem_reg_17__19_ ( .D(n8310), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[531]) );
  SDFFR_X2 mem_reg_17__18_ ( .D(n8311), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[530]) );
  SDFFR_X2 mem_reg_17__17_ ( .D(n8312), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[529]) );
  SDFFR_X2 mem_reg_17__15_ ( .D(n8314), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[527]) );
  SDFFR_X2 mem_reg_17__10_ ( .D(n8319), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[522]) );
  SDFFR_X2 mem_reg_18__31_ ( .D(n8333), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[575]) );
  SDFFR_X2 mem_reg_18__30_ ( .D(n8334), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[574]) );
  SDFFR_X2 mem_reg_18__23_ ( .D(n8341), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[567]) );
  SDFFR_X2 mem_reg_18__22_ ( .D(n8342), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[566]) );
  SDFFR_X2 mem_reg_18__21_ ( .D(n8343), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[565]) );
  SDFFR_X2 mem_reg_18__20_ ( .D(n8344), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[564]) );
  SDFFR_X2 mem_reg_18__19_ ( .D(n8345), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[563]) );
  SDFFR_X2 mem_reg_18__18_ ( .D(n8346), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[562]) );
  SDFFR_X2 mem_reg_18__17_ ( .D(n8347), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[561]) );
  SDFFR_X2 mem_reg_18__15_ ( .D(n8350), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[559]) );
  SDFFR_X2 mem_reg_18__10_ ( .D(n8355), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[554]) );
  SDFFR_X2 mem_reg_19__31_ ( .D(n8369), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[607]) );
  SDFFR_X2 mem_reg_19__30_ ( .D(n8370), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[606]) );
  SDFFR_X2 mem_reg_19__23_ ( .D(n8377), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[599]) );
  SDFFR_X2 mem_reg_19__22_ ( .D(n8378), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[598]) );
  SDFFR_X2 mem_reg_19__20_ ( .D(n8380), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[596]) );
  SDFFR_X2 mem_reg_19__19_ ( .D(n8381), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[595]) );
  SDFFR_X2 mem_reg_19__18_ ( .D(n8382), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[594]) );
  SDFFR_X2 mem_reg_19__17_ ( .D(n8383), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[593]) );
  SDFFR_X2 mem_reg_19__15_ ( .D(n8385), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[591]) );
  SDFFR_X2 mem_reg_19__10_ ( .D(n8390), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[586]) );
  SDFFR_X2 mem_reg_20__31_ ( .D(n8439), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[639]) );
  SDFFR_X2 mem_reg_20__30_ ( .D(n8440), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[638]) );
  SDFFR_X2 mem_reg_20__23_ ( .D(n8447), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[631]) );
  SDFFR_X2 mem_reg_20__22_ ( .D(n8448), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[630]) );
  SDFFR_X2 mem_reg_20__20_ ( .D(n8450), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[628]) );
  SDFFR_X2 mem_reg_20__19_ ( .D(n8451), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[627]) );
  SDFFR_X2 mem_reg_20__18_ ( .D(n8452), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[626]) );
  SDFFR_X2 mem_reg_20__17_ ( .D(n8453), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[625]) );
  SDFFR_X2 mem_reg_20__15_ ( .D(n8455), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[623]) );
  SDFFR_X2 mem_reg_20__10_ ( .D(n8460), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[618]) );
  SDFFR_X2 mem_reg_21__31_ ( .D(n8474), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[671]) );
  SDFFR_X2 mem_reg_21__30_ ( .D(n8475), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[670]) );
  SDFFR_X2 mem_reg_21__23_ ( .D(n8482), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[663]) );
  SDFFR_X2 mem_reg_21__22_ ( .D(n8483), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[662]) );
  SDFFR_X2 mem_reg_21__21_ ( .D(n8484), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[661]) );
  SDFFR_X2 mem_reg_21__20_ ( .D(n8485), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[660]) );
  SDFFR_X2 mem_reg_21__19_ ( .D(n8486), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[659]) );
  SDFFR_X2 mem_reg_21__18_ ( .D(n8487), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[658]) );
  SDFFR_X2 mem_reg_21__17_ ( .D(n8488), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[657]) );
  SDFFR_X2 mem_reg_21__15_ ( .D(n8490), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[655]) );
  SDFFR_X2 mem_reg_21__10_ ( .D(n8495), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[650]) );
  SDFFR_X2 mem_reg_22__31_ ( .D(n8509), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[703]) );
  SDFFR_X2 mem_reg_22__30_ ( .D(n8510), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[702]) );
  SDFFR_X2 mem_reg_22__23_ ( .D(n8517), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[695]) );
  SDFFR_X2 mem_reg_22__22_ ( .D(n8518), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[694]) );
  SDFFR_X2 mem_reg_22__20_ ( .D(n8520), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[692]) );
  SDFFR_X2 mem_reg_22__19_ ( .D(n8521), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[691]) );
  SDFFR_X2 mem_reg_22__18_ ( .D(n8522), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[690]) );
  SDFFR_X2 mem_reg_22__17_ ( .D(n8523), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[689]) );
  SDFFR_X2 mem_reg_22__15_ ( .D(n8525), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[687]) );
  SDFFR_X2 mem_reg_22__10_ ( .D(n8530), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[682]) );
  SDFFR_X2 mem_reg_23__31_ ( .D(n8544), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[735]) );
  SDFFR_X2 mem_reg_23__30_ ( .D(n8545), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[734]) );
  SDFFR_X2 mem_reg_23__23_ ( .D(n8552), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[727]) );
  SDFFR_X2 mem_reg_23__22_ ( .D(n8553), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[726]) );
  SDFFR_X2 mem_reg_23__21_ ( .D(n8554), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[725]) );
  SDFFR_X2 mem_reg_23__20_ ( .D(n8555), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[724]) );
  SDFFR_X2 mem_reg_23__19_ ( .D(n8556), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[723]) );
  SDFFR_X2 mem_reg_23__18_ ( .D(n8557), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[722]) );
  SDFFR_X2 mem_reg_23__17_ ( .D(n8558), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[721]) );
  SDFFR_X2 mem_reg_23__15_ ( .D(n8560), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[719]) );
  SDFFR_X2 mem_reg_23__10_ ( .D(n8565), .SI(1'b0), .SE(1'b0), .CK(n8576), .RN(
        rst_n), .Q(mem[714]) );
  SDFFR_X2 mem_reg_24__31_ ( .D(n8579), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[767]) );
  SDFFR_X2 mem_reg_24__30_ ( .D(n8580), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[766]) );
  SDFFR_X2 mem_reg_24__27_ ( .D(n8583), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[763]) );
  SDFFR_X2 mem_reg_24__26_ ( .D(n8584), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[762]) );
  SDFFR_X2 mem_reg_24__24_ ( .D(n8586), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[760]) );
  SDFFR_X2 mem_reg_24__23_ ( .D(n8587), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[759]) );
  SDFFR_X2 mem_reg_24__22_ ( .D(n8588), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[758]) );
  SDFFR_X2 mem_reg_24__21_ ( .D(n8589), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[757]) );
  SDFFR_X2 mem_reg_24__20_ ( .D(n8590), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[756]) );
  SDFFR_X2 mem_reg_24__18_ ( .D(n8592), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[754]) );
  SDFFR_X2 mem_reg_24__14_ ( .D(n8596), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[750]) );
  SDFFR_X2 mem_reg_25__31_ ( .D(n8614), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[799]) );
  SDFFR_X2 mem_reg_25__30_ ( .D(n8615), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[798]) );
  SDFFR_X2 mem_reg_25__27_ ( .D(n8617), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[795]) );
  SDFFR_X2 mem_reg_25__26_ ( .D(n8618), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[794]) );
  SDFFR_X2 mem_reg_25__24_ ( .D(n8620), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[792]) );
  SDFFR_X2 mem_reg_25__23_ ( .D(n8621), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[791]) );
  SDFFR_X2 mem_reg_25__22_ ( .D(n8622), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[790]) );
  SDFFR_X2 mem_reg_25__21_ ( .D(n8623), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[789]) );
  SDFFR_X2 mem_reg_25__20_ ( .D(n8624), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[788]) );
  SDFFR_X2 mem_reg_25__19_ ( .D(n8625), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[787]) );
  SDFFR_X2 mem_reg_25__18_ ( .D(n8626), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[786]) );
  SDFFR_X2 mem_reg_25__17_ ( .D(n8627), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[785]) );
  SDFFR_X2 mem_reg_25__15_ ( .D(n8629), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[783]) );
  SDFFR_X2 mem_reg_25__14_ ( .D(n8630), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[782]) );
  SDFFR_X2 mem_reg_26__31_ ( .D(n8648), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[831]) );
  SDFFR_X2 mem_reg_26__30_ ( .D(n8649), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[830]) );
  SDFFR_X2 mem_reg_26__27_ ( .D(n8652), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[827]) );
  SDFFR_X2 mem_reg_26__26_ ( .D(n8653), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[826]) );
  SDFFR_X2 mem_reg_26__24_ ( .D(n8655), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[824]) );
  SDFFR_X2 mem_reg_26__23_ ( .D(n8656), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[823]) );
  SDFFR_X2 mem_reg_26__22_ ( .D(n8657), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[822]) );
  SDFFR_X2 mem_reg_26__21_ ( .D(n8658), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[821]) );
  SDFFR_X2 mem_reg_26__20_ ( .D(n8659), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[820]) );
  SDFFR_X2 mem_reg_26__19_ ( .D(n8660), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[819]) );
  SDFFR_X2 mem_reg_26__18_ ( .D(n8661), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[818]) );
  SDFFR_X2 mem_reg_26__17_ ( .D(n8662), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[817]) );
  SDFFR_X2 mem_reg_26__14_ ( .D(n8665), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[814]) );
  SDFFR_X2 mem_reg_27__31_ ( .D(n8683), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[863]) );
  SDFFR_X2 mem_reg_27__30_ ( .D(n8684), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[862]) );
  SDFFR_X2 mem_reg_27__23_ ( .D(n8691), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[855]) );
  SDFFR_X2 mem_reg_27__22_ ( .D(n8692), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[854]) );
  SDFFR_X2 mem_reg_27__20_ ( .D(n8694), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[852]) );
  SDFFR_X2 mem_reg_27__19_ ( .D(n8695), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[851]) );
  SDFFR_X2 mem_reg_27__18_ ( .D(n8696), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[850]) );
  SDFFR_X2 mem_reg_27__17_ ( .D(n8697), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[849]) );
  SDFFR_X2 mem_reg_27__15_ ( .D(n8699), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[847]) );
  SDFFR_X2 mem_reg_27__10_ ( .D(n8704), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[842]) );
  SDFFR_X2 mem_reg_28__31_ ( .D(n8718), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[895]) );
  SDFFR_X2 mem_reg_28__30_ ( .D(n8719), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[894]) );
  SDFFR_X2 mem_reg_28__27_ ( .D(n8722), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[891]) );
  SDFFR_X2 mem_reg_28__26_ ( .D(n8723), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[890]) );
  SDFFR_X2 mem_reg_28__24_ ( .D(n8725), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[888]) );
  SDFFR_X2 mem_reg_28__23_ ( .D(n8726), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[887]) );
  SDFFR_X2 mem_reg_28__21_ ( .D(n8728), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[885]) );
  SDFFR_X2 mem_reg_28__20_ ( .D(n8729), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[884]) );
  SDFFR_X2 mem_reg_28__19_ ( .D(n8730), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[883]) );
  SDFFR_X2 mem_reg_28__18_ ( .D(n8731), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[882]) );
  SDFFR_X2 mem_reg_28__17_ ( .D(n8732), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[881]) );
  SDFFR_X2 mem_reg_28__15_ ( .D(n8734), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[879]) );
  SDFFR_X2 mem_reg_28__14_ ( .D(n8735), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[878]) );
  SDFFR_X2 mem_reg_29__31_ ( .D(n8753), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[927]) );
  SDFFR_X2 mem_reg_29__30_ ( .D(n8754), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[926]) );
  SDFFR_X2 mem_reg_29__23_ ( .D(n8761), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[919]) );
  SDFFR_X2 mem_reg_29__22_ ( .D(n8762), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[918]) );
  SDFFR_X2 mem_reg_29__20_ ( .D(n8764), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[916]) );
  SDFFR_X2 mem_reg_29__19_ ( .D(n8765), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[915]) );
  SDFFR_X2 mem_reg_29__18_ ( .D(n8766), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[914]) );
  SDFFR_X2 mem_reg_29__17_ ( .D(n8767), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[913]) );
  SDFFR_X2 mem_reg_29__15_ ( .D(n8769), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[911]) );
  SDFFR_X2 mem_reg_29__10_ ( .D(n8774), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[906]) );
  SDFFR_X2 mem_reg_30__31_ ( .D(n8823), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[959]) );
  SDFFR_X2 mem_reg_30__30_ ( .D(n8824), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[958]) );
  SDFFR_X2 mem_reg_30__27_ ( .D(n8827), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[955]) );
  SDFFR_X2 mem_reg_30__26_ ( .D(n8828), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[954]) );
  SDFFR_X2 mem_reg_30__24_ ( .D(n8830), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[952]) );
  SDFFR_X2 mem_reg_30__23_ ( .D(n8831), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[951]) );
  SDFFR_X2 mem_reg_30__22_ ( .D(n8832), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[950]) );
  SDFFR_X2 mem_reg_30__21_ ( .D(n8833), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[949]) );
  SDFFR_X2 mem_reg_30__20_ ( .D(n8834), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[948]) );
  SDFFR_X2 mem_reg_30__19_ ( .D(n8835), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[947]) );
  SDFFR_X2 mem_reg_30__18_ ( .D(n8836), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[946]) );
  SDFFR_X2 mem_reg_30__17_ ( .D(n8837), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[945]) );
  SDFFR_X2 mem_reg_30__15_ ( .D(n8839), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[943]) );
  SDFFR_X2 mem_reg_30__14_ ( .D(n8840), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[942]) );
  SDFFR_X2 mem_reg_31__24_ ( .D(n8869), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[984]) );
  SDFFR_X2 mem_reg_31__21_ ( .D(n8873), .SI(1'b0), .SE(1'b0), .CK(n8912), .RN(
        rst_n), .Q(mem[981]) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_0 clk_gate_mem_reg_9__0_ ( 
        .CLK(clk), .EN(n9198), .ENCLK(n9196), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_1 clk_gate_mem_reg_8__0_ ( 
        .CLK(clk), .EN(n9143), .ENCLK(n9141), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_2 clk_gate_mem_reg_7__0_ ( 
        .CLK(clk), .EN(n9108), .ENCLK(n9106), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_3 clk_gate_mem_reg_6__0_ ( 
        .CLK(clk), .EN(n9056), .ENCLK(n9054), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_4 clk_gate_mem_reg_5__0_ ( 
        .CLK(clk), .EN(n9020), .ENCLK(n9018), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_5 clk_gate_mem_reg_4__0_ ( 
        .CLK(clk), .EN(n8985), .ENCLK(n8983), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_6 clk_gate_mem_reg_3__0_ ( 
        .CLK(clk), .EN(n8950), .ENCLK(n8948), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_7 clk_gate_mem_reg_31__0_ ( 
        .CLK(clk), .EN(n8914), .ENCLK(n8912), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_8 clk_gate_mem_reg_30__0_ ( 
        .CLK(clk), .EN(n8858), .ENCLK(n8856), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_9 clk_gate_mem_reg_2__0_ ( 
        .CLK(clk), .EN(n8822), .ENCLK(n8820), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_10 clk_gate_mem_reg_29__0_ ( 
        .CLK(clk), .EN(n8787), .ENCLK(n8785), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_11 clk_gate_mem_reg_28__0_ ( 
        .CLK(clk), .EN(n8752), .ENCLK(n8750), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_12 clk_gate_mem_reg_27__0_ ( 
        .CLK(clk), .EN(n8717), .ENCLK(n8715), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_13 clk_gate_mem_reg_26__0_ ( 
        .CLK(clk), .EN(n8682), .ENCLK(n8680), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_14 clk_gate_mem_reg_25__0_ ( 
        .CLK(clk), .EN(n8647), .ENCLK(n8645), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_15 clk_gate_mem_reg_24__0_ ( 
        .CLK(clk), .EN(n8613), .ENCLK(n8611), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_16 clk_gate_mem_reg_23__0_ ( 
        .CLK(clk), .EN(n8578), .ENCLK(n8576), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_17 clk_gate_mem_reg_22__0_ ( 
        .CLK(clk), .EN(n8543), .ENCLK(n8541), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_18 clk_gate_mem_reg_21__0_ ( 
        .CLK(clk), .EN(n8508), .ENCLK(n8506), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_19 clk_gate_mem_reg_20__0_ ( 
        .CLK(clk), .EN(n8473), .ENCLK(n8471), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_20 clk_gate_mem_reg_1__0_ ( 
        .CLK(clk), .EN(n8438), .ENCLK(n8436), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_21 clk_gate_mem_reg_19__0_ ( 
        .CLK(clk), .EN(n8403), .ENCLK(n8401), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_22 clk_gate_mem_reg_18__0_ ( 
        .CLK(clk), .EN(n8368), .ENCLK(n8366), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_23 clk_gate_mem_reg_17__0_ ( 
        .CLK(clk), .EN(n8332), .ENCLK(n8330), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_24 clk_gate_mem_reg_16__0_ ( 
        .CLK(clk), .EN(n8297), .ENCLK(n8295), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_25 clk_gate_mem_reg_15__0_ ( 
        .CLK(clk), .EN(n8262), .ENCLK(n8260), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_26 clk_gate_mem_reg_14__0_ ( 
        .CLK(clk), .EN(n8227), .ENCLK(n8225), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_27 clk_gate_mem_reg_13__0_ ( 
        .CLK(clk), .EN(n8192), .ENCLK(n8190), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_28 clk_gate_mem_reg_12__0_ ( 
        .CLK(clk), .EN(n8157), .ENCLK(n8155), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_29 clk_gate_mem_reg_11__0_ ( 
        .CLK(clk), .EN(n8122), .ENCLK(n8120), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0_30 clk_gate_mem_reg_10__0_ ( 
        .CLK(clk), .EN(n8087), .ENCLK(n8085), .TE(1'b0) );
  SDFFR_X2 mem_reg_24__25_ ( .D(n8585), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[761]) );
  SDFFR_X2 mem_reg_25__25_ ( .D(n8619), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[793]) );
  SDFFR_X2 mem_reg_26__25_ ( .D(n8654), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[825]) );
  SDFFR_X2 mem_reg_28__25_ ( .D(n8724), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[889]) );
  SDFFR_X2 mem_reg_30__25_ ( .D(n8829), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[953]) );
  SDFFR_X2 mem_reg_24__28_ ( .D(n8582), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[764]) );
  SDFFR_X2 mem_reg_25__28_ ( .D(n4800), .SI(1'b0), .SE(1'b0), .CK(n8645), .RN(
        rst_n), .Q(mem[796]) );
  SDFFR_X2 mem_reg_26__28_ ( .D(n8651), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[828]) );
  SDFFR_X2 mem_reg_28__28_ ( .D(n8721), .SI(1'b0), .SE(1'b0), .CK(n8750), .RN(
        rst_n), .Q(mem[892]) );
  SDFFR_X2 mem_reg_30__28_ ( .D(n8826), .SI(1'b0), .SE(1'b0), .CK(n8856), .RN(
        rst_n), .Q(mem[956]) );
  SDFFR_X2 mem_reg_1__27_ ( .D(n8408), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[27]) );
  SDFFR_X2 mem_reg_2__27_ ( .D(n8792), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[59]) );
  SDFFR_X2 mem_reg_3__27_ ( .D(n8919), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[91]) );
  SDFFR_X2 mem_reg_5__27_ ( .D(n8990), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[155]) );
  SDFFR_X2 mem_reg_15__17_ ( .D(n8242), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[465]) );
  SDFFR_X2 mem_reg_15__23_ ( .D(n8236), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[471]) );
  SDFFR_X2 mem_reg_15__20_ ( .D(n8239), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[468]) );
  SDFFR_X2 mem_reg_15__19_ ( .D(n8240), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[467]) );
  AND2_X2 U1773 ( .A1(n2260), .A2(n2259), .ZN(n2263) );
  SDFFR_X2 mem_reg_6__20_ ( .D(n9033), .SI(1'b0), .SE(1'b0), .CK(n9054), .RN(
        rst_n), .Q(mem[180]) );
  AND2_X4 U1011 ( .A1(n1631), .A2(n3770), .ZN(n1629) );
  SDFFR_X2 mem_reg_1__20_ ( .D(n8415), .SI(1'b0), .SE(1'b0), .CK(n8436), .RN(
        rst_n), .Q(mem[20]) );
  SDFFR_X2 mem_reg_2__20_ ( .D(n8799), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[52]) );
  SDFFR_X2 mem_reg_3__20_ ( .D(n8927), .SI(1'b0), .SE(1'b0), .CK(n8948), .RN(
        rst_n), .Q(mem[84]) );
  SDFFR_X2 mem_reg_5__20_ ( .D(n8997), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[148]) );
  SDFFR_X2 mem_reg_4__20_ ( .D(n8962), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[116]) );
  SDFFR_X2 mem_reg_5__23_ ( .D(n8994), .SI(1'b0), .SE(1'b0), .CK(n9018), .RN(
        rst_n), .Q(mem[151]) );
  SDFFR_X2 mem_reg_26__7_ ( .D(n8672), .SI(1'b0), .SE(1'b0), .CK(n8680), .RN(
        rst_n), .Q(mem[807]) );
  SDFFR_X2 mem_reg_24__7_ ( .D(n8603), .SI(1'b0), .SE(1'b0), .CK(n8611), .RN(
        rst_n), .Q(mem[743]) );
  SDFFR_X2 mem_reg_20__7_ ( .D(n8463), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[615]) );
  SDFFR_X2 mem_reg_18__7_ ( .D(n8358), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[551]) );
  SDFFR_X2 mem_reg_16__7_ ( .D(n8287), .SI(1'b0), .SE(1'b0), .CK(n8295), .RN(
        rst_n), .Q(mem[487]) );
  SDFFR_X2 mem_reg_14__7_ ( .D(n8217), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[423]) );
  SDFFR_X2 mem_reg_10__7_ ( .D(n8077), .SI(1'b0), .SE(1'b0), .CK(n8085), .RN(
        rst_n), .Q(mem[295]) );
  SDFFR_X2 mem_reg_8__7_ ( .D(n9133), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[231]) );
  SDFFR_X2 mem_reg_18__5_ ( .D(n8360), .SI(1'b0), .SE(1'b0), .CK(n8366), .RN(
        rst_n), .Q(mem[549]) );
  SDFFR_X2 mem_reg_14__5_ ( .D(n8219), .SI(1'b0), .SE(1'b0), .CK(n8225), .RN(
        rst_n), .Q(mem[421]) );
  SDFFR_X2 mem_reg_11__5_ ( .D(n8114), .SI(1'b0), .SE(1'b0), .CK(n8120), .RN(
        rst_n), .Q(mem[325]) );
  SDFFR_X2 mem_reg_8__5_ ( .D(n9135), .SI(1'b0), .SE(1'b0), .CK(n9141), .RN(
        rst_n), .Q(mem[229]) );
  SDFFR_X2 mem_reg_4__5_ ( .D(n8977), .SI(1'b0), .SE(1'b0), .CK(n8983), .RN(
        rst_n), .Q(mem[101]) );
  SDFFR_X2 mem_reg_2__5_ ( .D(n8814), .SI(1'b0), .SE(1'b0), .CK(n8820), .RN(
        rst_n), .Q(mem[37]) );
  SDFFR_X2 mem_reg_21__11_ ( .D(n8494), .SI(1'b0), .SE(1'b0), .CK(n8506), .RN(
        rst_n), .Q(mem[651]) );
  AND2_X1 U230 ( .A1(n1691), .A2(n1708), .ZN(n3210) );
  BUF_X1 U66 ( .A(n3092), .Z(n3593) );
  AND2_X2 U1103 ( .A1(n1705), .A2(n1708), .ZN(n2162) );
  BUF_X1 U1115 ( .A(n3131), .Z(n3578) );
  BUF_X1 U67 ( .A(n3092), .Z(n3363) );
  BUF_X1 U186 ( .A(n3195), .Z(n1088) );
  BUF_X2 U53 ( .A(n3188), .Z(n1070) );
  BUF_X1 U113 ( .A(n1811), .Z(n1025) );
  AND2_X2 U1018 ( .A1(n1631), .A2(n3845), .ZN(n1634) );
  BUF_X2 U56 ( .A(n3194), .Z(n1068) );
  BUF_X2 U77 ( .A(n3189), .Z(n1071) );
  BUF_X1 U114 ( .A(n1811), .Z(n1026) );
  BUF_X1 U104 ( .A(n2156), .Z(n1018) );
  BUF_X1 U115 ( .A(n1811), .Z(n1027) );
  BUF_X1 U76 ( .A(n2154), .Z(n3383) );
  BUF_X1 U64 ( .A(n3189), .Z(n3162) );
  BUF_X1 U52 ( .A(n3194), .Z(n3167) );
  BUF_X1 U91 ( .A(n3075), .Z(n1006) );
  BUF_X1 U63 ( .A(n3176), .Z(n1084) );
  BUF_X1 U100 ( .A(n3078), .Z(n1014) );
  BUF_X1 U59 ( .A(n3207), .Z(n996) );
  BUF_X1 U62 ( .A(n3176), .Z(n1085) );
  BUF_X1 U86 ( .A(n2146), .Z(n1081) );
  BUF_X1 U94 ( .A(n2148), .Z(n1009) );
  BUF_X1 U102 ( .A(n3078), .Z(n1016) );
  BUF_X1 U92 ( .A(n3075), .Z(n1007) );
  CLKBUF_X2 U150 ( .A(n1786), .Z(n1033) );
  INV_X2 U3153 ( .A(wdata_b_i[18]), .ZN(n4444) );
  BUF_X1 U13 ( .A(n3195), .Z(n1086) );
  BUF_X1 U55 ( .A(n2163), .Z(n3512) );
  BUF_X1 U68 ( .A(n2163), .Z(n3234) );
  BUF_X2 U229 ( .A(n2170), .Z(n3455) );
  BUF_X1 U105 ( .A(n2156), .Z(n1019) );
  CLKBUF_X2 U151 ( .A(n1750), .Z(n1055) );
  CLKBUF_X2 U149 ( .A(n1415), .Z(n1056) );
  CLKBUF_X2 U159 ( .A(n1394), .Z(n3010) );
  CLKBUF_X2 U141 ( .A(n1429), .Z(n1047) );
  CLKBUF_X2 U129 ( .A(n1511), .Z(n1040) );
  CLKBUF_X2 U161 ( .A(n2067), .Z(n2578) );
  CLKBUF_X2 U126 ( .A(n1516), .Z(n1050) );
  BUF_X1 U144 ( .A(n1740), .Z(n2062) );
  CLKBUF_X2 U134 ( .A(n1401), .Z(n1044) );
  BUF_X1 U143 ( .A(n1745), .Z(n2668) );
  BUF_X1 U145 ( .A(n1752), .Z(n2433) );
  CLKBUF_X2 U139 ( .A(n1431), .Z(n1052) );
  CLKBUF_X2 U135 ( .A(n1739), .Z(n1048) );
  BUF_X1 U148 ( .A(n1424), .Z(n2874) );
  BUF_X1 U125 ( .A(n1403), .Z(n2869) );
  CLKBUF_X2 U137 ( .A(n1738), .Z(n1049) );
  CLKBUF_X2 U127 ( .A(n1409), .Z(n1054) );
  CLKBUF_X2 U124 ( .A(n1751), .Z(n1045) );
  CLKBUF_X2 U131 ( .A(n1430), .Z(n1041) );
  CLKBUF_X2 U138 ( .A(n1396), .Z(n1051) );
  BUF_X1 U140 ( .A(n1461), .Z(n2705) );
  BUF_X1 U146 ( .A(n1395), .Z(n3016) );
  CLKBUF_X2 U160 ( .A(n1474), .Z(n2750) );
  CLKBUF_X2 U133 ( .A(n1776), .Z(n1046) );
  CLKBUF_X2 U132 ( .A(n1402), .Z(n1039) );
  CLKBUF_X2 U130 ( .A(n1781), .Z(n1042) );
  CLKBUF_X2 U142 ( .A(n1521), .Z(n1053) );
  BUF_X1 U128 ( .A(n1452), .Z(n3015) );
  CLKBUF_X2 U136 ( .A(n1408), .Z(n1043) );
  INV_X1 U3124 ( .A(wdata_b_i[7]), .ZN(n4422) );
  BUF_X2 U1042 ( .A(wdata_b_i[6]), .Z(n4420) );
  INV_X1 U1780 ( .A(wdata_b_i[1]), .ZN(n4410) );
  INV_X1 U3166 ( .A(wdata_b_i[23]), .ZN(n4452) );
  SDFFR_X2 mem_reg_15__21_ ( .D(n8238), .SI(1'b0), .SE(1'b0), .CK(n8260), .RN(
        rst_n), .Q(mem[469]) );
  SDFFR_X2 mem_reg_17__21_ ( .D(n8308), .SI(1'b0), .SE(1'b0), .CK(n8330), .RN(
        rst_n), .Q(mem[533]) );
  SDFFR_X2 mem_reg_19__21_ ( .D(n8379), .SI(1'b0), .SE(1'b0), .CK(n8401), .RN(
        rst_n), .Q(mem[597]) );
  SDFFR_X2 mem_reg_20__21_ ( .D(n8449), .SI(1'b0), .SE(1'b0), .CK(n8471), .RN(
        rst_n), .Q(mem[629]) );
  SDFFR_X2 mem_reg_22__21_ ( .D(n8519), .SI(1'b0), .SE(1'b0), .CK(n8541), .RN(
        rst_n), .Q(mem[693]) );
  SDFFR_X2 mem_reg_27__21_ ( .D(n8693), .SI(1'b0), .SE(1'b0), .CK(n8715), .RN(
        rst_n), .Q(mem[853]) );
  SDFFR_X2 mem_reg_29__21_ ( .D(n8763), .SI(1'b0), .SE(1'b0), .CK(n8785), .RN(
        rst_n), .Q(mem[917]) );
  BUF_X2 U90 ( .A(n3075), .Z(n1005) );
  BUF_X1 U65 ( .A(n2163), .Z(n3579) );
  BUF_X1 U16 ( .A(n3114), .Z(n3517) );
  BUF_X1 U101 ( .A(n3078), .Z(n1015) );
  BUF_X1 U14 ( .A(n2170), .Z(n3594) );
  BUF_X1 U93 ( .A(n2148), .Z(n1008) );
  INV_X1 U3 ( .A(n4037), .ZN(n8881) );
  CLKBUF_X2 U4 ( .A(n2146), .Z(n1082) );
  BUF_X1 U5 ( .A(n4452), .Z(n4385) );
  BUF_X1 U6 ( .A(wdata_b_i[8]), .Z(n4774) );
  BUF_X2 U7 ( .A(n3210), .Z(n4729) );
  BUF_X2 U8 ( .A(n3210), .Z(n4730) );
  CLKBUF_X1 U9 ( .A(n4043), .Z(n4004) );
  INV_X1 U10 ( .A(wdata_b_i[21]), .ZN(n4449) );
  INV_X1 U17 ( .A(n4470), .ZN(n4731) );
  INV_X1 U18 ( .A(n4795), .ZN(n4732) );
  INV_X1 U19 ( .A(n4441), .ZN(n4734) );
  BUF_X1 U20 ( .A(n2148), .Z(n1010) );
  BUF_X2 U21 ( .A(n1028), .Z(n4736) );
  BUF_X1 U22 ( .A(n3195), .Z(n1087) );
  AND2_X1 U23 ( .A1(raddr_a_i[0]), .A2(n4773), .ZN(n1717) );
  INV_X1 U24 ( .A(n4382), .ZN(n9068) );
  INV_X1 U25 ( .A(n4382), .ZN(n9159) );
  INV_X1 U26 ( .A(n4798), .ZN(n9178) );
  INV_X1 U27 ( .A(n4436), .ZN(n9172) );
  INV_X1 U28 ( .A(n4432), .ZN(n9085) );
  INV_X1 U29 ( .A(n4452), .ZN(n8871) );
  INV_X1 U30 ( .A(n4436), .ZN(n8887) );
  INV_X1 U31 ( .A(n4439), .ZN(n9081) );
  INV_X1 U32 ( .A(n4439), .ZN(n8885) );
  INV_X1 U33 ( .A(n4798), .ZN(n8894) );
  INV_X1 U34 ( .A(n4470), .ZN(n9146) );
  BUF_X1 U35 ( .A(n4043), .Z(n4382) );
  BUF_X1 U36 ( .A(wdata_b_i[29]), .Z(n4803) );
  INV_X1 U37 ( .A(n4804), .ZN(n9164) );
  INV_X1 U38 ( .A(n4004), .ZN(n4737) );
  INV_X1 U39 ( .A(n4426), .ZN(n9091) );
  INV_X1 U40 ( .A(n4424), .ZN(n8898) );
  BUF_X1 U41 ( .A(wdata_b_i[29]), .Z(n4796) );
  INV_X1 U42 ( .A(n4804), .ZN(n8877) );
  INV_X1 U43 ( .A(n4470), .ZN(n8861) );
  BUF_X1 U44 ( .A(wdata_b_i[31]), .Z(n4784) );
  INV_X1 U45 ( .A(n4785), .ZN(n9184) );
  INV_X1 U46 ( .A(n4412), .ZN(n9191) );
  INV_X1 U48 ( .A(n4408), .ZN(n9195) );
  INV_X1 U60 ( .A(wdata_b_i[24]), .ZN(n4047) );
  INV_X1 U69 ( .A(n4414), .ZN(n8906) );
  INV_X1 U78 ( .A(n4441), .ZN(n8349) );
  BUF_X1 U79 ( .A(wdata_b_i[31]), .Z(n4789) );
  INV_X1 U80 ( .A(n4410), .ZN(n8910) );
  BUF_X2 U82 ( .A(n2146), .Z(n1080) );
  INV_X2 U84 ( .A(n4751), .ZN(n4822) );
  INV_X2 U85 ( .A(n4759), .ZN(n4814) );
  INV_X2 U95 ( .A(n4760), .ZN(n4813) );
  INV_X2 U99 ( .A(n1624), .ZN(n4744) );
  INV_X2 U112 ( .A(n4752), .ZN(n4807) );
  INV_X2 U118 ( .A(n4747), .ZN(n4745) );
  INV_X2 U120 ( .A(n4749), .ZN(n4746) );
  AND2_X1 U122 ( .A1(n1689), .A2(n1691), .ZN(n2163) );
  OR2_X1 U123 ( .A1(n1688), .A2(raddr_a_i[3]), .ZN(n1696) );
  NAND2_X1 U156 ( .A1(raddr_a_i[1]), .A2(raddr_a_i[0]), .ZN(n1724) );
  NOR2_X1 U157 ( .A1(n1709), .A2(n1095), .ZN(n2147) );
  NAND2_X1 U162 ( .A1(raddr_c_i[1]), .A2(n1344), .ZN(n1364) );
  AND2_X2 U164 ( .A1(n3845), .A2(n1636), .ZN(n1640) );
  AND2_X2 U168 ( .A1(n3770), .A2(n1643), .ZN(n1617) );
  AND2_X2 U173 ( .A1(n3845), .A2(n1643), .ZN(n1647) );
  AND2_X2 U175 ( .A1(n3846), .A2(n3845), .ZN(n3851) );
  INV_X2 U176 ( .A(n4756), .ZN(n4809) );
  INV_X2 U180 ( .A(n4762), .ZN(n4811) );
  INV_X2 U181 ( .A(n4757), .ZN(n4808) );
  INV_X2 U182 ( .A(n4763), .ZN(n4810) );
  INV_X2 U183 ( .A(n4767), .ZN(n4817) );
  INV_X2 U184 ( .A(n4765), .ZN(n4819) );
  INV_X2 U185 ( .A(n4761), .ZN(n4812) );
  INV_X2 U187 ( .A(n4755), .ZN(n4820) );
  INV_X2 U188 ( .A(n4758), .ZN(n4815) );
  INV_X2 U189 ( .A(n4768), .ZN(n4816) );
  INV_X2 U190 ( .A(n4766), .ZN(n4818) );
  INV_X2 U191 ( .A(n4750), .ZN(n4823) );
  INV_X2 U192 ( .A(n4764), .ZN(n4821) );
  AND2_X1 U193 ( .A1(n3770), .A2(n1636), .ZN(n1624) );
  OR2_X1 U194 ( .A1(n2479), .A2(n2539), .ZN(n4747) );
  INV_X1 U195 ( .A(n4748), .ZN(n4825) );
  OR2_X1 U196 ( .A1(n1601), .A2(n2479), .ZN(n4748) );
  OR2_X1 U197 ( .A1(n2479), .A2(n1591), .ZN(n4749) );
  OR2_X1 U198 ( .A1(n2479), .A2(n2546), .ZN(n4750) );
  OR2_X1 U199 ( .A1(n1585), .A2(n2479), .ZN(n4751) );
  OR2_X1 U200 ( .A1(n2479), .A2(n1608), .ZN(n4752) );
  OR2_X1 U202 ( .A1(n2540), .A2(n2539), .ZN(n4753) );
  INV_X2 U203 ( .A(n4753), .ZN(n4826) );
  INV_X1 U204 ( .A(n4754), .ZN(n4824) );
  OR2_X1 U205 ( .A1(n2540), .A2(n2546), .ZN(n4754) );
  OR2_X1 U207 ( .A1(n1601), .A2(n2540), .ZN(n4755) );
  OR2_X1 U209 ( .A1(n2540), .A2(n1608), .ZN(n4756) );
  OR2_X1 U212 ( .A1(n2540), .A2(n1591), .ZN(n4757) );
  OR2_X1 U213 ( .A1(n2547), .A2(n1601), .ZN(n4758) );
  OR2_X1 U215 ( .A1(n2547), .A2(n2539), .ZN(n4759) );
  OR2_X1 U216 ( .A1(n2547), .A2(n2546), .ZN(n4760) );
  OR2_X1 U217 ( .A1(n1585), .A2(n2547), .ZN(n4761) );
  OR2_X1 U225 ( .A1(n2547), .A2(n1608), .ZN(n4762) );
  OR2_X1 U231 ( .A1(n2547), .A2(n1591), .ZN(n4763) );
  OR2_X1 U238 ( .A1(n3769), .A2(n2546), .ZN(n4764) );
  OR2_X1 U239 ( .A1(n3769), .A2(n1591), .ZN(n4765) );
  OR2_X1 U240 ( .A1(n3769), .A2(n1601), .ZN(n4766) );
  OR2_X1 U241 ( .A1(n3769), .A2(n1608), .ZN(n4767) );
  OR2_X1 U242 ( .A1(n1585), .A2(n3769), .ZN(n4768) );
  AND4_X1 U243 ( .A1(n2923), .A2(n2922), .A3(n2921), .A4(n2920), .ZN(n4769) );
  AND4_X1 U244 ( .A1(n2911), .A2(n2910), .A3(n2909), .A4(n2908), .ZN(n4770) );
  AND4_X1 U245 ( .A1(n2915), .A2(n2914), .A3(n2913), .A4(n2912), .ZN(n4771) );
  AND4_X1 U246 ( .A1(n2919), .A2(n2918), .A3(n2917), .A4(n2916), .ZN(n4772) );
  INV_X1 U247 ( .A(raddr_a_i[1]), .ZN(n4773) );
  OR2_X1 U248 ( .A1(n4444), .A2(n4757), .ZN(n5365) );
  INV_X1 U249 ( .A(n4441), .ZN(n8883) );
  INV_X1 U250 ( .A(n4799), .ZN(n4775) );
  INV_X1 U251 ( .A(n4799), .ZN(n4776) );
  OR2_X1 U252 ( .A1(n4799), .A2(n4777), .ZN(n5137) );
  INV_X1 U253 ( .A(n1647), .ZN(n4777) );
  INV_X1 U254 ( .A(n4799), .ZN(n9157) );
  INV_X1 U255 ( .A(n4422), .ZN(n8848) );
  OR2_X1 U256 ( .A1(n4002), .A2(n4778), .ZN(n5163) );
  INV_X1 U257 ( .A(n1640), .ZN(n4778) );
  OR2_X1 U258 ( .A1(n4444), .A2(n7797), .ZN(n5181) );
  INV_X1 U259 ( .A(n4422), .ZN(n4779) );
  INV_X1 U260 ( .A(n4422), .ZN(n4780) );
  INV_X1 U261 ( .A(n4422), .ZN(n9182) );
  INV_X1 U262 ( .A(n4430), .ZN(n4781) );
  INV_X1 U263 ( .A(n4430), .ZN(n8892) );
  INV_X1 U264 ( .A(wdata_b_i[25]), .ZN(n4011) );
  INV_X1 U265 ( .A(n4430), .ZN(n4782) );
  INV_X1 U266 ( .A(n4426), .ZN(n4783) );
  INV_X1 U267 ( .A(wdata_b_i[6]), .ZN(n4785) );
  INV_X1 U268 ( .A(n4410), .ZN(n4786) );
  INV_X1 U269 ( .A(n4410), .ZN(n9193) );
  INV_X1 U270 ( .A(n4004), .ZN(n4788) );
  INV_X1 U271 ( .A(n4416), .ZN(n4787) );
  INV_X1 U272 ( .A(n4416), .ZN(n8904) );
  OR2_X1 U273 ( .A1(n4385), .A2(n4753), .ZN(n4971) );
  NAND2_X1 U274 ( .A1(n4797), .A2(n3774), .ZN(n5143) );
  INV_X1 U275 ( .A(n4408), .ZN(n4790) );
  INV_X1 U276 ( .A(n4408), .ZN(n4791) );
  INV_X1 U277 ( .A(n4444), .ZN(n9076) );
  BUF_X1 U278 ( .A(n4447), .Z(n4002) );
  INV_X1 U279 ( .A(n4444), .ZN(n4792) );
  INV_X1 U280 ( .A(n4444), .ZN(n4793) );
  OR2_X1 U281 ( .A1(n4444), .A2(n4794), .ZN(n5173) );
  INV_X1 U282 ( .A(n3851), .ZN(n4794) );
  INV_X1 U283 ( .A(n4444), .ZN(n8879) );
  INV_X1 U284 ( .A(wdata_b_i[27]), .ZN(n4795) );
  INV_X1 U285 ( .A(n4799), .ZN(n4797) );
  INV_X1 U286 ( .A(n4040), .ZN(n9074) );
  INV_X2 U287 ( .A(n4434), .ZN(n9174) );
  INV_X1 U288 ( .A(wdata_b_i[10]), .ZN(n4798) );
  INV_X1 U289 ( .A(wdata_b_i[23]), .ZN(n4799) );
  OR2_X1 U290 ( .A1(n4801), .A2(n4802), .ZN(n4800) );
  AND2_X1 U291 ( .A1(wdata_b_i[28]), .A2(n1647), .ZN(n4801) );
  AND2_X1 U292 ( .A1(n4618), .A2(n7704), .ZN(n4802) );
  INV_X1 U293 ( .A(wdata_b_i[28]), .ZN(n4017) );
  INV_X1 U294 ( .A(wdata_b_i[19]), .ZN(n4804) );
  INV_X2 U295 ( .A(n4449), .ZN(n9070) );
  INV_X1 U296 ( .A(n4374), .ZN(n4805) );
  INV_X1 U297 ( .A(n4374), .ZN(n4806) );
  INV_X1 U298 ( .A(n4374), .ZN(n9168) );
  INV_X1 U299 ( .A(wdata_b_i[0]), .ZN(n4408) );
  INV_X1 U307 ( .A(n4002), .ZN(n9072) );
  NAND4_X1 U308 ( .A1(n4772), .A2(n4769), .A3(n4770), .A4(n4771), .ZN(
        rdata_a_o[1]) );
  OR2_X1 U309 ( .A1(n4040), .A2(n4753), .ZN(n4991) );
  INV_X1 U310 ( .A(n3774), .ZN(n4827) );
  AND2_X4 U311 ( .A1(n3846), .A2(n3770), .ZN(n3774) );
  INV_X2 U312 ( .A(n4444), .ZN(n9166) );
  OR2_X1 U313 ( .A1(n4374), .A2(n4753), .ZN(n5049) );
  BUF_X1 U314 ( .A(n4447), .Z(n4380) );
  INV_X2 U326 ( .A(n4047), .ZN(n8923) );
  NAND2_X1 U328 ( .A1(n4829), .A2(n4828), .ZN(n8053) );
  NAND2_X1 U854 ( .A1(n4477), .A2(n7362), .ZN(n4828) );
  NAND2_X1 U858 ( .A1(n4789), .A2(n4816), .ZN(n4829) );
  NAND2_X1 U866 ( .A1(n4831), .A2(n4830), .ZN(n8088) );
  NAND2_X1 U867 ( .A1(n4477), .A2(n7384), .ZN(n4830) );
  NAND2_X1 U868 ( .A1(n4784), .A2(n4822), .ZN(n4831) );
  NAND2_X1 U869 ( .A1(n4833), .A2(n4832), .ZN(n8298) );
  NAND2_X1 U871 ( .A1(n4477), .A2(n7494), .ZN(n4832) );
  NAND2_X1 U876 ( .A1(n4784), .A2(n4746), .ZN(n4833) );
  NAND2_X1 U877 ( .A1(n4835), .A2(n4834), .ZN(n8333) );
  NAND2_X1 U878 ( .A1(n4477), .A2(n7517), .ZN(n4834) );
  NAND2_X1 U879 ( .A1(n4784), .A2(n4817), .ZN(n4835) );
  NAND2_X1 U882 ( .A1(n4837), .A2(n4836), .ZN(n8369) );
  NAND2_X1 U888 ( .A1(n4477), .A2(n7539), .ZN(n4836) );
  NAND2_X1 U889 ( .A1(n4784), .A2(n4807), .ZN(n4837) );
  NAND2_X1 U890 ( .A1(n4839), .A2(n4838), .ZN(n8727) );
  NAND2_X1 U891 ( .A1(wdata_a_i[22]), .A2(n7783), .ZN(n4838) );
  NAND2_X1 U895 ( .A1(n9068), .A2(n1634), .ZN(n4839) );
  NAND2_X1 U898 ( .A1(n4841), .A2(n4840), .ZN(n8123) );
  NAND2_X1 U899 ( .A1(n4477), .A2(n7405), .ZN(n4840) );
  NAND2_X1 U900 ( .A1(n4784), .A2(n4815), .ZN(n4841) );
  NAND2_X1 U901 ( .A1(n4843), .A2(n4842), .ZN(n9109) );
  NAND2_X1 U902 ( .A1(n4477), .A2(n8008), .ZN(n4842) );
  NAND2_X1 U904 ( .A1(n4784), .A2(n4818), .ZN(n4843) );
  NAND2_X1 U908 ( .A1(n4845), .A2(n4844), .ZN(n8951) );
  NAND2_X1 U909 ( .A1(wdata_a_i[31]), .A2(n7914), .ZN(n4844) );
  NAND2_X1 U910 ( .A1(n4784), .A2(n4814), .ZN(n4845) );
  NAND2_X1 U911 ( .A1(n4847), .A2(n4846), .ZN(n9021) );
  NAND2_X1 U913 ( .A1(wdata_a_i[31]), .A2(n7959), .ZN(n4846) );
  NAND2_X1 U916 ( .A1(n4784), .A2(n4813), .ZN(n4847) );
  BUF_X2 U917 ( .A(n4037), .Z(n4374) );
  NAND2_X1 U918 ( .A1(n4849), .A2(n4848), .ZN(n8404) );
  NAND2_X1 U919 ( .A1(wdata_a_i[31]), .A2(n7562), .ZN(n4848) );
  NAND2_X1 U920 ( .A1(n4784), .A2(n4745), .ZN(n4849) );
  NAND2_X1 U923 ( .A1(n4851), .A2(n4850), .ZN(n8788) );
  NAND2_X1 U924 ( .A1(wdata_a_i[31]), .A2(n7822), .ZN(n4850) );
  NAND2_X1 U925 ( .A1(n4784), .A2(n4821), .ZN(n4851) );
  NAND2_X1 U926 ( .A1(n4853), .A2(n4852), .ZN(n8915) );
  NAND2_X1 U927 ( .A1(wdata_a_i[31]), .A2(n7892), .ZN(n4852) );
  NAND2_X1 U930 ( .A1(n4784), .A2(n4823), .ZN(n4853) );
  NAND2_X1 U931 ( .A1(n4855), .A2(n4854), .ZN(n8986) );
  NAND2_X1 U932 ( .A1(wdata_a_i[31]), .A2(n7937), .ZN(n4854) );
  NAND2_X1 U933 ( .A1(n4784), .A2(n4826), .ZN(n4855) );
  NAND2_X1 U934 ( .A1(n4857), .A2(n4856), .ZN(n8158) );
  NAND2_X1 U935 ( .A1(n4477), .A2(n7427), .ZN(n4856) );
  NAND2_X1 U941 ( .A1(n4784), .A2(n4820), .ZN(n4857) );
  NAND2_X1 U942 ( .A1(n4859), .A2(n4858), .ZN(n8069) );
  NAND2_X1 U943 ( .A1(wdata_a_i[15]), .A2(n7366), .ZN(n4858) );
  NAND2_X1 U944 ( .A1(n8885), .A2(n4816), .ZN(n4859) );
  NAND2_X1 U945 ( .A1(n4861), .A2(n4860), .ZN(n8104) );
  NAND2_X1 U948 ( .A1(wdata_a_i[15]), .A2(n7398), .ZN(n4860) );
  NAND2_X1 U949 ( .A1(n9081), .A2(n4822), .ZN(n4861) );
  NAND2_X1 U950 ( .A1(n4863), .A2(n4862), .ZN(n8139) );
  NAND2_X1 U951 ( .A1(wdata_a_i[15]), .A2(n7409), .ZN(n4862) );
  NAND2_X1 U952 ( .A1(n9081), .A2(n4815), .ZN(n4863) );
  NAND2_X1 U957 ( .A1(n4865), .A2(n4864), .ZN(n8174) );
  NAND2_X1 U958 ( .A1(wdata_a_i[15]), .A2(n7442), .ZN(n4864) );
  NAND2_X1 U959 ( .A1(n9081), .A2(n4820), .ZN(n4865) );
  NAND2_X1 U960 ( .A1(n4867), .A2(n4866), .ZN(n8209) );
  NAND2_X1 U961 ( .A1(wdata_a_i[15]), .A2(n7453), .ZN(n4866) );
  NAND2_X1 U962 ( .A1(n8885), .A2(n4812), .ZN(n4867) );
  NAND2_X1 U965 ( .A1(n4869), .A2(n4868), .ZN(n8279) );
  NAND2_X1 U966 ( .A1(wdata_a_i[15]), .A2(n7476), .ZN(n4868) );
  NAND2_X1 U967 ( .A1(n8885), .A2(n4819), .ZN(n4869) );
  NAND2_X1 U968 ( .A1(n4871), .A2(n4870), .ZN(n8314) );
  NAND2_X1 U969 ( .A1(wdata_a_i[15]), .A2(n7499), .ZN(n4870) );
  NAND2_X1 U972 ( .A1(n9081), .A2(n4746), .ZN(n4871) );
  NAND2_X1 U973 ( .A1(n4873), .A2(n4872), .ZN(n8350) );
  NAND2_X1 U974 ( .A1(wdata_a_i[15]), .A2(n7521), .ZN(n4872) );
  NAND2_X1 U975 ( .A1(n9081), .A2(n4817), .ZN(n4873) );
  NAND2_X1 U976 ( .A1(n4875), .A2(n4874), .ZN(n8385) );
  NAND2_X1 U979 ( .A1(wdata_a_i[15]), .A2(n7544), .ZN(n4874) );
  NAND2_X1 U980 ( .A1(n9081), .A2(n4807), .ZN(n4875) );
  NAND2_X1 U981 ( .A1(n4877), .A2(n4876), .ZN(n8484) );
  NAND2_X1 U982 ( .A1(wdata_a_i[21]), .A2(n7610), .ZN(n4876) );
  NAND2_X1 U983 ( .A1(wdata_b_i[21]), .A2(n4808), .ZN(n4877) );
  NAND2_X1 U986 ( .A1(n4879), .A2(n4878), .ZN(n8932) );
  NAND2_X1 U987 ( .A1(wdata_a_i[15]), .A2(n7907), .ZN(n4878) );
  NAND2_X1 U988 ( .A1(n8885), .A2(n4823), .ZN(n4879) );
  NAND2_X1 U989 ( .A1(n4881), .A2(n4880), .ZN(n9125) );
  NAND2_X1 U992 ( .A1(wdata_a_i[15]), .A2(n8012), .ZN(n4880) );
  NAND2_X1 U997 ( .A1(n8885), .A2(n4818), .ZN(n4881) );
  NAND2_X1 U998 ( .A1(n4883), .A2(n4882), .ZN(n8623) );
  NAND2_X1 U999 ( .A1(wdata_a_i[21]), .A2(n7712), .ZN(n4882) );
  NAND2_X1 U1000 ( .A1(n9070), .A2(n1647), .ZN(n4883) );
  NAND2_X1 U1003 ( .A1(n4885), .A2(n4884), .ZN(n8728) );
  NAND2_X1 U1005 ( .A1(wdata_a_i[21]), .A2(n7784), .ZN(n4884) );
  NAND2_X1 U1007 ( .A1(n9070), .A2(n1634), .ZN(n4885) );
  NAND2_X1 U1008 ( .A1(n4887), .A2(n4886), .ZN(n8833) );
  NAND2_X1 U1009 ( .A1(wdata_a_i[21]), .A2(n7855), .ZN(n4886) );
  NAND2_X1 U1013 ( .A1(n9070), .A2(n1629), .ZN(n4887) );
  NAND2_X1 U1014 ( .A1(n4889), .A2(n4888), .ZN(n8873) );
  NAND2_X1 U1015 ( .A1(wdata_a_i[21]), .A2(n7891), .ZN(n4888) );
  NAND2_X1 U1016 ( .A1(n9070), .A2(n1624), .ZN(n4889) );
  NAND2_X1 U1017 ( .A1(n4891), .A2(n4890), .ZN(n8972) );
  NAND2_X1 U1020 ( .A1(wdata_a_i[10]), .A2(n7921), .ZN(n4890) );
  NAND2_X1 U1021 ( .A1(n8894), .A2(n4814), .ZN(n4891) );
  NAND2_X1 U1022 ( .A1(n4893), .A2(n4892), .ZN(n9043) );
  NAND2_X1 U1023 ( .A1(wdata_a_i[10]), .A2(n7967), .ZN(n4892) );
  NAND2_X1 U1024 ( .A1(n8894), .A2(n4813), .ZN(n4893) );
  NAND2_X1 U1025 ( .A1(n4895), .A2(n4894), .ZN(n8420) );
  NAND2_X1 U1029 ( .A1(wdata_a_i[15]), .A2(n7577), .ZN(n4894) );
  NAND2_X1 U1030 ( .A1(n8885), .A2(n4745), .ZN(n4895) );
  NAND2_X1 U1031 ( .A1(n4897), .A2(n4896), .ZN(n8804) );
  NAND2_X1 U1032 ( .A1(wdata_a_i[15]), .A2(n7837), .ZN(n4896) );
  NAND2_X1 U1033 ( .A1(n8885), .A2(n4821), .ZN(n4897) );
  NAND2_X1 U1037 ( .A1(n4899), .A2(n4898), .ZN(n8967) );
  NAND2_X1 U1039 ( .A1(wdata_a_i[15]), .A2(n7919), .ZN(n4898) );
  NAND2_X1 U1040 ( .A1(n9081), .A2(n4814), .ZN(n4899) );
  NAND2_X1 U1041 ( .A1(n4901), .A2(n4900), .ZN(n9002) );
  NAND2_X1 U1043 ( .A1(wdata_a_i[15]), .A2(n7952), .ZN(n4900) );
  NAND2_X1 U1044 ( .A1(wdata_b_i[15]), .A2(n4826), .ZN(n4901) );
  NAND2_X1 U1045 ( .A1(n4903), .A2(n4902), .ZN(n9038) );
  NAND2_X1 U1046 ( .A1(wdata_a_i[15]), .A2(n7965), .ZN(n4902) );
  NAND2_X1 U1047 ( .A1(n8885), .A2(n4813), .ZN(n4903) );
  NAND2_X1 U1048 ( .A1(n4905), .A2(n4904), .ZN(n9059) );
  NAND2_X1 U1049 ( .A1(n4468), .A2(n7986), .ZN(n4904) );
  NAND2_X1 U1050 ( .A1(n4803), .A2(n4824), .ZN(n4905) );
  NAND2_X1 U1051 ( .A1(n4907), .A2(n4906), .ZN(n8063) );
  NAND2_X1 U1052 ( .A1(wdata_a_i[21]), .A2(n7364), .ZN(n4906) );
  NAND2_X1 U1053 ( .A1(wdata_b_i[21]), .A2(n4816), .ZN(n4907) );
  NAND2_X1 U1054 ( .A1(n4909), .A2(n4908), .ZN(n8074) );
  NAND2_X1 U1055 ( .A1(wdata_a_i[10]), .A2(n7368), .ZN(n4908) );
  NAND2_X1 U1056 ( .A1(n9178), .A2(n4816), .ZN(n4909) );
  NAND2_X1 U1057 ( .A1(n4911), .A2(n4910), .ZN(n8417) );
  NAND2_X1 U1058 ( .A1(wdata_a_i[18]), .A2(n7573), .ZN(n4910) );
  NAND2_X1 U1059 ( .A1(n9076), .A2(n4745), .ZN(n4911) );
  NAND2_X1 U1060 ( .A1(n4913), .A2(n4912), .ZN(n8801) );
  NAND2_X1 U1061 ( .A1(wdata_a_i[18]), .A2(n7833), .ZN(n4912) );
  NAND2_X1 U1062 ( .A1(n9076), .A2(n4821), .ZN(n4913) );
  NAND2_X1 U1063 ( .A1(n4915), .A2(n4914), .ZN(n8926) );
  NAND2_X1 U1064 ( .A1(wdata_a_i[21]), .A2(n7902), .ZN(n4914) );
  NAND2_X1 U1065 ( .A1(n9032), .A2(n4823), .ZN(n4915) );
  NAND2_X1 U1066 ( .A1(n4917), .A2(n4916), .ZN(n8929) );
  NAND2_X1 U1067 ( .A1(wdata_a_i[18]), .A2(n7903), .ZN(n4916) );
  NAND2_X1 U1068 ( .A1(n9076), .A2(n4823), .ZN(n4917) );
  NAND2_X1 U1069 ( .A1(n4919), .A2(n4918), .ZN(n8961) );
  NAND2_X1 U1070 ( .A1(wdata_a_i[21]), .A2(n7916), .ZN(n4918) );
  NAND2_X1 U1071 ( .A1(n9070), .A2(n4814), .ZN(n4919) );
  NAND2_X1 U1072 ( .A1(n4921), .A2(n4920), .ZN(n8964) );
  NAND2_X1 U1073 ( .A1(wdata_a_i[18]), .A2(n7917), .ZN(n4920) );
  NAND2_X1 U1074 ( .A1(n9076), .A2(n4814), .ZN(n4921) );
  NAND2_X1 U1102 ( .A1(n4923), .A2(n4922), .ZN(n8996) );
  NAND2_X1 U1107 ( .A1(wdata_a_i[21]), .A2(n7947), .ZN(n4922) );
  NAND2_X1 U1113 ( .A1(n9070), .A2(n4826), .ZN(n4923) );
  NAND2_X1 U1114 ( .A1(n4925), .A2(n4924), .ZN(n8999) );
  NAND2_X1 U1192 ( .A1(wdata_a_i[18]), .A2(n7948), .ZN(n4924) );
  NAND2_X1 U1193 ( .A1(n9166), .A2(n4826), .ZN(n4925) );
  NAND2_X1 U1194 ( .A1(n4927), .A2(n4926), .ZN(n9035) );
  NAND2_X1 U1195 ( .A1(wdata_a_i[18]), .A2(n7963), .ZN(n4926) );
  NAND2_X1 U1196 ( .A1(n9166), .A2(n4813), .ZN(n4927) );
  NAND2_X1 U1197 ( .A1(n4929), .A2(n4928), .ZN(n8144) );
  NAND2_X1 U1198 ( .A1(wdata_a_i[10]), .A2(n7411), .ZN(n4928) );
  NAND2_X1 U1199 ( .A1(n9178), .A2(n4815), .ZN(n4929) );
  NAND2_X1 U1200 ( .A1(n4931), .A2(n4930), .ZN(n8214) );
  NAND2_X1 U1201 ( .A1(wdata_a_i[10]), .A2(n7455), .ZN(n4930) );
  NAND2_X1 U1202 ( .A1(n9178), .A2(n4812), .ZN(n4931) );
  NAND2_X1 U1203 ( .A1(n4933), .A2(n4932), .ZN(n8284) );
  NAND2_X1 U1204 ( .A1(wdata_a_i[10]), .A2(n7478), .ZN(n4932) );
  NAND2_X1 U1205 ( .A1(n9178), .A2(n4819), .ZN(n4933) );
  NAND2_X1 U1206 ( .A1(n4935), .A2(n4934), .ZN(n8319) );
  NAND2_X1 U1207 ( .A1(wdata_a_i[10]), .A2(n7501), .ZN(n4934) );
  NAND2_X1 U1208 ( .A1(n9178), .A2(n4746), .ZN(n4935) );
  NAND2_X1 U1209 ( .A1(n4937), .A2(n4936), .ZN(n8355) );
  NAND2_X1 U1210 ( .A1(wdata_a_i[10]), .A2(n7523), .ZN(n4936) );
  NAND2_X1 U1211 ( .A1(n9178), .A2(n4817), .ZN(n4937) );
  NAND2_X1 U1212 ( .A1(n4939), .A2(n4938), .ZN(n8390) );
  NAND2_X1 U1213 ( .A1(wdata_a_i[10]), .A2(n7546), .ZN(n4938) );
  NAND2_X1 U1214 ( .A1(n9178), .A2(n4807), .ZN(n4939) );
  NAND2_X1 U1215 ( .A1(n4941), .A2(n4940), .ZN(n8415) );
  NAND2_X1 U1216 ( .A1(wdata_a_i[20]), .A2(n7572), .ZN(n4940) );
  NAND2_X1 U1217 ( .A1(n9072), .A2(n4745), .ZN(n4941) );
  NAND2_X1 U1218 ( .A1(n4943), .A2(n4942), .ZN(n8799) );
  NAND2_X1 U1219 ( .A1(wdata_a_i[20]), .A2(n7832), .ZN(n4942) );
  NAND2_X1 U1220 ( .A1(n8875), .A2(n4821), .ZN(n4943) );
  NAND2_X1 U1221 ( .A1(n4945), .A2(n4944), .ZN(n8927) );
  NAND2_X1 U1436 ( .A1(wdata_a_i[20]), .A2(n7902), .ZN(n4944) );
  NAND2_X1 U1437 ( .A1(n9162), .A2(n4823), .ZN(n4945) );
  NAND2_X1 U1438 ( .A1(n4947), .A2(n4946), .ZN(n8997) );
  NAND2_X1 U1439 ( .A1(wdata_a_i[20]), .A2(n7947), .ZN(n4946) );
  NAND2_X1 U1440 ( .A1(n8875), .A2(n4826), .ZN(n4947) );
  NAND2_X1 U1441 ( .A1(n4949), .A2(n4948), .ZN(n9130) );
  NAND2_X1 U1442 ( .A1(wdata_a_i[10]), .A2(n8014), .ZN(n4948) );
  NAND2_X1 U1443 ( .A1(n9178), .A2(n4818), .ZN(n4949) );
  NAND2_X1 U1444 ( .A1(n4951), .A2(n4950), .ZN(n8406) );
  NAND2_X1 U1445 ( .A1(wdata_a_i[29]), .A2(n7564), .ZN(n4950) );
  NAND2_X1 U1446 ( .A1(n4803), .A2(n4745), .ZN(n4951) );
  NAND2_X1 U1447 ( .A1(n4953), .A2(n4952), .ZN(n8790) );
  NAND2_X1 U1448 ( .A1(wdata_a_i[29]), .A2(n7824), .ZN(n4952) );
  NAND2_X1 U1449 ( .A1(n4803), .A2(n4821), .ZN(n4953) );
  NAND2_X1 U1450 ( .A1(n4955), .A2(n4954), .ZN(n8988) );
  NAND2_X1 U1451 ( .A1(wdata_a_i[29]), .A2(n7939), .ZN(n4954) );
  NAND2_X1 U1452 ( .A1(n4803), .A2(n4826), .ZN(n4955) );
  NAND2_X1 U1453 ( .A1(n4957), .A2(n4956), .ZN(n8090) );
  NAND2_X1 U1454 ( .A1(n4468), .A2(n7386), .ZN(n4956) );
  NAND2_X1 U1455 ( .A1(n4803), .A2(n4822), .ZN(n4957) );
  NAND2_X1 U1456 ( .A1(n4959), .A2(n4958), .ZN(n8917) );
  NAND2_X1 U1457 ( .A1(n4468), .A2(n7893), .ZN(n4958) );
  NAND2_X1 U1458 ( .A1(n4803), .A2(n4823), .ZN(n4959) );
  NAND2_X1 U1459 ( .A1(n4961), .A2(n4960), .ZN(n8412) );
  NAND2_X1 U1460 ( .A1(wdata_a_i[23]), .A2(n7571), .ZN(n4960) );
  NAND2_X1 U1461 ( .A1(n9157), .A2(n4745), .ZN(n4961) );
  NAND2_X1 U1462 ( .A1(n4963), .A2(n4962), .ZN(n8591) );
  NAND2_X1 U1463 ( .A1(wdata_a_i[19]), .A2(n7690), .ZN(n4962) );
  NAND2_X1 U1464 ( .A1(n8877), .A2(n3851), .ZN(n4963) );
  NAND2_X1 U1465 ( .A1(n4965), .A2(n4964), .ZN(n8796) );
  NAND2_X1 U1466 ( .A1(wdata_a_i[23]), .A2(n7831), .ZN(n4964) );
  NAND2_X1 U1467 ( .A1(n4775), .A2(n4821), .ZN(n4965) );
  NAND2_X1 U1468 ( .A1(n4967), .A2(n4966), .ZN(n8924) );
  NAND2_X1 U1469 ( .A1(wdata_a_i[23]), .A2(n7901), .ZN(n4966) );
  NAND2_X1 U1470 ( .A1(n4797), .A2(n4823), .ZN(n4967) );
  NAND2_X1 U1471 ( .A1(n4969), .A2(n4968), .ZN(n8959) );
  NAND2_X1 U1472 ( .A1(wdata_a_i[23]), .A2(n7915), .ZN(n4968) );
  NAND2_X1 U1473 ( .A1(n9157), .A2(n4814), .ZN(n4969) );
  NAND2_X1 U1474 ( .A1(n4971), .A2(n4970), .ZN(n8994) );
  NAND2_X1 U1475 ( .A1(wdata_a_i[23]), .A2(n7946), .ZN(n4970) );
  NAND2_X1 U1476 ( .A1(n4973), .A2(n4972), .ZN(n9029) );
  NAND2_X1 U1477 ( .A1(wdata_a_i[23]), .A2(n7960), .ZN(n4972) );
  NAND2_X1 U1478 ( .A1(n9157), .A2(n4813), .ZN(n4973) );
  NAND2_X1 U1479 ( .A1(n4975), .A2(n4974), .ZN(n8416) );
  NAND2_X1 U1481 ( .A1(wdata_a_i[19]), .A2(n7573), .ZN(n4974) );
  NAND2_X1 U1482 ( .A1(n9074), .A2(n4745), .ZN(n4975) );
  NAND2_X1 U1483 ( .A1(n4977), .A2(n4976), .ZN(n8460) );
  NAND2_X1 U1484 ( .A1(wdata_a_i[10]), .A2(n7592), .ZN(n4976) );
  NAND2_X1 U1485 ( .A1(n8894), .A2(n4810), .ZN(n4977) );
  NAND2_X1 U1507 ( .A1(n4979), .A2(n4978), .ZN(n8495) );
  NAND2_X1 U1508 ( .A1(wdata_a_i[10]), .A2(n7615), .ZN(n4978) );
  NAND2_X1 U1509 ( .A1(n8894), .A2(n4808), .ZN(n4979) );
  NAND2_X1 U1510 ( .A1(n4981), .A2(n4980), .ZN(n8530) );
  NAND2_X1 U1511 ( .A1(wdata_a_i[10]), .A2(n7639), .ZN(n4980) );
  NAND2_X1 U1512 ( .A1(n8894), .A2(n4811), .ZN(n4981) );
  NAND2_X1 U1513 ( .A1(n4983), .A2(n4982), .ZN(n8565) );
  NAND2_X1 U1514 ( .A1(wdata_a_i[10]), .A2(n7662), .ZN(n4982) );
  NAND2_X1 U1515 ( .A1(n8894), .A2(n4809), .ZN(n4983) );
  NAND2_X1 U1516 ( .A1(n4985), .A2(n4984), .ZN(n8800) );
  NAND2_X1 U1517 ( .A1(wdata_a_i[19]), .A2(n7833), .ZN(n4984) );
  NAND2_X1 U1518 ( .A1(n9074), .A2(n4821), .ZN(n4985) );
  NAND2_X1 U1519 ( .A1(n4987), .A2(n4986), .ZN(n8928) );
  NAND2_X1 U1520 ( .A1(wdata_a_i[19]), .A2(n7903), .ZN(n4986) );
  NAND2_X1 U1521 ( .A1(n9074), .A2(n4823), .ZN(n4987) );
  NAND2_X1 U1522 ( .A1(n4989), .A2(n4988), .ZN(n8963) );
  NAND2_X1 U1523 ( .A1(wdata_a_i[19]), .A2(n7916), .ZN(n4988) );
  NAND2_X1 U1524 ( .A1(n9164), .A2(n4814), .ZN(n4989) );
  NAND2_X1 U1525 ( .A1(n4991), .A2(n4990), .ZN(n8998) );
  NAND2_X1 U1526 ( .A1(wdata_a_i[19]), .A2(n7948), .ZN(n4990) );
  NAND2_X1 U1527 ( .A1(n4993), .A2(n4992), .ZN(n9034) );
  NAND2_X1 U1528 ( .A1(wdata_a_i[19]), .A2(n7962), .ZN(n4992) );
  NAND2_X1 U1529 ( .A1(n8877), .A2(n4813), .ZN(n4993) );
  NAND2_X1 U1530 ( .A1(n4995), .A2(n4994), .ZN(n8704) );
  NAND2_X1 U1531 ( .A1(wdata_a_i[10]), .A2(n7757), .ZN(n4994) );
  NAND2_X1 U1532 ( .A1(n8894), .A2(n1617), .ZN(n4995) );
  NAND2_X1 U1533 ( .A1(n4997), .A2(n4996), .ZN(n8774) );
  NAND2_X1 U1534 ( .A1(wdata_a_i[10]), .A2(n7806), .ZN(n4996) );
  NAND2_X1 U1535 ( .A1(n8894), .A2(n1640), .ZN(n4997) );
  NAND2_X1 U1536 ( .A1(n4999), .A2(n4998), .ZN(n8093) );
  NAND2_X1 U1537 ( .A1(n4459), .A2(n7388), .ZN(n4998) );
  NAND2_X1 U1538 ( .A1(n8867), .A2(n4822), .ZN(n4999) );
  NAND2_X1 U1539 ( .A1(n5001), .A2(n5000), .ZN(n8163) );
  NAND2_X1 U1540 ( .A1(n4459), .A2(n7432), .ZN(n5000) );
  NAND2_X1 U1541 ( .A1(n9152), .A2(n4820), .ZN(n5001) );
  INV_X2 U1542 ( .A(n4380), .ZN(n9162) );
  NAND2_X1 U1543 ( .A1(n5003), .A2(n5002), .ZN(n8405) );
  NAND2_X1 U1544 ( .A1(wdata_a_i[30]), .A2(n7562), .ZN(n5002) );
  NAND2_X1 U1545 ( .A1(n8861), .A2(n4745), .ZN(n5003) );
  NAND2_X1 U1589 ( .A1(n5005), .A2(n5004), .ZN(n8789) );
  NAND2_X1 U1590 ( .A1(wdata_a_i[30]), .A2(n7822), .ZN(n5004) );
  NAND2_X1 U1591 ( .A1(n4731), .A2(n4821), .ZN(n5005) );
  NAND2_X1 U1592 ( .A1(n5007), .A2(n5006), .ZN(n8952) );
  NAND2_X1 U1593 ( .A1(wdata_a_i[30]), .A2(n7914), .ZN(n5006) );
  NAND2_X1 U1718 ( .A1(n4731), .A2(n4814), .ZN(n5007) );
  NAND2_X1 U1719 ( .A1(n5009), .A2(n5008), .ZN(n8987) );
  NAND2_X1 U1720 ( .A1(wdata_a_i[30]), .A2(n7937), .ZN(n5008) );
  NAND2_X1 U1721 ( .A1(n4731), .A2(n4826), .ZN(n5009) );
  NAND2_X1 U1722 ( .A1(n5011), .A2(n5010), .ZN(n9022) );
  NAND2_X1 U1766 ( .A1(wdata_a_i[30]), .A2(n7960), .ZN(n5010) );
  NAND2_X1 U1767 ( .A1(n4731), .A2(n4813), .ZN(n5011) );
  NAND2_X1 U1768 ( .A1(n5013), .A2(n5012), .ZN(n8916) );
  NAND2_X1 U1769 ( .A1(n4623), .A2(n7893), .ZN(n5012) );
  NAND2_X1 U1770 ( .A1(n9146), .A2(n4823), .ZN(n5013) );
  NAND2_X1 U1771 ( .A1(n5015), .A2(n5014), .ZN(n8588) );
  NAND2_X1 U1774 ( .A1(wdata_a_i[22]), .A2(n7688), .ZN(n5014) );
  NAND2_X1 U1776 ( .A1(n4737), .A2(n3851), .ZN(n5015) );
  NAND2_X1 U1777 ( .A1(n5017), .A2(n5016), .ZN(n8622) );
  NAND2_X1 U1778 ( .A1(wdata_a_i[22]), .A2(n7711), .ZN(n5016) );
  NAND2_X1 U1779 ( .A1(n4788), .A2(n1647), .ZN(n5017) );
  NAND2_X1 U1781 ( .A1(n5019), .A2(n5018), .ZN(n8657) );
  NAND2_X1 U1782 ( .A1(wdata_a_i[22]), .A2(n7735), .ZN(n5018) );
  NAND2_X1 U1783 ( .A1(n4737), .A2(n3774), .ZN(n5019) );
  NAND2_X1 U1784 ( .A1(n5021), .A2(n5020), .ZN(n8692) );
  NAND2_X1 U1785 ( .A1(wdata_a_i[22]), .A2(n7750), .ZN(n5020) );
  NAND2_X1 U1786 ( .A1(n4737), .A2(n1617), .ZN(n5021) );
  NAND2_X1 U1787 ( .A1(n5023), .A2(n5022), .ZN(n8762) );
  NAND2_X1 U1788 ( .A1(wdata_a_i[22]), .A2(n7799), .ZN(n5022) );
  NAND2_X1 U1789 ( .A1(n4788), .A2(n1640), .ZN(n5023) );
  NAND2_X1 U1790 ( .A1(n5025), .A2(n5024), .ZN(n8832) );
  NAND2_X1 U1791 ( .A1(wdata_a_i[22]), .A2(n7854), .ZN(n5024) );
  NAND2_X1 U1792 ( .A1(n4737), .A2(n1629), .ZN(n5025) );
  NAND2_X1 U1793 ( .A1(n5027), .A2(n5026), .ZN(n8342) );
  NAND2_X1 U1794 ( .A1(wdata_a_i[22]), .A2(n7518), .ZN(n5026) );
  NAND2_X1 U1795 ( .A1(n9068), .A2(n4817), .ZN(n5027) );
  NAND2_X1 U1796 ( .A1(n5029), .A2(n5028), .ZN(n8413) );
  NAND2_X1 U1797 ( .A1(wdata_a_i[22]), .A2(n7571), .ZN(n5028) );
  NAND2_X1 U1798 ( .A1(n9068), .A2(n4745), .ZN(n5029) );
  NAND2_X1 U1799 ( .A1(n5031), .A2(n5030), .ZN(n8797) );
  NAND2_X1 U1800 ( .A1(wdata_a_i[22]), .A2(n7831), .ZN(n5030) );
  NAND2_X1 U1801 ( .A1(n9068), .A2(n4821), .ZN(n5031) );
  NAND2_X1 U1802 ( .A1(n5033), .A2(n5032), .ZN(n8925) );
  NAND2_X1 U1803 ( .A1(wdata_a_i[22]), .A2(n7901), .ZN(n5032) );
  NAND2_X1 U1804 ( .A1(n9068), .A2(n4823), .ZN(n5033) );
  NAND2_X1 U1805 ( .A1(n5035), .A2(n5034), .ZN(n8960) );
  NAND2_X1 U1806 ( .A1(wdata_a_i[22]), .A2(n7915), .ZN(n5034) );
  NAND2_X1 U1807 ( .A1(n9068), .A2(n4814), .ZN(n5035) );
  NAND2_X1 U1808 ( .A1(n5037), .A2(n5036), .ZN(n8995) );
  NAND2_X1 U1809 ( .A1(wdata_a_i[22]), .A2(n7946), .ZN(n5036) );
  NAND2_X1 U1810 ( .A1(n9159), .A2(n4826), .ZN(n5037) );
  NAND2_X1 U1811 ( .A1(n5039), .A2(n5038), .ZN(n9030) );
  NAND2_X1 U1812 ( .A1(wdata_a_i[22]), .A2(n7962), .ZN(n5038) );
  NAND2_X1 U1982 ( .A1(n9068), .A2(n4813), .ZN(n5039) );
  NAND2_X1 U1983 ( .A1(n5041), .A2(n5040), .ZN(n8418) );
  NAND2_X1 U1984 ( .A1(wdata_a_i[17]), .A2(n7575), .ZN(n5040) );
  NAND2_X1 U1985 ( .A1(n9078), .A2(n4745), .ZN(n5041) );
  NAND2_X1 U1986 ( .A1(n5043), .A2(n5042), .ZN(n8802) );
  NAND2_X1 U1987 ( .A1(wdata_a_i[17]), .A2(n7835), .ZN(n5042) );
  NAND2_X1 U1988 ( .A1(n9078), .A2(n4821), .ZN(n5043) );
  NAND2_X1 U1989 ( .A1(n5045), .A2(n5044), .ZN(n8930) );
  NAND2_X1 U1990 ( .A1(wdata_a_i[17]), .A2(n7905), .ZN(n5044) );
  NAND2_X1 U1991 ( .A1(n9078), .A2(n4823), .ZN(n5045) );
  NAND2_X1 U1992 ( .A1(n5047), .A2(n5046), .ZN(n8965) );
  NAND2_X1 U1993 ( .A1(wdata_a_i[17]), .A2(n7917), .ZN(n5046) );
  NAND2_X1 U1994 ( .A1(n4805), .A2(n4814), .ZN(n5047) );
  NAND2_X1 U1995 ( .A1(n5049), .A2(n5048), .ZN(n9000) );
  NAND2_X1 U1996 ( .A1(wdata_a_i[17]), .A2(n7950), .ZN(n5048) );
  NAND2_X1 U1997 ( .A1(n5051), .A2(n5050), .ZN(n9036) );
  NAND2_X1 U1998 ( .A1(wdata_a_i[17]), .A2(n7963), .ZN(n5050) );
  NAND2_X1 U1999 ( .A1(n4806), .A2(n4813), .ZN(n5051) );
  NAND2_X1 U2000 ( .A1(n5053), .A2(n5052), .ZN(n8593) );
  NAND2_X1 U2001 ( .A1(wdata_a_i[17]), .A2(n7692), .ZN(n5052) );
  NAND2_X1 U2002 ( .A1(n8881), .A2(n3851), .ZN(n5053) );
  NAND2_X1 U2003 ( .A1(n5055), .A2(n5054), .ZN(n8579) );
  NAND2_X1 U2004 ( .A1(n4477), .A2(n7678), .ZN(n5054) );
  NAND2_X1 U2005 ( .A1(n4789), .A2(n3851), .ZN(n5055) );
  NAND2_X1 U2006 ( .A1(n5057), .A2(n5056), .ZN(n8614) );
  NAND2_X1 U2007 ( .A1(n4477), .A2(n7702), .ZN(n5056) );
  NAND2_X1 U2008 ( .A1(n4789), .A2(n1647), .ZN(n5057) );
  NAND2_X1 U2009 ( .A1(n5059), .A2(n5058), .ZN(n8648) );
  NAND2_X1 U2010 ( .A1(n4477), .A2(n7725), .ZN(n5058) );
  NAND2_X1 U2011 ( .A1(n4789), .A2(n3774), .ZN(n5059) );
  NAND2_X1 U2012 ( .A1(n5061), .A2(n5060), .ZN(n8683) );
  NAND2_X1 U2013 ( .A1(n4477), .A2(n7749), .ZN(n5060) );
  NAND2_X1 U2014 ( .A1(n4789), .A2(n1617), .ZN(n5061) );
  NAND2_X1 U2015 ( .A1(n5063), .A2(n5062), .ZN(n8718) );
  NAND2_X1 U2016 ( .A1(n4477), .A2(n7773), .ZN(n5062) );
  NAND2_X1 U2017 ( .A1(n4789), .A2(n1634), .ZN(n5063) );
  NAND2_X1 U2018 ( .A1(n5065), .A2(n5064), .ZN(n8753) );
  NAND2_X1 U2019 ( .A1(n4477), .A2(n7798), .ZN(n5064) );
  NAND2_X1 U2020 ( .A1(n4789), .A2(n1640), .ZN(n5065) );
  NAND2_X1 U2021 ( .A1(n5067), .A2(n5066), .ZN(n8823) );
  NAND2_X1 U2022 ( .A1(n4477), .A2(n7844), .ZN(n5066) );
  NAND2_X1 U2023 ( .A1(n4789), .A2(n1629), .ZN(n5067) );
  INV_X2 U2024 ( .A(n4380), .ZN(n8875) );
  NAND2_X1 U2025 ( .A1(n5069), .A2(n5068), .ZN(n8649) );
  NAND2_X1 U2026 ( .A1(n4623), .A2(n7725), .ZN(n5068) );
  NAND2_X1 U2027 ( .A1(n8861), .A2(n3774), .ZN(n5069) );
  NAND2_X1 U2028 ( .A1(n5071), .A2(n5070), .ZN(n8719) );
  NAND2_X1 U2029 ( .A1(n4623), .A2(n7773), .ZN(n5070) );
  NAND2_X1 U2030 ( .A1(n8861), .A2(n1634), .ZN(n5071) );
  NAND2_X1 U2031 ( .A1(n5073), .A2(n5072), .ZN(n8824) );
  NAND2_X1 U2032 ( .A1(n4623), .A2(n7844), .ZN(n5072) );
  NAND2_X1 U2033 ( .A1(n8861), .A2(n1629), .ZN(n5073) );
  NAND2_X1 U2034 ( .A1(n5075), .A2(n5074), .ZN(n8062) );
  NAND2_X1 U2036 ( .A1(wdata_a_i[22]), .A2(n7363), .ZN(n5074) );
  NAND2_X1 U2039 ( .A1(n9159), .A2(n4816), .ZN(n5075) );
  NAND2_X1 U2040 ( .A1(n5077), .A2(n5076), .ZN(n8097) );
  NAND2_X1 U2041 ( .A1(wdata_a_i[22]), .A2(n7392), .ZN(n5076) );
  NAND2_X1 U2042 ( .A1(n9159), .A2(n4822), .ZN(n5077) );
  NAND2_X1 U2043 ( .A1(n5079), .A2(n5078), .ZN(n8132) );
  NAND2_X1 U2044 ( .A1(wdata_a_i[22]), .A2(n7406), .ZN(n5078) );
  NAND2_X1 U2046 ( .A1(n9159), .A2(n4815), .ZN(n5079) );
  NAND2_X1 U2047 ( .A1(n5081), .A2(n5080), .ZN(n8167) );
  NAND2_X1 U2048 ( .A1(wdata_a_i[22]), .A2(n7436), .ZN(n5080) );
  NAND2_X1 U2049 ( .A1(n9068), .A2(n4820), .ZN(n5081) );
  NAND2_X1 U2050 ( .A1(n5083), .A2(n5082), .ZN(n8202) );
  NAND2_X1 U2052 ( .A1(wdata_a_i[22]), .A2(n7450), .ZN(n5082) );
  NAND2_X1 U2055 ( .A1(n9159), .A2(n4812), .ZN(n5083) );
  NAND2_X1 U2056 ( .A1(n5085), .A2(n5084), .ZN(n8272) );
  NAND2_X1 U2057 ( .A1(wdata_a_i[22]), .A2(n7473), .ZN(n5084) );
  NAND2_X1 U2058 ( .A1(n9159), .A2(n4819), .ZN(n5085) );
  NAND2_X1 U2059 ( .A1(n5087), .A2(n5086), .ZN(n8307) );
  NAND2_X1 U2102 ( .A1(wdata_a_i[22]), .A2(n7495), .ZN(n5086) );
  NAND2_X1 U2106 ( .A1(n9159), .A2(n4746), .ZN(n5087) );
  NAND2_X1 U2107 ( .A1(n5089), .A2(n5088), .ZN(n8378) );
  NAND2_X1 U2108 ( .A1(wdata_a_i[22]), .A2(n7540), .ZN(n5088) );
  NAND2_X1 U2109 ( .A1(n9159), .A2(n4807), .ZN(n5089) );
  NAND2_X1 U2110 ( .A1(n5091), .A2(n5090), .ZN(n9118) );
  NAND2_X1 U2113 ( .A1(wdata_a_i[22]), .A2(n8009), .ZN(n5090) );
  NAND2_X1 U2114 ( .A1(n9159), .A2(n4818), .ZN(n5091) );
  NAND2_X1 U2115 ( .A1(n5093), .A2(n5092), .ZN(n8054) );
  NAND2_X1 U2116 ( .A1(n4472), .A2(n7362), .ZN(n5092) );
  NAND2_X1 U2117 ( .A1(n9146), .A2(n4816), .ZN(n5093) );
  NAND2_X1 U2118 ( .A1(n5095), .A2(n5094), .ZN(n8089) );
  NAND2_X1 U2120 ( .A1(n4472), .A2(n7384), .ZN(n5094) );
  NAND2_X1 U2121 ( .A1(n9146), .A2(n4822), .ZN(n5095) );
  NAND2_X1 U2122 ( .A1(n5097), .A2(n5096), .ZN(n8124) );
  NAND2_X1 U2123 ( .A1(n4472), .A2(n7405), .ZN(n5096) );
  NAND2_X1 U2124 ( .A1(n9146), .A2(n4815), .ZN(n5097) );
  NAND2_X1 U2125 ( .A1(n5099), .A2(n5098), .ZN(n8159) );
  NAND2_X1 U2128 ( .A1(n4472), .A2(n7427), .ZN(n5098) );
  NAND2_X1 U2129 ( .A1(n9146), .A2(n4820), .ZN(n5099) );
  NAND2_X1 U2130 ( .A1(n5101), .A2(n5100), .ZN(n8194) );
  NAND2_X1 U2131 ( .A1(n4472), .A2(n7449), .ZN(n5100) );
  NAND2_X1 U2468 ( .A1(n9146), .A2(n4812), .ZN(n5101) );
  NAND2_X1 U2473 ( .A1(n5103), .A2(n5102), .ZN(n8264) );
  NAND2_X1 U2478 ( .A1(n4472), .A2(n7472), .ZN(n5102) );
  NAND2_X1 U2483 ( .A1(n9146), .A2(n4819), .ZN(n5103) );
  NAND2_X1 U2484 ( .A1(n5105), .A2(n5104), .ZN(n8299) );
  NAND2_X1 U2485 ( .A1(n4472), .A2(n7494), .ZN(n5104) );
  NAND2_X1 U2486 ( .A1(n9146), .A2(n4746), .ZN(n5105) );
  NAND2_X1 U2487 ( .A1(n5107), .A2(n5106), .ZN(n8334) );
  NAND2_X1 U2488 ( .A1(n4472), .A2(n7517), .ZN(n5106) );
  NAND2_X1 U2489 ( .A1(n9146), .A2(n4817), .ZN(n5107) );
  NAND2_X1 U2490 ( .A1(n5109), .A2(n5108), .ZN(n8370) );
  NAND2_X1 U2491 ( .A1(n4472), .A2(n7539), .ZN(n5108) );
  NAND2_X1 U2492 ( .A1(n9146), .A2(n4807), .ZN(n5109) );
  NAND2_X1 U2493 ( .A1(n5111), .A2(n5110), .ZN(n8580) );
  NAND2_X1 U2494 ( .A1(n4623), .A2(n7678), .ZN(n5110) );
  NAND2_X1 U2495 ( .A1(n8861), .A2(n3851), .ZN(n5111) );
  NAND2_X1 U2496 ( .A1(n5113), .A2(n5112), .ZN(n8615) );
  NAND2_X1 U2497 ( .A1(n4623), .A2(n7702), .ZN(n5112) );
  NAND2_X1 U2498 ( .A1(n8861), .A2(n1647), .ZN(n5113) );
  NAND2_X1 U2499 ( .A1(n5115), .A2(n5114), .ZN(n8684) );
  NAND2_X1 U2500 ( .A1(n4623), .A2(n7749), .ZN(n5114) );
  NAND2_X1 U2501 ( .A1(n8861), .A2(n1617), .ZN(n5115) );
  NAND2_X1 U2502 ( .A1(n5117), .A2(n5116), .ZN(n8754) );
  NAND2_X1 U2503 ( .A1(n4623), .A2(n7798), .ZN(n5116) );
  NAND2_X1 U2504 ( .A1(n8861), .A2(n1640), .ZN(n5117) );
  NAND2_X1 U2505 ( .A1(n5119), .A2(n5118), .ZN(n9110) );
  NAND2_X1 U2506 ( .A1(n4472), .A2(n8008), .ZN(n5118) );
  NAND2_X1 U2507 ( .A1(n9146), .A2(n4818), .ZN(n5119) );
  NAND2_X1 U2508 ( .A1(n5121), .A2(n5120), .ZN(n8625) );
  NAND2_X1 U2509 ( .A1(wdata_a_i[19]), .A2(n7713), .ZN(n5120) );
  NAND2_X1 U2510 ( .A1(n8877), .A2(n1647), .ZN(n5121) );
  NAND2_X1 U2511 ( .A1(n5123), .A2(n5122), .ZN(n8660) );
  NAND2_X1 U2512 ( .A1(wdata_a_i[19]), .A2(n7737), .ZN(n5122) );
  NAND2_X1 U2513 ( .A1(n9074), .A2(n3774), .ZN(n5123) );
  NAND2_X1 U2514 ( .A1(n5125), .A2(n5124), .ZN(n8695) );
  NAND2_X1 U2515 ( .A1(wdata_a_i[19]), .A2(n7751), .ZN(n5124) );
  NAND2_X1 U2516 ( .A1(n8877), .A2(n1617), .ZN(n5125) );
  NAND2_X1 U2517 ( .A1(n5127), .A2(n5126), .ZN(n8730) );
  NAND2_X1 U2518 ( .A1(wdata_a_i[19]), .A2(n7785), .ZN(n5126) );
  NAND2_X1 U2519 ( .A1(n8877), .A2(n1634), .ZN(n5127) );
  NAND2_X1 U2520 ( .A1(n5129), .A2(n5128), .ZN(n8765) );
  NAND2_X1 U2521 ( .A1(wdata_a_i[19]), .A2(n7800), .ZN(n5128) );
  NAND2_X1 U2522 ( .A1(n8877), .A2(n1640), .ZN(n5129) );
  NAND2_X1 U2523 ( .A1(n5131), .A2(n5130), .ZN(n8835) );
  NAND2_X1 U2524 ( .A1(wdata_a_i[19]), .A2(n7856), .ZN(n5130) );
  NAND2_X1 U2525 ( .A1(n8877), .A2(n1629), .ZN(n5131) );
  NAND2_X1 U2526 ( .A1(n5133), .A2(n5132), .ZN(n8587) );
  NAND2_X1 U2527 ( .A1(wdata_a_i[23]), .A2(n7688), .ZN(n5132) );
  NAND2_X1 U3116 ( .A1(n8871), .A2(n3851), .ZN(n5133) );
  NAND2_X1 U3117 ( .A1(n5135), .A2(n5134), .ZN(n8590) );
  NAND2_X1 U3118 ( .A1(wdata_a_i[20]), .A2(n7689), .ZN(n5134) );
  NAND2_X1 U3119 ( .A1(n8875), .A2(n3851), .ZN(n5135) );
  NAND2_X1 U3120 ( .A1(n5137), .A2(n5136), .ZN(n8621) );
  NAND2_X1 U3121 ( .A1(wdata_a_i[23]), .A2(n7711), .ZN(n5136) );
  NAND2_X1 U3122 ( .A1(n5139), .A2(n5138), .ZN(n8624) );
  NAND2_X1 U3123 ( .A1(wdata_a_i[20]), .A2(n7712), .ZN(n5138) );
  NAND2_X1 U3126 ( .A1(n8875), .A2(n1647), .ZN(n5139) );
  NAND2_X1 U3127 ( .A1(n5141), .A2(n5140), .ZN(n8627) );
  NAND2_X1 U3128 ( .A1(wdata_a_i[17]), .A2(n7715), .ZN(n5140) );
  NAND2_X1 U3129 ( .A1(n8881), .A2(n1647), .ZN(n5141) );
  NAND2_X1 U3130 ( .A1(n5143), .A2(n5142), .ZN(n8656) );
  NAND2_X1 U3131 ( .A1(wdata_a_i[23]), .A2(n7735), .ZN(n5142) );
  NAND2_X1 U3132 ( .A1(n5145), .A2(n5144), .ZN(n8659) );
  NAND2_X1 U3133 ( .A1(wdata_a_i[20]), .A2(n7736), .ZN(n5144) );
  NAND2_X1 U3134 ( .A1(n9072), .A2(n3774), .ZN(n5145) );
  NAND2_X1 U3135 ( .A1(n5147), .A2(n5146), .ZN(n8662) );
  NAND2_X1 U3136 ( .A1(wdata_a_i[17]), .A2(n7739), .ZN(n5146) );
  NAND2_X1 U3137 ( .A1(n8881), .A2(n3774), .ZN(n5147) );
  NAND2_X1 U3138 ( .A1(n5149), .A2(n5148), .ZN(n8691) );
  NAND2_X1 U3139 ( .A1(wdata_a_i[23]), .A2(n7750), .ZN(n5148) );
  NAND2_X1 U3140 ( .A1(n8871), .A2(n1617), .ZN(n5149) );
  NAND2_X1 U3142 ( .A1(n5151), .A2(n5150), .ZN(n8694) );
  NAND2_X1 U3143 ( .A1(wdata_a_i[20]), .A2(n7751), .ZN(n5150) );
  NAND2_X1 U3145 ( .A1(n8875), .A2(n1617), .ZN(n5151) );
  NAND2_X1 U3146 ( .A1(n5153), .A2(n5152), .ZN(n8697) );
  NAND2_X1 U3148 ( .A1(wdata_a_i[17]), .A2(n7752), .ZN(n5152) );
  NAND2_X1 U3149 ( .A1(n8881), .A2(n1617), .ZN(n5153) );
  NAND2_X1 U3151 ( .A1(n5155), .A2(n5154), .ZN(n8726) );
  NAND2_X1 U3152 ( .A1(wdata_a_i[23]), .A2(n7783), .ZN(n5154) );
  NAND2_X1 U3154 ( .A1(n8871), .A2(n1634), .ZN(n5155) );
  NAND2_X1 U3155 ( .A1(n5157), .A2(n5156), .ZN(n8729) );
  NAND2_X1 U3157 ( .A1(wdata_a_i[20]), .A2(n7784), .ZN(n5156) );
  NAND2_X1 U3158 ( .A1(n8875), .A2(n1634), .ZN(n5157) );
  NAND2_X1 U3160 ( .A1(n5159), .A2(n5158), .ZN(n8732) );
  NAND2_X1 U3161 ( .A1(wdata_a_i[17]), .A2(n7787), .ZN(n5158) );
  NAND2_X1 U3163 ( .A1(n8881), .A2(n1634), .ZN(n5159) );
  NAND2_X1 U3164 ( .A1(n5161), .A2(n5160), .ZN(n8761) );
  NAND2_X1 U3165 ( .A1(wdata_a_i[23]), .A2(n7799), .ZN(n5160) );
  NAND2_X1 U3167 ( .A1(n8871), .A2(n1640), .ZN(n5161) );
  NAND2_X1 U3168 ( .A1(n5163), .A2(n5162), .ZN(n8764) );
  NAND2_X1 U3169 ( .A1(wdata_a_i[20]), .A2(n7800), .ZN(n5162) );
  NAND2_X1 U3170 ( .A1(n5165), .A2(n5164), .ZN(n8767) );
  NAND2_X1 U3171 ( .A1(wdata_a_i[17]), .A2(n7801), .ZN(n5164) );
  NAND2_X1 U3172 ( .A1(n8881), .A2(n1640), .ZN(n5165) );
  NAND2_X1 U3173 ( .A1(n5167), .A2(n5166), .ZN(n8831) );
  NAND2_X1 U3175 ( .A1(wdata_a_i[23]), .A2(n7854), .ZN(n5166) );
  NAND2_X1 U3176 ( .A1(n8871), .A2(n1629), .ZN(n5167) );
  NAND2_X1 U3178 ( .A1(n5169), .A2(n5168), .ZN(n8834) );
  NAND2_X1 U3179 ( .A1(wdata_a_i[20]), .A2(n7855), .ZN(n5168) );
  NAND2_X1 U3180 ( .A1(n8875), .A2(n1629), .ZN(n5169) );
  NAND2_X1 U3181 ( .A1(n5171), .A2(n5170), .ZN(n8837) );
  NAND2_X1 U3182 ( .A1(wdata_a_i[17]), .A2(n7858), .ZN(n5170) );
  NAND2_X1 U3183 ( .A1(n8881), .A2(n1629), .ZN(n5171) );
  NAND2_X1 U3184 ( .A1(n5173), .A2(n5172), .ZN(n8592) );
  NAND2_X1 U3186 ( .A1(wdata_a_i[18]), .A2(n7690), .ZN(n5172) );
  NAND2_X1 U3187 ( .A1(n5175), .A2(n5174), .ZN(n8626) );
  NAND2_X1 U3188 ( .A1(wdata_a_i[18]), .A2(n7713), .ZN(n5174) );
  NAND2_X1 U3189 ( .A1(n4792), .A2(n1647), .ZN(n5175) );
  NAND2_X1 U3190 ( .A1(n5177), .A2(n5176), .ZN(n8661) );
  NAND2_X1 U3191 ( .A1(wdata_a_i[18]), .A2(n7737), .ZN(n5176) );
  NAND2_X1 U3192 ( .A1(n9166), .A2(n3774), .ZN(n5177) );
  NAND2_X1 U3193 ( .A1(n5179), .A2(n5178), .ZN(n8696) );
  NAND2_X1 U3194 ( .A1(wdata_a_i[18]), .A2(n7752), .ZN(n5178) );
  NAND2_X1 U3195 ( .A1(n4792), .A2(n1617), .ZN(n5179) );
  NAND2_X1 U3196 ( .A1(n5181), .A2(n5180), .ZN(n8731) );
  NAND2_X1 U3197 ( .A1(wdata_a_i[18]), .A2(n7785), .ZN(n5180) );
  NAND2_X1 U3198 ( .A1(n5183), .A2(n5182), .ZN(n8766) );
  NAND2_X1 U3199 ( .A1(wdata_a_i[18]), .A2(n7801), .ZN(n5182) );
  NAND2_X1 U3200 ( .A1(n4792), .A2(n1640), .ZN(n5183) );
  NAND2_X1 U3201 ( .A1(n5185), .A2(n5184), .ZN(n8836) );
  NAND2_X1 U3202 ( .A1(wdata_a_i[18]), .A2(n7856), .ZN(n5184) );
  NAND2_X1 U3203 ( .A1(n4793), .A2(n1629), .ZN(n5185) );
  NAND2_X1 U3204 ( .A1(n5187), .A2(n5186), .ZN(n8193) );
  NAND2_X1 U3205 ( .A1(n4477), .A2(n7449), .ZN(n5186) );
  NAND2_X1 U3206 ( .A1(n4784), .A2(n4812), .ZN(n5187) );
  NAND2_X1 U3207 ( .A1(n5189), .A2(n5188), .ZN(n8263) );
  NAND2_X1 U3208 ( .A1(n4477), .A2(n7472), .ZN(n5188) );
  NAND2_X1 U3209 ( .A1(n4789), .A2(n4819), .ZN(n5189) );
  NAND2_X1 U3210 ( .A1(n5191), .A2(n5190), .ZN(n8439) );
  NAND2_X1 U3211 ( .A1(n4477), .A2(n7584), .ZN(n5190) );
  NAND2_X1 U3212 ( .A1(n4789), .A2(n4810), .ZN(n5191) );
  NAND2_X1 U3213 ( .A1(n5193), .A2(n5192), .ZN(n8474) );
  NAND2_X1 U3214 ( .A1(n4477), .A2(n7608), .ZN(n5192) );
  NAND2_X1 U3215 ( .A1(n4789), .A2(n4808), .ZN(n5193) );
  NAND2_X1 U3216 ( .A1(n5195), .A2(n5194), .ZN(n8509) );
  NAND2_X1 U3217 ( .A1(n4477), .A2(n7631), .ZN(n5194) );
  NAND2_X1 U3218 ( .A1(n4789), .A2(n4811), .ZN(n5195) );
  NAND2_X1 U3219 ( .A1(n5197), .A2(n5196), .ZN(n8544) );
  NAND2_X1 U3220 ( .A1(n4477), .A2(n7655), .ZN(n5196) );
  NAND2_X1 U3221 ( .A1(n4789), .A2(n4809), .ZN(n5197) );
  NAND2_X1 U3222 ( .A1(n5199), .A2(n5198), .ZN(n8589) );
  NAND2_X1 U3223 ( .A1(wdata_a_i[21]), .A2(n7689), .ZN(n5198) );
  NAND2_X1 U3224 ( .A1(n9032), .A2(n3851), .ZN(n5199) );
  NAND2_X1 U3225 ( .A1(n5201), .A2(n5200), .ZN(n8658) );
  NAND2_X1 U3226 ( .A1(wdata_a_i[21]), .A2(n7736), .ZN(n5200) );
  NAND2_X1 U3227 ( .A1(n9032), .A2(n3774), .ZN(n5201) );
  NAND2_X1 U3228 ( .A1(n5203), .A2(n5202), .ZN(n8098) );
  NAND2_X1 U3229 ( .A1(wdata_a_i[21]), .A2(n7393), .ZN(n5202) );
  NAND2_X1 U3230 ( .A1(n9070), .A2(n4822), .ZN(n5203) );
  NAND2_X1 U3231 ( .A1(n5205), .A2(n5204), .ZN(n8133) );
  NAND2_X1 U3232 ( .A1(wdata_a_i[21]), .A2(n7407), .ZN(n5204) );
  NAND2_X1 U3233 ( .A1(n9070), .A2(n4815), .ZN(n5205) );
  NAND2_X1 U3234 ( .A1(n5207), .A2(n5206), .ZN(n8168) );
  NAND2_X1 U3235 ( .A1(wdata_a_i[21]), .A2(n7437), .ZN(n5206) );
  NAND2_X1 U3236 ( .A1(n9070), .A2(n4820), .ZN(n5207) );
  NAND2_X1 U3237 ( .A1(n5209), .A2(n5208), .ZN(n8203) );
  NAND2_X1 U3238 ( .A1(wdata_a_i[21]), .A2(n7451), .ZN(n5208) );
  NAND2_X1 U3239 ( .A1(wdata_b_i[21]), .A2(n4812), .ZN(n5209) );
  NAND2_X1 U3240 ( .A1(n5211), .A2(n5210), .ZN(n8273) );
  NAND2_X1 U3241 ( .A1(wdata_a_i[21]), .A2(n7474), .ZN(n5210) );
  NAND2_X1 U3242 ( .A1(n9070), .A2(n4819), .ZN(n5211) );
  NAND2_X1 U3243 ( .A1(n5213), .A2(n5212), .ZN(n8343) );
  NAND2_X1 U3244 ( .A1(wdata_a_i[21]), .A2(n7519), .ZN(n5212) );
  NAND2_X1 U3245 ( .A1(wdata_b_i[21]), .A2(n4817), .ZN(n5213) );
  NAND2_X1 U3246 ( .A1(n5215), .A2(n5214), .ZN(n8414) );
  NAND2_X1 U3247 ( .A1(wdata_a_i[21]), .A2(n7572), .ZN(n5214) );
  NAND2_X1 U3248 ( .A1(n9032), .A2(n4745), .ZN(n5215) );
  NAND2_X1 U3249 ( .A1(n5217), .A2(n5216), .ZN(n8554) );
  NAND2_X1 U3250 ( .A1(wdata_a_i[21]), .A2(n7657), .ZN(n5216) );
  NAND2_X1 U3251 ( .A1(wdata_b_i[21]), .A2(n4809), .ZN(n5217) );
  NAND2_X1 U3252 ( .A1(n5219), .A2(n5218), .ZN(n8798) );
  NAND2_X1 U3253 ( .A1(wdata_a_i[21]), .A2(n7832), .ZN(n5218) );
  NAND2_X1 U3254 ( .A1(n9070), .A2(n4821), .ZN(n5219) );
  NAND2_X1 U3255 ( .A1(n5221), .A2(n5220), .ZN(n9119) );
  NAND2_X1 U3256 ( .A1(wdata_a_i[21]), .A2(n8010), .ZN(n5220) );
  NAND2_X1 U3257 ( .A1(n9070), .A2(n4818), .ZN(n5221) );
  NAND2_X1 U3258 ( .A1(n5223), .A2(n5222), .ZN(n8448) );
  NAND2_X1 U3259 ( .A1(wdata_a_i[22]), .A2(n7585), .ZN(n5222) );
  NAND2_X1 U3260 ( .A1(n4737), .A2(n4810), .ZN(n5223) );
  NAND2_X1 U3261 ( .A1(n5225), .A2(n5224), .ZN(n8483) );
  NAND2_X1 U3262 ( .A1(wdata_a_i[22]), .A2(n7609), .ZN(n5224) );
  NAND2_X1 U3263 ( .A1(n4788), .A2(n4808), .ZN(n5225) );
  NAND2_X1 U3264 ( .A1(n5227), .A2(n5226), .ZN(n8518) );
  NAND2_X1 U3265 ( .A1(wdata_a_i[22]), .A2(n7632), .ZN(n5226) );
  NAND2_X1 U3266 ( .A1(n4737), .A2(n4811), .ZN(n5227) );
  NAND2_X1 U3267 ( .A1(n5229), .A2(n5228), .ZN(n8553) );
  NAND2_X1 U3268 ( .A1(wdata_a_i[22]), .A2(n7656), .ZN(n5228) );
  NAND2_X1 U3269 ( .A1(n4788), .A2(n4809), .ZN(n5229) );
  NAND2_X1 U3270 ( .A1(n5231), .A2(n5230), .ZN(n8065) );
  NAND2_X1 U3271 ( .A1(wdata_a_i[19]), .A2(n7365), .ZN(n5230) );
  NAND2_X1 U3272 ( .A1(n9164), .A2(n4816), .ZN(n5231) );
  NAND2_X1 U3273 ( .A1(n5233), .A2(n5232), .ZN(n8135) );
  NAND2_X1 U3274 ( .A1(wdata_a_i[19]), .A2(n7408), .ZN(n5232) );
  NAND2_X1 U3275 ( .A1(n9074), .A2(n4815), .ZN(n5233) );
  NAND2_X1 U3276 ( .A1(n5235), .A2(n5234), .ZN(n8205) );
  NAND2_X1 U3277 ( .A1(wdata_a_i[19]), .A2(n7452), .ZN(n5234) );
  NAND2_X1 U3278 ( .A1(n9074), .A2(n4812), .ZN(n5235) );
  NAND2_X1 U3279 ( .A1(n5237), .A2(n5236), .ZN(n8275) );
  NAND2_X1 U3280 ( .A1(wdata_a_i[19]), .A2(n7475), .ZN(n5236) );
  NAND2_X1 U3281 ( .A1(n9164), .A2(n4819), .ZN(n5237) );
  NAND2_X1 U3282 ( .A1(n5239), .A2(n5238), .ZN(n8310) );
  NAND2_X1 U3283 ( .A1(wdata_a_i[19]), .A2(n7496), .ZN(n5238) );
  NAND2_X1 U3284 ( .A1(n9164), .A2(n4746), .ZN(n5239) );
  NAND2_X1 U3285 ( .A1(n5241), .A2(n5240), .ZN(n8451) );
  NAND2_X1 U3286 ( .A1(wdata_a_i[19]), .A2(n7586), .ZN(n5240) );
  NAND2_X1 U3287 ( .A1(n8877), .A2(n4810), .ZN(n5241) );
  NAND2_X1 U3288 ( .A1(n5243), .A2(n5242), .ZN(n8453) );
  NAND2_X1 U3289 ( .A1(wdata_a_i[17]), .A2(n7587), .ZN(n5242) );
  NAND2_X1 U3290 ( .A1(n8881), .A2(n4810), .ZN(n5243) );
  NAND2_X1 U3291 ( .A1(n5245), .A2(n5244), .ZN(n8486) );
  NAND2_X1 U3292 ( .A1(wdata_a_i[19]), .A2(n7611), .ZN(n5244) );
  NAND2_X1 U3293 ( .A1(n8877), .A2(n4808), .ZN(n5245) );
  NAND2_X1 U3294 ( .A1(n5247), .A2(n5246), .ZN(n8488) );
  NAND2_X1 U3295 ( .A1(wdata_a_i[17]), .A2(n7613), .ZN(n5246) );
  NAND2_X1 U3296 ( .A1(n8881), .A2(n4808), .ZN(n5247) );
  NAND2_X1 U3297 ( .A1(n5249), .A2(n5248), .ZN(n8521) );
  NAND2_X1 U3298 ( .A1(wdata_a_i[19]), .A2(n7633), .ZN(n5248) );
  NAND2_X1 U3299 ( .A1(n8877), .A2(n4811), .ZN(n5249) );
  NAND2_X1 U3300 ( .A1(n5251), .A2(n5250), .ZN(n8523) );
  NAND2_X1 U3301 ( .A1(wdata_a_i[17]), .A2(n7634), .ZN(n5250) );
  NAND2_X1 U3302 ( .A1(n8881), .A2(n4811), .ZN(n5251) );
  NAND2_X1 U3303 ( .A1(n5253), .A2(n5252), .ZN(n8556) );
  NAND2_X1 U3304 ( .A1(wdata_a_i[19]), .A2(n7658), .ZN(n5252) );
  NAND2_X1 U3305 ( .A1(n8877), .A2(n4809), .ZN(n5253) );
  NAND2_X1 U3306 ( .A1(n5255), .A2(n5254), .ZN(n8558) );
  NAND2_X1 U3307 ( .A1(wdata_a_i[17]), .A2(n7660), .ZN(n5254) );
  NAND2_X1 U3308 ( .A1(n8881), .A2(n4809), .ZN(n5255) );
  NAND2_X1 U3309 ( .A1(n5257), .A2(n5256), .ZN(n9121) );
  NAND2_X1 U3310 ( .A1(wdata_a_i[19]), .A2(n8011), .ZN(n5256) );
  NAND2_X1 U3311 ( .A1(n9164), .A2(n4818), .ZN(n5257) );
  NAND2_X1 U3312 ( .A1(n5259), .A2(n5258), .ZN(n8061) );
  NAND2_X1 U3313 ( .A1(wdata_a_i[23]), .A2(n7363), .ZN(n5258) );
  NAND2_X1 U3314 ( .A1(n4797), .A2(n4816), .ZN(n5259) );
  NAND2_X1 U3315 ( .A1(n5261), .A2(n5260), .ZN(n8064) );
  NAND2_X1 U3316 ( .A1(wdata_a_i[20]), .A2(n7364), .ZN(n5260) );
  NAND2_X1 U3317 ( .A1(n9162), .A2(n4816), .ZN(n5261) );
  NAND2_X1 U3318 ( .A1(n5263), .A2(n5262), .ZN(n8067) );
  NAND2_X1 U3319 ( .A1(wdata_a_i[17]), .A2(n7366), .ZN(n5262) );
  NAND2_X1 U3320 ( .A1(n4806), .A2(n4816), .ZN(n5263) );
  NAND2_X1 U3321 ( .A1(n5265), .A2(n5264), .ZN(n8096) );
  NAND2_X1 U3322 ( .A1(wdata_a_i[23]), .A2(n7392), .ZN(n5264) );
  NAND2_X1 U3323 ( .A1(n4775), .A2(n4822), .ZN(n5265) );
  NAND2_X1 U3324 ( .A1(n5267), .A2(n5266), .ZN(n8099) );
  NAND2_X1 U3325 ( .A1(wdata_a_i[20]), .A2(n7393), .ZN(n5266) );
  NAND2_X1 U3326 ( .A1(n9162), .A2(n4822), .ZN(n5267) );
  NAND2_X1 U3327 ( .A1(n5269), .A2(n5268), .ZN(n8100) );
  NAND2_X1 U3328 ( .A1(wdata_a_i[19]), .A2(n7394), .ZN(n5268) );
  NAND2_X1 U3329 ( .A1(n9164), .A2(n4822), .ZN(n5269) );
  NAND2_X1 U3330 ( .A1(n5271), .A2(n5270), .ZN(n8102) );
  NAND2_X1 U3331 ( .A1(wdata_a_i[17]), .A2(n7396), .ZN(n5270) );
  NAND2_X1 U3332 ( .A1(n9168), .A2(n4822), .ZN(n5271) );
  NAND2_X1 U3333 ( .A1(n5273), .A2(n5272), .ZN(n8131) );
  NAND2_X1 U3334 ( .A1(wdata_a_i[23]), .A2(n7406), .ZN(n5272) );
  NAND2_X1 U3335 ( .A1(n4776), .A2(n4815), .ZN(n5273) );
  NAND2_X1 U3336 ( .A1(n5275), .A2(n5274), .ZN(n8134) );
  NAND2_X1 U3337 ( .A1(wdata_a_i[20]), .A2(n7407), .ZN(n5274) );
  NAND2_X1 U3338 ( .A1(n9162), .A2(n4815), .ZN(n5275) );
  NAND2_X1 U3339 ( .A1(n5277), .A2(n5276), .ZN(n8137) );
  NAND2_X1 U3340 ( .A1(wdata_a_i[17]), .A2(n7409), .ZN(n5276) );
  NAND2_X1 U3341 ( .A1(n9078), .A2(n4815), .ZN(n5277) );
  NAND2_X1 U3342 ( .A1(n5279), .A2(n5278), .ZN(n8166) );
  NAND2_X1 U3343 ( .A1(wdata_a_i[23]), .A2(n7436), .ZN(n5278) );
  NAND2_X1 U3344 ( .A1(n4776), .A2(n4820), .ZN(n5279) );
  NAND2_X1 U3345 ( .A1(n5281), .A2(n5280), .ZN(n8169) );
  NAND2_X1 U3346 ( .A1(wdata_a_i[20]), .A2(n7437), .ZN(n5280) );
  NAND2_X1 U3347 ( .A1(n9162), .A2(n4820), .ZN(n5281) );
  NAND2_X1 U3348 ( .A1(n5283), .A2(n5282), .ZN(n8170) );
  NAND2_X1 U3349 ( .A1(wdata_a_i[19]), .A2(n7438), .ZN(n5282) );
  NAND2_X1 U3350 ( .A1(n9164), .A2(n4820), .ZN(n5283) );
  NAND2_X1 U3351 ( .A1(n5285), .A2(n5284), .ZN(n8172) );
  NAND2_X1 U3352 ( .A1(wdata_a_i[17]), .A2(n7440), .ZN(n5284) );
  NAND2_X1 U3353 ( .A1(n9168), .A2(n4820), .ZN(n5285) );
  NAND2_X1 U3354 ( .A1(n5287), .A2(n5286), .ZN(n8201) );
  NAND2_X1 U3355 ( .A1(wdata_a_i[23]), .A2(n7450), .ZN(n5286) );
  NAND2_X1 U3356 ( .A1(n4776), .A2(n4812), .ZN(n5287) );
  NAND2_X1 U3357 ( .A1(n5289), .A2(n5288), .ZN(n8204) );
  NAND2_X1 U3358 ( .A1(wdata_a_i[20]), .A2(n7451), .ZN(n5288) );
  NAND2_X1 U3359 ( .A1(n9162), .A2(n4812), .ZN(n5289) );
  NAND2_X1 U3360 ( .A1(n5291), .A2(n5290), .ZN(n8207) );
  NAND2_X1 U3361 ( .A1(wdata_a_i[17]), .A2(n7453), .ZN(n5290) );
  NAND2_X1 U3362 ( .A1(n9078), .A2(n4812), .ZN(n5291) );
  NAND2_X1 U3363 ( .A1(n5293), .A2(n5292), .ZN(n8271) );
  NAND2_X1 U3364 ( .A1(wdata_a_i[23]), .A2(n7473), .ZN(n5292) );
  NAND2_X1 U3365 ( .A1(n4775), .A2(n4819), .ZN(n5293) );
  NAND2_X1 U3366 ( .A1(n5295), .A2(n5294), .ZN(n8274) );
  NAND2_X1 U3367 ( .A1(wdata_a_i[20]), .A2(n7474), .ZN(n5294) );
  NAND2_X1 U3368 ( .A1(n9162), .A2(n4819), .ZN(n5295) );
  NAND2_X1 U3369 ( .A1(n5297), .A2(n5296), .ZN(n8277) );
  NAND2_X1 U3370 ( .A1(wdata_a_i[17]), .A2(n7476), .ZN(n5296) );
  NAND2_X1 U3371 ( .A1(n4805), .A2(n4819), .ZN(n5297) );
  NAND2_X1 U3372 ( .A1(n5299), .A2(n5298), .ZN(n8306) );
  NAND2_X1 U3373 ( .A1(wdata_a_i[23]), .A2(n7495), .ZN(n5298) );
  NAND2_X1 U3374 ( .A1(n9157), .A2(n4746), .ZN(n5299) );
  NAND2_X1 U3375 ( .A1(n5301), .A2(n5300), .ZN(n8309) );
  NAND2_X1 U3376 ( .A1(wdata_a_i[20]), .A2(n7496), .ZN(n5300) );
  NAND2_X1 U3377 ( .A1(n9162), .A2(n4746), .ZN(n5301) );
  NAND2_X1 U3378 ( .A1(n5303), .A2(n5302), .ZN(n8312) );
  NAND2_X1 U3379 ( .A1(wdata_a_i[17]), .A2(n7497), .ZN(n5302) );
  NAND2_X1 U3380 ( .A1(n9168), .A2(n4746), .ZN(n5303) );
  NAND2_X1 U3381 ( .A1(n5305), .A2(n5304), .ZN(n8341) );
  NAND2_X1 U3382 ( .A1(wdata_a_i[23]), .A2(n7518), .ZN(n5304) );
  NAND2_X1 U3383 ( .A1(n4797), .A2(n4817), .ZN(n5305) );
  NAND2_X1 U3384 ( .A1(n5307), .A2(n5306), .ZN(n8344) );
  NAND2_X1 U3385 ( .A1(wdata_a_i[20]), .A2(n7519), .ZN(n5306) );
  NAND2_X1 U3386 ( .A1(n9162), .A2(n4817), .ZN(n5307) );
  NAND2_X1 U3387 ( .A1(n5309), .A2(n5308), .ZN(n8345) );
  NAND2_X1 U3388 ( .A1(wdata_a_i[19]), .A2(n7520), .ZN(n5308) );
  NAND2_X1 U3389 ( .A1(n9164), .A2(n4817), .ZN(n5309) );
  NAND2_X1 U3390 ( .A1(n5311), .A2(n5310), .ZN(n8347) );
  NAND2_X1 U3391 ( .A1(wdata_a_i[17]), .A2(n7521), .ZN(n5310) );
  NAND2_X1 U3392 ( .A1(n4806), .A2(n4817), .ZN(n5311) );
  NAND2_X1 U3393 ( .A1(n5313), .A2(n5312), .ZN(n8377) );
  NAND2_X1 U3394 ( .A1(wdata_a_i[23]), .A2(n7540), .ZN(n5312) );
  NAND2_X1 U3395 ( .A1(n4775), .A2(n4807), .ZN(n5313) );
  NAND2_X1 U3396 ( .A1(n5315), .A2(n5314), .ZN(n8380) );
  NAND2_X1 U3397 ( .A1(wdata_a_i[20]), .A2(n7541), .ZN(n5314) );
  NAND2_X1 U3398 ( .A1(n9162), .A2(n4807), .ZN(n5315) );
  NAND2_X1 U3399 ( .A1(n5317), .A2(n5316), .ZN(n8381) );
  NAND2_X1 U3400 ( .A1(wdata_a_i[19]), .A2(n7541), .ZN(n5316) );
  NAND2_X1 U3401 ( .A1(n9164), .A2(n4807), .ZN(n5317) );
  NAND2_X1 U3402 ( .A1(n5319), .A2(n5318), .ZN(n8383) );
  NAND2_X1 U3403 ( .A1(wdata_a_i[17]), .A2(n7542), .ZN(n5318) );
  NAND2_X1 U3404 ( .A1(n4805), .A2(n4807), .ZN(n5319) );
  NAND2_X1 U3405 ( .A1(n5321), .A2(n5320), .ZN(n9117) );
  NAND2_X1 U3406 ( .A1(wdata_a_i[23]), .A2(n8009), .ZN(n5320) );
  NAND2_X1 U3407 ( .A1(n4776), .A2(n4818), .ZN(n5321) );
  NAND2_X1 U3408 ( .A1(n5323), .A2(n5322), .ZN(n9120) );
  NAND2_X1 U3409 ( .A1(wdata_a_i[20]), .A2(n8010), .ZN(n5322) );
  NAND2_X1 U3410 ( .A1(n9162), .A2(n4818), .ZN(n5323) );
  NAND2_X1 U3411 ( .A1(n5325), .A2(n5324), .ZN(n9123) );
  NAND2_X1 U3412 ( .A1(wdata_a_i[17]), .A2(n8012), .ZN(n5324) );
  NAND2_X1 U3413 ( .A1(n4805), .A2(n4818), .ZN(n5325) );
  NAND2_X1 U3414 ( .A1(n5327), .A2(n5326), .ZN(n8066) );
  NAND2_X1 U3416 ( .A1(wdata_a_i[18]), .A2(n7365), .ZN(n5326) );
  NAND2_X1 U3418 ( .A1(n9166), .A2(n4816), .ZN(n5327) );
  NAND2_X1 U3419 ( .A1(n5329), .A2(n5328), .ZN(n8101) );
  NAND2_X1 U3420 ( .A1(wdata_a_i[18]), .A2(n7394), .ZN(n5328) );
  NAND2_X1 U3421 ( .A1(n9166), .A2(n4822), .ZN(n5329) );
  NAND2_X1 U3422 ( .A1(n5331), .A2(n5330), .ZN(n8136) );
  NAND2_X1 U3423 ( .A1(wdata_a_i[18]), .A2(n7408), .ZN(n5330) );
  NAND2_X1 U3424 ( .A1(n9166), .A2(n4815), .ZN(n5331) );
  NAND2_X1 U3425 ( .A1(n5333), .A2(n5332), .ZN(n8171) );
  NAND2_X1 U3426 ( .A1(wdata_a_i[18]), .A2(n7438), .ZN(n5332) );
  NAND2_X1 U3427 ( .A1(n9166), .A2(n4820), .ZN(n5333) );
  NAND2_X1 U3428 ( .A1(n5335), .A2(n5334), .ZN(n8206) );
  NAND2_X1 U3429 ( .A1(wdata_a_i[18]), .A2(n7452), .ZN(n5334) );
  NAND2_X1 U3430 ( .A1(n9166), .A2(n4812), .ZN(n5335) );
  NAND2_X1 U3431 ( .A1(n5337), .A2(n5336), .ZN(n8276) );
  NAND2_X1 U3432 ( .A1(wdata_a_i[18]), .A2(n7475), .ZN(n5336) );
  NAND2_X1 U3433 ( .A1(n9166), .A2(n4819), .ZN(n5337) );
  NAND2_X1 U3434 ( .A1(n5339), .A2(n5338), .ZN(n8311) );
  NAND2_X1 U3435 ( .A1(wdata_a_i[18]), .A2(n7497), .ZN(n5338) );
  NAND2_X1 U3436 ( .A1(n9166), .A2(n4746), .ZN(n5339) );
  NAND2_X1 U3437 ( .A1(n5341), .A2(n5340), .ZN(n8346) );
  NAND2_X1 U3438 ( .A1(wdata_a_i[18]), .A2(n7520), .ZN(n5340) );
  NAND2_X1 U3439 ( .A1(n9166), .A2(n4817), .ZN(n5341) );
  NAND2_X1 U3440 ( .A1(n5343), .A2(n5342), .ZN(n8382) );
  NAND2_X1 U3441 ( .A1(wdata_a_i[18]), .A2(n7542), .ZN(n5342) );
  NAND2_X1 U3442 ( .A1(n4793), .A2(n4807), .ZN(n5343) );
  NAND2_X1 U3443 ( .A1(n5345), .A2(n5344), .ZN(n8447) );
  NAND2_X1 U3444 ( .A1(wdata_a_i[23]), .A2(n7585), .ZN(n5344) );
  NAND2_X1 U3445 ( .A1(n4776), .A2(n4810), .ZN(n5345) );
  NAND2_X1 U3446 ( .A1(n5347), .A2(n5346), .ZN(n8450) );
  NAND2_X1 U3447 ( .A1(wdata_a_i[20]), .A2(n7586), .ZN(n5346) );
  NAND2_X1 U3448 ( .A1(n8875), .A2(n4810), .ZN(n5347) );
  NAND2_X1 U3449 ( .A1(n5349), .A2(n5348), .ZN(n8482) );
  NAND2_X1 U3450 ( .A1(wdata_a_i[23]), .A2(n7609), .ZN(n5348) );
  NAND2_X1 U3451 ( .A1(n4775), .A2(n4808), .ZN(n5349) );
  NAND2_X1 U3452 ( .A1(n5351), .A2(n5350), .ZN(n8485) );
  NAND2_X1 U3453 ( .A1(wdata_a_i[20]), .A2(n7610), .ZN(n5350) );
  NAND2_X1 U3454 ( .A1(n8875), .A2(n4808), .ZN(n5351) );
  NAND2_X1 U3455 ( .A1(n5353), .A2(n5352), .ZN(n8517) );
  NAND2_X1 U3456 ( .A1(wdata_a_i[23]), .A2(n7632), .ZN(n5352) );
  NAND2_X1 U3457 ( .A1(n4776), .A2(n4811), .ZN(n5353) );
  NAND2_X1 U3458 ( .A1(n5355), .A2(n5354), .ZN(n8520) );
  NAND2_X1 U3459 ( .A1(wdata_a_i[20]), .A2(n7633), .ZN(n5354) );
  NAND2_X1 U3460 ( .A1(n8875), .A2(n4811), .ZN(n5355) );
  NAND2_X1 U3461 ( .A1(n5357), .A2(n5356), .ZN(n8552) );
  NAND2_X1 U3462 ( .A1(wdata_a_i[23]), .A2(n7656), .ZN(n5356) );
  NAND2_X1 U3463 ( .A1(n4797), .A2(n4809), .ZN(n5357) );
  NAND2_X1 U3464 ( .A1(n5359), .A2(n5358), .ZN(n8555) );
  NAND2_X1 U3465 ( .A1(wdata_a_i[20]), .A2(n7657), .ZN(n5358) );
  NAND2_X1 U3466 ( .A1(n8875), .A2(n4809), .ZN(n5359) );
  NAND2_X1 U3467 ( .A1(n5361), .A2(n5360), .ZN(n9122) );
  NAND2_X1 U3468 ( .A1(wdata_a_i[18]), .A2(n8011), .ZN(n5360) );
  NAND2_X1 U3469 ( .A1(n9166), .A2(n4818), .ZN(n5361) );
  NAND2_X1 U3470 ( .A1(n5363), .A2(n5362), .ZN(n8452) );
  NAND2_X1 U3471 ( .A1(wdata_a_i[18]), .A2(n7587), .ZN(n5362) );
  NAND2_X1 U3472 ( .A1(n4793), .A2(n4810), .ZN(n5363) );
  NAND2_X1 U3473 ( .A1(n5365), .A2(n5364), .ZN(n8487) );
  NAND2_X1 U3474 ( .A1(wdata_a_i[18]), .A2(n7611), .ZN(n5364) );
  NAND2_X1 U3475 ( .A1(n5367), .A2(n5366), .ZN(n8522) );
  NAND2_X1 U3476 ( .A1(wdata_a_i[18]), .A2(n7634), .ZN(n5366) );
  NAND2_X1 U3477 ( .A1(n4792), .A2(n4811), .ZN(n5367) );
  NAND2_X1 U3478 ( .A1(n5369), .A2(n5368), .ZN(n8557) );
  NAND2_X1 U3479 ( .A1(wdata_a_i[18]), .A2(n7658), .ZN(n5368) );
  NAND2_X1 U3480 ( .A1(n8879), .A2(n4809), .ZN(n5369) );
  NAND2_X1 U3481 ( .A1(n5371), .A2(n5370), .ZN(n8440) );
  NAND2_X1 U3482 ( .A1(n4623), .A2(n7584), .ZN(n5370) );
  NAND2_X1 U3483 ( .A1(n8861), .A2(n4810), .ZN(n5371) );
  NAND2_X1 U3484 ( .A1(n5373), .A2(n5372), .ZN(n8475) );
  NAND2_X1 U3485 ( .A1(n4623), .A2(n7608), .ZN(n5372) );
  NAND2_X1 U3486 ( .A1(n8861), .A2(n4808), .ZN(n5373) );
  NAND2_X1 U3487 ( .A1(n5375), .A2(n5374), .ZN(n8510) );
  NAND2_X1 U3488 ( .A1(n4623), .A2(n7631), .ZN(n5374) );
  NAND2_X1 U3489 ( .A1(n8861), .A2(n4811), .ZN(n5375) );
  NAND2_X1 U3490 ( .A1(n5377), .A2(n5376), .ZN(n8545) );
  NAND2_X1 U3491 ( .A1(n4623), .A2(n7655), .ZN(n5376) );
  NAND2_X1 U3492 ( .A1(n8861), .A2(n4809), .ZN(n5377) );
  INV_X1 U3493 ( .A(wdata_b_i[31]), .ZN(n4474) );
  INV_X2 U3494 ( .A(n4047), .ZN(n9155) );
  INV_X1 U3495 ( .A(wdata_b_i[9]), .ZN(n4426) );
  NOR2_X1 U5481 ( .A1(n1546), .A2(n4816), .ZN(n7362) );
  MUX2_X1 U5482 ( .A(n4468), .B(n4803), .S(n4816), .Z(n8055) );
  MUX2_X1 U5483 ( .A(n4618), .B(wdata_b_i[28]), .S(n4816), .Z(n8056) );
  MUX2_X1 U5484 ( .A(n4394), .B(n4732), .S(n4816), .Z(n8057) );
  MUX2_X1 U5485 ( .A(n4459), .B(n8867), .S(n4816), .Z(n8058) );
  MUX2_X1 U5486 ( .A(n4614), .B(wdata_b_i[25]), .S(n4816), .Z(n8059) );
  MUX2_X1 U5487 ( .A(n4386), .B(n9155), .S(n4816), .Z(n8060) );
  NOR2_X1 U5488 ( .A1(n1546), .A2(n4816), .ZN(n7363) );
  NOR2_X1 U5489 ( .A1(n1546), .A2(n4816), .ZN(n7364) );
  NOR2_X1 U5490 ( .A1(n1546), .A2(n4816), .ZN(n7365) );
  MUX2_X1 U5491 ( .A(wdata_a_i[16]), .B(n8349), .S(n4816), .Z(n8068) );
  NOR2_X1 U5492 ( .A1(n1546), .A2(n4816), .ZN(n7366) );
  MUX2_X1 U5493 ( .A(wdata_a_i[14]), .B(n9172), .S(n4816), .Z(n8070) );
  MUX2_X1 U5494 ( .A(wdata_a_i[13]), .B(n9174), .S(n4816), .Z(n8071) );
  MUX2_X1 U5495 ( .A(wdata_a_i[12]), .B(n9085), .S(n4816), .Z(n8072) );
  INV_X1 U5496 ( .A(n7367), .ZN(n8073) );
  AOI22_X1 U5497 ( .A1(wdata_a_i[11]), .A2(n7368), .B1(n4816), .B2(n8892), 
        .ZN(n7367) );
  NOR2_X1 U5498 ( .A1(n1546), .A2(n4816), .ZN(n7368) );
  INV_X1 U5499 ( .A(n7369), .ZN(n8075) );
  AOI22_X1 U5500 ( .A1(wdata_a_i[9]), .A2(n7371), .B1(n4816), .B2(n9091), .ZN(
        n7369) );
  INV_X1 U5501 ( .A(n7370), .ZN(n8076) );
  AOI22_X1 U5502 ( .A1(wdata_a_i[8]), .A2(n7371), .B1(n4816), .B2(n4774), .ZN(
        n7370) );
  NOR2_X1 U5503 ( .A1(n1546), .A2(n4816), .ZN(n7371) );
  INV_X1 U5504 ( .A(n7372), .ZN(n8077) );
  AOI22_X1 U5505 ( .A1(n4486), .A2(n7374), .B1(n4816), .B2(n4780), .ZN(n7372)
         );
  INV_X1 U5506 ( .A(n7373), .ZN(n8078) );
  AOI22_X1 U5507 ( .A1(wdata_a_i[6]), .A2(n7374), .B1(n4816), .B2(n9184), .ZN(
        n7373) );
  NOR2_X1 U5508 ( .A1(n1546), .A2(n4816), .ZN(n7374) );
  INV_X1 U5509 ( .A(n7375), .ZN(n8079) );
  AOI22_X1 U5510 ( .A1(wdata_a_i[5]), .A2(n7377), .B1(n4816), .B2(n9186), .ZN(
        n7375) );
  INV_X1 U5511 ( .A(n7376), .ZN(n8080) );
  AOI22_X1 U5512 ( .A1(wdata_a_i[4]), .A2(n7377), .B1(n4816), .B2(n4787), .ZN(
        n7376) );
  NOR2_X1 U5513 ( .A1(n1546), .A2(n4816), .ZN(n7377) );
  INV_X1 U5514 ( .A(n7378), .ZN(n8081) );
  AOI22_X1 U5515 ( .A1(wdata_a_i[3]), .A2(n7380), .B1(n4816), .B2(n9189), .ZN(
        n7378) );
  INV_X1 U5516 ( .A(n7379), .ZN(n8082) );
  AOI22_X1 U5517 ( .A1(wdata_a_i[2]), .A2(n7380), .B1(n4816), .B2(n9191), .ZN(
        n7379) );
  NOR2_X1 U5518 ( .A1(n1546), .A2(n4816), .ZN(n7380) );
  INV_X1 U5519 ( .A(n7381), .ZN(n8083) );
  AOI22_X1 U5520 ( .A1(wdata_a_i[1]), .A2(n7383), .B1(n4816), .B2(n9193), .ZN(
        n7381) );
  INV_X1 U5521 ( .A(n7382), .ZN(n8084) );
  AOI22_X1 U5522 ( .A1(wdata_a_i[0]), .A2(n7383), .B1(n4816), .B2(n4790), .ZN(
        n7382) );
  NOR2_X1 U5523 ( .A1(n1546), .A2(n4816), .ZN(n7383) );
  OR2_X1 U5524 ( .A1(n1548), .A2(n4816), .ZN(n8087) );
  NOR2_X1 U5525 ( .A1(n1587), .A2(n4822), .ZN(n7384) );
  INV_X1 U5526 ( .A(n7385), .ZN(n8091) );
  AOI22_X1 U5527 ( .A1(n4618), .A2(n7386), .B1(n4822), .B2(wdata_b_i[28]), 
        .ZN(n7385) );
  NOR2_X1 U5528 ( .A1(n1587), .A2(n4822), .ZN(n7386) );
  INV_X1 U5529 ( .A(n7387), .ZN(n8092) );
  AOI22_X1 U5530 ( .A1(n4394), .A2(n7388), .B1(n4822), .B2(n9150), .ZN(n7387)
         );
  NOR2_X1 U5531 ( .A1(n1587), .A2(n4822), .ZN(n7388) );
  INV_X1 U5532 ( .A(n7389), .ZN(n8094) );
  AOI22_X1 U5533 ( .A1(n4614), .A2(n7391), .B1(n4822), .B2(wdata_b_i[25]), 
        .ZN(n7389) );
  INV_X1 U5534 ( .A(n7390), .ZN(n8095) );
  AOI22_X1 U5535 ( .A1(n4386), .A2(n7391), .B1(n4822), .B2(n9155), .ZN(n7390)
         );
  NOR2_X1 U5536 ( .A1(n1587), .A2(n4822), .ZN(n7391) );
  NOR2_X1 U5537 ( .A1(n1587), .A2(n4822), .ZN(n7392) );
  NOR2_X1 U5538 ( .A1(n1587), .A2(n4822), .ZN(n7393) );
  NOR2_X1 U5539 ( .A1(n1587), .A2(n4822), .ZN(n7394) );
  INV_X1 U5540 ( .A(n7395), .ZN(n8103) );
  AOI22_X1 U5541 ( .A1(wdata_a_i[16]), .A2(n7396), .B1(n4822), .B2(n8349), 
        .ZN(n7395) );
  NOR2_X1 U5542 ( .A1(n1587), .A2(n4822), .ZN(n7396) );
  MUX2_X1 U5543 ( .A(wdata_a_i[14]), .B(n9172), .S(n4822), .Z(n8105) );
  MUX2_X1 U5544 ( .A(wdata_a_i[13]), .B(n9174), .S(n4822), .Z(n8106) );
  MUX2_X1 U5545 ( .A(wdata_a_i[12]), .B(n9085), .S(n4822), .Z(n8107) );
  MUX2_X1 U5546 ( .A(wdata_a_i[11]), .B(n4782), .S(n4822), .Z(n8108) );
  MUX2_X1 U5547 ( .A(wdata_a_i[10]), .B(n9178), .S(n4822), .Z(n8109) );
  MUX2_X1 U5548 ( .A(wdata_a_i[9]), .B(n4783), .S(n4822), .Z(n8110) );
  MUX2_X1 U5549 ( .A(wdata_a_i[8]), .B(n8898), .S(n4822), .Z(n8111) );
  MUX2_X1 U5550 ( .A(n4486), .B(n4779), .S(n4822), .Z(n8112) );
  MUX2_X1 U5551 ( .A(wdata_a_i[6]), .B(n9184), .S(n4822), .Z(n8113) );
  INV_X1 U5552 ( .A(n7397), .ZN(n8114) );
  AOI22_X1 U5553 ( .A1(wdata_a_i[5]), .A2(n7398), .B1(n4822), .B2(n9096), .ZN(
        n7397) );
  NOR2_X1 U5554 ( .A1(n1587), .A2(n4822), .ZN(n7398) );
  INV_X1 U5555 ( .A(n7399), .ZN(n8115) );
  AOI22_X1 U5556 ( .A1(wdata_a_i[4]), .A2(n7401), .B1(n4822), .B2(n9098), .ZN(
        n7399) );
  MUX2_X1 U5557 ( .A(wdata_a_i[3]), .B(n9100), .S(n4822), .Z(n8116) );
  INV_X1 U5558 ( .A(n7400), .ZN(n8117) );
  AOI22_X1 U5559 ( .A1(wdata_a_i[2]), .A2(n7401), .B1(n4822), .B2(n9191), .ZN(
        n7400) );
  NOR2_X1 U5560 ( .A1(n1587), .A2(n4822), .ZN(n7401) );
  INV_X1 U5561 ( .A(n7402), .ZN(n8118) );
  AOI22_X1 U5562 ( .A1(wdata_a_i[1]), .A2(n7404), .B1(n4822), .B2(n9193), .ZN(
        n7402) );
  INV_X1 U5563 ( .A(n7403), .ZN(n8119) );
  AOI22_X1 U5564 ( .A1(wdata_a_i[0]), .A2(n7404), .B1(n4822), .B2(n4791), .ZN(
        n7403) );
  NOR2_X1 U5565 ( .A1(n1587), .A2(n4822), .ZN(n7404) );
  NAND2_X1 U5566 ( .A1(n1587), .A2(n4751), .ZN(n8122) );
  NOR2_X1 U5567 ( .A1(n1577), .A2(n4815), .ZN(n7405) );
  MUX2_X1 U5568 ( .A(n4468), .B(n4803), .S(n4815), .Z(n8125) );
  MUX2_X1 U5569 ( .A(n4618), .B(wdata_b_i[28]), .S(n4815), .Z(n8126) );
  MUX2_X1 U5570 ( .A(n4394), .B(n8865), .S(n4815), .Z(n8127) );
  MUX2_X1 U5571 ( .A(n4459), .B(n9152), .S(n4815), .Z(n8128) );
  MUX2_X1 U5572 ( .A(n4614), .B(wdata_b_i[25]), .S(n4815), .Z(n8129) );
  MUX2_X1 U5573 ( .A(n4386), .B(n9155), .S(n4815), .Z(n8130) );
  NOR2_X1 U5574 ( .A1(n1577), .A2(n4815), .ZN(n7406) );
  NOR2_X1 U5575 ( .A1(n1577), .A2(n4815), .ZN(n7407) );
  NOR2_X1 U5576 ( .A1(n1577), .A2(n4815), .ZN(n7408) );
  MUX2_X1 U5577 ( .A(wdata_a_i[16]), .B(n4734), .S(n4815), .Z(n8138) );
  NOR2_X1 U5578 ( .A1(n1577), .A2(n4815), .ZN(n7409) );
  MUX2_X1 U5579 ( .A(wdata_a_i[14]), .B(n9172), .S(n4815), .Z(n8140) );
  MUX2_X1 U5580 ( .A(wdata_a_i[13]), .B(n9174), .S(n4815), .Z(n8141) );
  MUX2_X1 U5581 ( .A(wdata_a_i[12]), .B(n9085), .S(n4815), .Z(n8142) );
  INV_X1 U5582 ( .A(n7410), .ZN(n8143) );
  AOI22_X1 U5583 ( .A1(wdata_a_i[11]), .A2(n7411), .B1(n4815), .B2(n9087), 
        .ZN(n7410) );
  NOR2_X1 U5584 ( .A1(n1577), .A2(n4815), .ZN(n7411) );
  INV_X1 U5585 ( .A(n7412), .ZN(n8145) );
  AOI22_X1 U5586 ( .A1(wdata_a_i[9]), .A2(n7414), .B1(n4815), .B2(n9091), .ZN(
        n7412) );
  INV_X1 U5587 ( .A(n7413), .ZN(n8146) );
  AOI22_X1 U5588 ( .A1(wdata_a_i[8]), .A2(n7414), .B1(n4815), .B2(n4774), .ZN(
        n7413) );
  NOR2_X1 U5589 ( .A1(n1577), .A2(n4815), .ZN(n7414) );
  INV_X1 U5590 ( .A(n7415), .ZN(n8147) );
  AOI22_X1 U5591 ( .A1(wdata_a_i[7]), .A2(n7417), .B1(n4815), .B2(n4779), .ZN(
        n7415) );
  INV_X1 U5592 ( .A(n7416), .ZN(n8148) );
  AOI22_X1 U5593 ( .A1(wdata_a_i[6]), .A2(n7417), .B1(n4815), .B2(n9184), .ZN(
        n7416) );
  NOR2_X1 U5594 ( .A1(n1577), .A2(n4815), .ZN(n7417) );
  INV_X1 U5595 ( .A(n7418), .ZN(n8149) );
  AOI22_X1 U5596 ( .A1(wdata_a_i[5]), .A2(n7420), .B1(n4815), .B2(n8902), .ZN(
        n7418) );
  INV_X1 U5597 ( .A(n7419), .ZN(n8150) );
  AOI22_X1 U5598 ( .A1(wdata_a_i[4]), .A2(n7420), .B1(n4815), .B2(n4787), .ZN(
        n7419) );
  NOR2_X1 U5599 ( .A1(n1577), .A2(n4815), .ZN(n7420) );
  INV_X1 U5600 ( .A(n7421), .ZN(n8151) );
  AOI22_X1 U5601 ( .A1(wdata_a_i[3]), .A2(n7423), .B1(n4815), .B2(n9189), .ZN(
        n7421) );
  INV_X1 U5602 ( .A(n7422), .ZN(n8152) );
  AOI22_X1 U5603 ( .A1(wdata_a_i[2]), .A2(n7423), .B1(n4815), .B2(n9191), .ZN(
        n7422) );
  NOR2_X1 U5604 ( .A1(n1577), .A2(n4815), .ZN(n7423) );
  INV_X1 U5605 ( .A(n7424), .ZN(n8153) );
  AOI22_X1 U5606 ( .A1(wdata_a_i[1]), .A2(n7426), .B1(n4815), .B2(n9193), .ZN(
        n7424) );
  INV_X1 U5607 ( .A(n7425), .ZN(n8154) );
  AOI22_X1 U5608 ( .A1(wdata_a_i[0]), .A2(n7426), .B1(n4815), .B2(n9195), .ZN(
        n7425) );
  NOR2_X1 U5609 ( .A1(n1577), .A2(n4815), .ZN(n7426) );
  OR2_X1 U5610 ( .A1(n1579), .A2(n4815), .ZN(n8157) );
  NOR2_X1 U5611 ( .A1(n1571), .A2(n4820), .ZN(n7427) );
  INV_X1 U5612 ( .A(n7428), .ZN(n8160) );
  AOI22_X1 U5613 ( .A1(n4468), .A2(n7430), .B1(n4820), .B2(n4796), .ZN(n7428)
         );
  INV_X1 U5614 ( .A(n7429), .ZN(n8161) );
  AOI22_X1 U5615 ( .A1(n4618), .A2(n7430), .B1(n4820), .B2(wdata_b_i[28]), 
        .ZN(n7429) );
  NOR2_X1 U5616 ( .A1(n1571), .A2(n4820), .ZN(n7430) );
  INV_X1 U5617 ( .A(n7431), .ZN(n8162) );
  AOI22_X1 U5618 ( .A1(n4394), .A2(n7432), .B1(n4820), .B2(n9150), .ZN(n7431)
         );
  NOR2_X1 U5619 ( .A1(n1571), .A2(n4820), .ZN(n7432) );
  INV_X1 U5620 ( .A(n7433), .ZN(n8164) );
  AOI22_X1 U5621 ( .A1(n4614), .A2(n7435), .B1(n4820), .B2(wdata_b_i[25]), 
        .ZN(n7433) );
  INV_X1 U5622 ( .A(n7434), .ZN(n8165) );
  AOI22_X1 U5623 ( .A1(n4386), .A2(n7435), .B1(n4820), .B2(n9155), .ZN(n7434)
         );
  NOR2_X1 U5624 ( .A1(n1571), .A2(n4820), .ZN(n7435) );
  NOR2_X1 U5625 ( .A1(n1571), .A2(n4820), .ZN(n7436) );
  NOR2_X1 U5626 ( .A1(n1571), .A2(n4820), .ZN(n7437) );
  NOR2_X1 U5627 ( .A1(n1571), .A2(n4820), .ZN(n7438) );
  INV_X1 U5628 ( .A(n7439), .ZN(n8173) );
  AOI22_X1 U5629 ( .A1(wdata_a_i[16]), .A2(n7440), .B1(n4820), .B2(n8349), 
        .ZN(n7439) );
  NOR2_X1 U5630 ( .A1(n1571), .A2(n4820), .ZN(n7440) );
  MUX2_X1 U5631 ( .A(wdata_a_i[14]), .B(n9172), .S(n4820), .Z(n8175) );
  MUX2_X1 U5632 ( .A(wdata_a_i[13]), .B(n9174), .S(n4820), .Z(n8176) );
  MUX2_X1 U5633 ( .A(wdata_a_i[12]), .B(n9085), .S(n4820), .Z(n8177) );
  MUX2_X1 U5634 ( .A(wdata_a_i[11]), .B(n4782), .S(n4820), .Z(n8178) );
  MUX2_X1 U5635 ( .A(wdata_a_i[10]), .B(n9178), .S(n4820), .Z(n8179) );
  MUX2_X1 U5636 ( .A(wdata_a_i[9]), .B(n4783), .S(n4820), .Z(n8180) );
  MUX2_X1 U5637 ( .A(wdata_a_i[8]), .B(n8898), .S(n4820), .Z(n8181) );
  MUX2_X1 U5638 ( .A(n4486), .B(n8848), .S(n4820), .Z(n8182) );
  INV_X1 U5639 ( .A(n7441), .ZN(n8183) );
  AOI22_X1 U5640 ( .A1(wdata_a_i[6]), .A2(n7442), .B1(n4820), .B2(n9184), .ZN(
        n7441) );
  NOR2_X1 U5641 ( .A1(n1571), .A2(n4820), .ZN(n7442) );
  MUX2_X1 U5642 ( .A(wdata_a_i[5]), .B(n9096), .S(n4820), .Z(n8184) );
  INV_X1 U5643 ( .A(n7443), .ZN(n8185) );
  AOI22_X1 U5644 ( .A1(wdata_a_i[4]), .A2(n7445), .B1(n4820), .B2(n9098), .ZN(
        n7443) );
  MUX2_X1 U5645 ( .A(wdata_a_i[3]), .B(n8906), .S(n4820), .Z(n8186) );
  INV_X1 U5646 ( .A(n7444), .ZN(n8187) );
  AOI22_X1 U5647 ( .A1(wdata_a_i[2]), .A2(n7445), .B1(n4820), .B2(n9191), .ZN(
        n7444) );
  NOR2_X1 U5648 ( .A1(n1571), .A2(n4820), .ZN(n7445) );
  INV_X1 U5649 ( .A(n7446), .ZN(n8188) );
  AOI22_X1 U5650 ( .A1(wdata_a_i[1]), .A2(n7448), .B1(n4820), .B2(n4786), .ZN(
        n7446) );
  INV_X1 U5651 ( .A(n7447), .ZN(n8189) );
  AOI22_X1 U5652 ( .A1(wdata_a_i[0]), .A2(n7448), .B1(n4820), .B2(n9195), .ZN(
        n7447) );
  NOR2_X1 U5653 ( .A1(n1571), .A2(n4820), .ZN(n7448) );
  NAND2_X1 U5654 ( .A1(n1571), .A2(n4755), .ZN(n8192) );
  NOR2_X1 U5655 ( .A1(n1581), .A2(n4812), .ZN(n7449) );
  MUX2_X1 U5656 ( .A(n4468), .B(n4803), .S(n4812), .Z(n8195) );
  MUX2_X1 U5657 ( .A(n4618), .B(wdata_b_i[28]), .S(n4812), .Z(n8196) );
  MUX2_X1 U5658 ( .A(n4394), .B(n4732), .S(n4812), .Z(n8197) );
  MUX2_X1 U5659 ( .A(n4459), .B(n8867), .S(n4812), .Z(n8198) );
  MUX2_X1 U5660 ( .A(n4614), .B(wdata_b_i[25]), .S(n4812), .Z(n8199) );
  MUX2_X1 U5661 ( .A(n4386), .B(n9155), .S(n4812), .Z(n8200) );
  NOR2_X1 U5662 ( .A1(n1581), .A2(n4812), .ZN(n7450) );
  NOR2_X1 U5663 ( .A1(n1581), .A2(n4812), .ZN(n7451) );
  NOR2_X1 U5664 ( .A1(n1581), .A2(n4812), .ZN(n7452) );
  MUX2_X1 U5665 ( .A(wdata_a_i[16]), .B(n8349), .S(n4812), .Z(n8208) );
  NOR2_X1 U5666 ( .A1(n1581), .A2(n4812), .ZN(n7453) );
  MUX2_X1 U5667 ( .A(wdata_a_i[14]), .B(n9172), .S(n4812), .Z(n8210) );
  MUX2_X1 U5668 ( .A(wdata_a_i[13]), .B(n9174), .S(n4812), .Z(n8211) );
  MUX2_X1 U5669 ( .A(wdata_a_i[12]), .B(n9085), .S(n4812), .Z(n8212) );
  INV_X1 U5670 ( .A(n7454), .ZN(n8213) );
  AOI22_X1 U5671 ( .A1(wdata_a_i[11]), .A2(n7455), .B1(n4812), .B2(n8892), 
        .ZN(n7454) );
  NOR2_X1 U5672 ( .A1(n1581), .A2(n4812), .ZN(n7455) );
  INV_X1 U5673 ( .A(n7456), .ZN(n8215) );
  AOI22_X1 U5674 ( .A1(wdata_a_i[9]), .A2(n7458), .B1(n4812), .B2(n9091), .ZN(
        n7456) );
  INV_X1 U5675 ( .A(n7457), .ZN(n8216) );
  AOI22_X1 U5676 ( .A1(wdata_a_i[8]), .A2(n7458), .B1(n4812), .B2(n4774), .ZN(
        n7457) );
  NOR2_X1 U5677 ( .A1(n1581), .A2(n4812), .ZN(n7458) );
  INV_X1 U5678 ( .A(n7459), .ZN(n8217) );
  AOI22_X1 U5679 ( .A1(n4486), .A2(n7461), .B1(n4812), .B2(n4779), .ZN(n7459)
         );
  INV_X1 U5680 ( .A(n7460), .ZN(n8218) );
  AOI22_X1 U5681 ( .A1(wdata_a_i[6]), .A2(n7461), .B1(n4812), .B2(n9184), .ZN(
        n7460) );
  NOR2_X1 U5682 ( .A1(n1581), .A2(n4812), .ZN(n7461) );
  INV_X1 U5683 ( .A(n7462), .ZN(n8219) );
  AOI22_X1 U5684 ( .A1(wdata_a_i[5]), .A2(n7464), .B1(n4812), .B2(n9096), .ZN(
        n7462) );
  INV_X1 U5685 ( .A(n7463), .ZN(n8220) );
  AOI22_X1 U5686 ( .A1(wdata_a_i[4]), .A2(n7464), .B1(n4812), .B2(n4787), .ZN(
        n7463) );
  NOR2_X1 U5687 ( .A1(n1581), .A2(n4812), .ZN(n7464) );
  INV_X1 U5688 ( .A(n7465), .ZN(n8221) );
  AOI22_X1 U5689 ( .A1(wdata_a_i[3]), .A2(n7467), .B1(n4812), .B2(n9189), .ZN(
        n7465) );
  INV_X1 U5690 ( .A(n7466), .ZN(n8222) );
  AOI22_X1 U5691 ( .A1(wdata_a_i[2]), .A2(n7467), .B1(n4812), .B2(n9191), .ZN(
        n7466) );
  NOR2_X1 U5692 ( .A1(n1581), .A2(n4812), .ZN(n7467) );
  INV_X1 U5693 ( .A(n7468), .ZN(n8223) );
  AOI22_X1 U5694 ( .A1(wdata_a_i[1]), .A2(n7470), .B1(n4812), .B2(n4786), .ZN(
        n7468) );
  INV_X1 U5695 ( .A(n7469), .ZN(n8224) );
  AOI22_X1 U5696 ( .A1(wdata_a_i[0]), .A2(n7470), .B1(n4812), .B2(n9195), .ZN(
        n7469) );
  NOR2_X1 U5697 ( .A1(n1581), .A2(n4812), .ZN(n7470) );
  OR2_X1 U5698 ( .A1(n4812), .A2(n1582), .ZN(n8227) );
  MUX2_X1 U5699 ( .A(wdata_a_i[31]), .B(n4789), .S(n2263), .Z(n8228) );
  MUX2_X1 U5700 ( .A(n4472), .B(n9146), .S(n2263), .Z(n8229) );
  MUX2_X1 U5701 ( .A(n4468), .B(n4803), .S(n2263), .Z(n8230) );
  MUX2_X1 U5702 ( .A(wdata_a_i[28]), .B(wdata_b_i[28]), .S(n2263), .Z(n8231)
         );
  MUX2_X1 U5703 ( .A(n4394), .B(n4732), .S(n2263), .Z(n8232) );
  MUX2_X1 U5704 ( .A(wdata_a_i[26]), .B(n8867), .S(n2263), .Z(n8233) );
  MUX2_X1 U5705 ( .A(wdata_a_i[25]), .B(wdata_b_i[25]), .S(n2263), .Z(n8234)
         );
  MUX2_X1 U5706 ( .A(n4386), .B(n9155), .S(n2263), .Z(n8235) );
  MUX2_X1 U5707 ( .A(wdata_a_i[23]), .B(n9157), .S(n2263), .Z(n8236) );
  MUX2_X1 U5708 ( .A(wdata_a_i[22]), .B(n9159), .S(n2263), .Z(n8237) );
  MUX2_X1 U5709 ( .A(wdata_a_i[21]), .B(n9032), .S(n2263), .Z(n8238) );
  MUX2_X1 U5710 ( .A(wdata_a_i[20]), .B(n9162), .S(n2263), .Z(n8239) );
  MUX2_X1 U5711 ( .A(wdata_a_i[19]), .B(n9164), .S(n2263), .Z(n8240) );
  MUX2_X1 U5712 ( .A(wdata_a_i[18]), .B(n9166), .S(n2263), .Z(n8241) );
  MUX2_X1 U5713 ( .A(wdata_a_i[17]), .B(n9078), .S(n2263), .Z(n8242) );
  MUX2_X1 U5714 ( .A(wdata_a_i[16]), .B(n8349), .S(n2263), .Z(n8243) );
  MUX2_X1 U5715 ( .A(wdata_a_i[15]), .B(n9081), .S(n2263), .Z(n8244) );
  MUX2_X1 U5716 ( .A(wdata_a_i[14]), .B(n9172), .S(n2263), .Z(n8245) );
  MUX2_X1 U5717 ( .A(wdata_a_i[13]), .B(n9174), .S(n2263), .Z(n8246) );
  MUX2_X1 U5718 ( .A(wdata_a_i[12]), .B(n9085), .S(n2263), .Z(n8247) );
  MUX2_X1 U5719 ( .A(wdata_a_i[11]), .B(n4782), .S(n2263), .Z(n8248) );
  MUX2_X1 U5720 ( .A(wdata_a_i[10]), .B(n9178), .S(n2263), .Z(n8249) );
  MUX2_X1 U5721 ( .A(wdata_a_i[9]), .B(n4783), .S(n2263), .Z(n8250) );
  MUX2_X1 U5722 ( .A(wdata_a_i[8]), .B(n8898), .S(n2263), .Z(n8251) );
  MUX2_X1 U5723 ( .A(n4486), .B(n4780), .S(n2263), .Z(n8252) );
  MUX2_X1 U5724 ( .A(wdata_a_i[6]), .B(n9184), .S(n2263), .Z(n8253) );
  MUX2_X1 U5725 ( .A(wdata_a_i[5]), .B(n8902), .S(n2263), .Z(n8254) );
  MUX2_X1 U5726 ( .A(wdata_a_i[4]), .B(n9098), .S(n2263), .Z(n8255) );
  MUX2_X1 U5727 ( .A(wdata_a_i[3]), .B(n8906), .S(n2263), .Z(n8256) );
  MUX2_X1 U5728 ( .A(wdata_a_i[2]), .B(n9191), .S(n2263), .Z(n8257) );
  MUX2_X1 U5729 ( .A(wdata_a_i[1]), .B(n4786), .S(n2263), .Z(n8258) );
  MUX2_X1 U5730 ( .A(wdata_a_i[0]), .B(n4790), .S(n2263), .Z(n8259) );
  NAND2_X1 U5731 ( .A1(n2264), .A2(n7471), .ZN(n8262) );
  INV_X1 U5732 ( .A(n2263), .ZN(n7471) );
  NOR2_X1 U5733 ( .A1(n1541), .A2(n4819), .ZN(n7472) );
  MUX2_X1 U5734 ( .A(n4468), .B(n4803), .S(n4819), .Z(n8265) );
  MUX2_X1 U5735 ( .A(n4618), .B(wdata_b_i[28]), .S(n4819), .Z(n8266) );
  MUX2_X1 U5736 ( .A(n4394), .B(n8865), .S(n4819), .Z(n8267) );
  MUX2_X1 U5737 ( .A(n4459), .B(n9152), .S(n4819), .Z(n8268) );
  MUX2_X1 U5738 ( .A(n4614), .B(wdata_b_i[25]), .S(n4819), .Z(n8269) );
  MUX2_X1 U5739 ( .A(n4386), .B(n9155), .S(n4819), .Z(n8270) );
  NOR2_X1 U5740 ( .A1(n1541), .A2(n4819), .ZN(n7473) );
  NOR2_X1 U5741 ( .A1(n1541), .A2(n4819), .ZN(n7474) );
  NOR2_X1 U5742 ( .A1(n1541), .A2(n4819), .ZN(n7475) );
  MUX2_X1 U5743 ( .A(wdata_a_i[16]), .B(n8349), .S(n4819), .Z(n8278) );
  NOR2_X1 U5744 ( .A1(n1541), .A2(n4819), .ZN(n7476) );
  MUX2_X1 U5745 ( .A(wdata_a_i[14]), .B(n9172), .S(n4819), .Z(n8280) );
  MUX2_X1 U5746 ( .A(wdata_a_i[13]), .B(n9174), .S(n4819), .Z(n8281) );
  MUX2_X1 U5747 ( .A(wdata_a_i[12]), .B(n9085), .S(n4819), .Z(n8282) );
  INV_X1 U5748 ( .A(n7477), .ZN(n8283) );
  AOI22_X1 U5749 ( .A1(wdata_a_i[11]), .A2(n7478), .B1(n4819), .B2(n4782), 
        .ZN(n7477) );
  NOR2_X1 U5750 ( .A1(n1541), .A2(n4819), .ZN(n7478) );
  INV_X1 U5751 ( .A(n7479), .ZN(n8285) );
  AOI22_X1 U5752 ( .A1(wdata_a_i[9]), .A2(n7481), .B1(n4819), .B2(n9091), .ZN(
        n7479) );
  INV_X1 U5753 ( .A(n7480), .ZN(n8286) );
  AOI22_X1 U5754 ( .A1(wdata_a_i[8]), .A2(n7481), .B1(n4819), .B2(n8898), .ZN(
        n7480) );
  NOR2_X1 U5755 ( .A1(n1541), .A2(n4819), .ZN(n7481) );
  INV_X1 U5756 ( .A(n7482), .ZN(n8287) );
  AOI22_X1 U5757 ( .A1(n4486), .A2(n7484), .B1(n4819), .B2(n8848), .ZN(n7482)
         );
  INV_X1 U5758 ( .A(n7483), .ZN(n8288) );
  AOI22_X1 U5759 ( .A1(wdata_a_i[6]), .A2(n7484), .B1(n4819), .B2(n9184), .ZN(
        n7483) );
  NOR2_X1 U5760 ( .A1(n1541), .A2(n4819), .ZN(n7484) );
  INV_X1 U5761 ( .A(n7485), .ZN(n8289) );
  AOI22_X1 U5762 ( .A1(wdata_a_i[5]), .A2(n7487), .B1(n4819), .B2(n8902), .ZN(
        n7485) );
  INV_X1 U5763 ( .A(n7486), .ZN(n8290) );
  AOI22_X1 U5764 ( .A1(wdata_a_i[4]), .A2(n7487), .B1(n4819), .B2(n9098), .ZN(
        n7486) );
  NOR2_X1 U5765 ( .A1(n1541), .A2(n4819), .ZN(n7487) );
  INV_X1 U5766 ( .A(n7488), .ZN(n8291) );
  AOI22_X1 U5767 ( .A1(wdata_a_i[3]), .A2(n7490), .B1(n4819), .B2(n9189), .ZN(
        n7488) );
  INV_X1 U5768 ( .A(n7489), .ZN(n8292) );
  AOI22_X1 U5769 ( .A1(wdata_a_i[2]), .A2(n7490), .B1(n4819), .B2(n9191), .ZN(
        n7489) );
  NOR2_X1 U5770 ( .A1(n1541), .A2(n4819), .ZN(n7490) );
  INV_X1 U5771 ( .A(n7491), .ZN(n8293) );
  AOI22_X1 U5772 ( .A1(wdata_a_i[1]), .A2(n7493), .B1(n4819), .B2(n4786), .ZN(
        n7491) );
  INV_X1 U5773 ( .A(n7492), .ZN(n8294) );
  AOI22_X1 U5774 ( .A1(wdata_a_i[0]), .A2(n7493), .B1(n4819), .B2(n9195), .ZN(
        n7492) );
  NOR2_X1 U5775 ( .A1(n1541), .A2(n4819), .ZN(n7493) );
  OR2_X1 U5776 ( .A1(n1543), .A2(n4819), .ZN(n8297) );
  NOR2_X1 U5777 ( .A1(n1592), .A2(n4746), .ZN(n7494) );
  MUX2_X1 U5778 ( .A(n4468), .B(n4803), .S(n4746), .Z(n8300) );
  MUX2_X1 U5779 ( .A(wdata_a_i[28]), .B(wdata_b_i[28]), .S(n4746), .Z(n8301)
         );
  MUX2_X1 U5780 ( .A(n4394), .B(n8865), .S(n4746), .Z(n8302) );
  MUX2_X1 U5781 ( .A(wdata_a_i[26]), .B(n9152), .S(n4746), .Z(n8303) );
  MUX2_X1 U5782 ( .A(wdata_a_i[25]), .B(wdata_b_i[25]), .S(n4746), .Z(n8304)
         );
  MUX2_X1 U5783 ( .A(n4386), .B(n9155), .S(n4746), .Z(n8305) );
  NOR2_X1 U5784 ( .A1(n1592), .A2(n4746), .ZN(n7495) );
  MUX2_X1 U5785 ( .A(wdata_a_i[21]), .B(n9032), .S(n4746), .Z(n8308) );
  NOR2_X1 U5786 ( .A1(n1592), .A2(n4746), .ZN(n7496) );
  NOR2_X1 U5787 ( .A1(n1592), .A2(n4746), .ZN(n7497) );
  INV_X1 U5788 ( .A(n7498), .ZN(n8313) );
  AOI22_X1 U5789 ( .A1(wdata_a_i[16]), .A2(n7499), .B1(n4746), .B2(n8349), 
        .ZN(n7498) );
  NOR2_X1 U5790 ( .A1(n1592), .A2(n4746), .ZN(n7499) );
  MUX2_X1 U5791 ( .A(wdata_a_i[14]), .B(n9172), .S(n4746), .Z(n8315) );
  MUX2_X1 U5792 ( .A(wdata_a_i[13]), .B(n9174), .S(n4746), .Z(n8316) );
  MUX2_X1 U5793 ( .A(wdata_a_i[12]), .B(n9085), .S(n4746), .Z(n8317) );
  INV_X1 U5794 ( .A(n7500), .ZN(n8318) );
  AOI22_X1 U5795 ( .A1(wdata_a_i[11]), .A2(n7501), .B1(n4746), .B2(n8892), 
        .ZN(n7500) );
  NOR2_X1 U5796 ( .A1(n1592), .A2(n4746), .ZN(n7501) );
  INV_X1 U5797 ( .A(n7502), .ZN(n8320) );
  AOI22_X1 U5798 ( .A1(wdata_a_i[9]), .A2(n7504), .B1(n4746), .B2(n9091), .ZN(
        n7502) );
  INV_X1 U5799 ( .A(n7503), .ZN(n8321) );
  AOI22_X1 U5800 ( .A1(wdata_a_i[8]), .A2(n7504), .B1(n4746), .B2(n4774), .ZN(
        n7503) );
  NOR2_X1 U5801 ( .A1(n1592), .A2(n4746), .ZN(n7504) );
  INV_X1 U5802 ( .A(n7505), .ZN(n8322) );
  AOI22_X1 U5803 ( .A1(n4486), .A2(n7507), .B1(n4746), .B2(n4780), .ZN(n7505)
         );
  INV_X1 U5804 ( .A(n7506), .ZN(n8323) );
  AOI22_X1 U5805 ( .A1(wdata_a_i[6]), .A2(n7507), .B1(n4746), .B2(n9184), .ZN(
        n7506) );
  NOR2_X1 U5806 ( .A1(n1592), .A2(n4746), .ZN(n7507) );
  INV_X1 U5807 ( .A(n7508), .ZN(n8324) );
  AOI22_X1 U5808 ( .A1(wdata_a_i[5]), .A2(n7510), .B1(n9186), .B2(n4746), .ZN(
        n7508) );
  INV_X1 U5809 ( .A(n7509), .ZN(n8325) );
  AOI22_X1 U5810 ( .A1(wdata_a_i[4]), .A2(n7510), .B1(n4746), .B2(n9098), .ZN(
        n7509) );
  NOR2_X1 U5811 ( .A1(n1592), .A2(n4746), .ZN(n7510) );
  INV_X1 U5812 ( .A(n7511), .ZN(n8326) );
  AOI22_X1 U5813 ( .A1(wdata_a_i[3]), .A2(n7513), .B1(n4746), .B2(n9189), .ZN(
        n7511) );
  INV_X1 U5814 ( .A(n7512), .ZN(n8327) );
  AOI22_X1 U5815 ( .A1(wdata_a_i[2]), .A2(n7513), .B1(n4746), .B2(n9191), .ZN(
        n7512) );
  NOR2_X1 U5816 ( .A1(n1592), .A2(n4746), .ZN(n7513) );
  INV_X1 U5817 ( .A(n7514), .ZN(n8328) );
  AOI22_X1 U5818 ( .A1(wdata_a_i[1]), .A2(n7516), .B1(n4746), .B2(n9193), .ZN(
        n7514) );
  INV_X1 U5819 ( .A(n7515), .ZN(n8329) );
  AOI22_X1 U5820 ( .A1(wdata_a_i[0]), .A2(n7516), .B1(n4746), .B2(n9195), .ZN(
        n7515) );
  NOR2_X1 U5821 ( .A1(n1592), .A2(n4746), .ZN(n7516) );
  OR2_X1 U5822 ( .A1(n4746), .A2(n1593), .ZN(n8332) );
  NOR2_X1 U5823 ( .A1(n1537), .A2(n4817), .ZN(n7517) );
  MUX2_X1 U5824 ( .A(n4468), .B(n4803), .S(n4817), .Z(n8335) );
  MUX2_X1 U5825 ( .A(n4618), .B(wdata_b_i[28]), .S(n4817), .Z(n8336) );
  MUX2_X1 U5826 ( .A(n4394), .B(n4732), .S(n4817), .Z(n8337) );
  MUX2_X1 U5827 ( .A(n4459), .B(n8867), .S(n4817), .Z(n8338) );
  MUX2_X1 U5828 ( .A(n4614), .B(wdata_b_i[25]), .S(n4817), .Z(n8339) );
  MUX2_X1 U5829 ( .A(n4386), .B(n9155), .S(n4817), .Z(n8340) );
  NOR2_X1 U5830 ( .A1(n1537), .A2(n4817), .ZN(n7518) );
  NOR2_X1 U5831 ( .A1(n1537), .A2(n4817), .ZN(n7519) );
  NOR2_X1 U5832 ( .A1(n1537), .A2(n4817), .ZN(n7520) );
  MUX2_X1 U5833 ( .A(wdata_a_i[16]), .B(n8349), .S(n4817), .Z(n8348) );
  NOR2_X1 U5834 ( .A1(n1537), .A2(n4817), .ZN(n7521) );
  MUX2_X1 U5835 ( .A(wdata_a_i[14]), .B(n9172), .S(n4817), .Z(n8351) );
  MUX2_X1 U5836 ( .A(wdata_a_i[13]), .B(n9174), .S(n4817), .Z(n8352) );
  MUX2_X1 U5837 ( .A(wdata_a_i[12]), .B(n9085), .S(n4817), .Z(n8353) );
  INV_X1 U5838 ( .A(n7522), .ZN(n8354) );
  AOI22_X1 U5839 ( .A1(wdata_a_i[11]), .A2(n7523), .B1(n4817), .B2(n4782), 
        .ZN(n7522) );
  NOR2_X1 U5840 ( .A1(n1537), .A2(n4817), .ZN(n7523) );
  INV_X1 U5841 ( .A(n7524), .ZN(n8356) );
  AOI22_X1 U5842 ( .A1(wdata_a_i[9]), .A2(n7526), .B1(n4817), .B2(n9091), .ZN(
        n7524) );
  INV_X1 U5843 ( .A(n7525), .ZN(n8357) );
  AOI22_X1 U5844 ( .A1(wdata_a_i[8]), .A2(n7526), .B1(n4817), .B2(n8898), .ZN(
        n7525) );
  NOR2_X1 U5845 ( .A1(n1537), .A2(n4817), .ZN(n7526) );
  INV_X1 U5846 ( .A(n7527), .ZN(n8358) );
  AOI22_X1 U5847 ( .A1(n4486), .A2(n7529), .B1(n4817), .B2(n4779), .ZN(n7527)
         );
  INV_X1 U5848 ( .A(n7528), .ZN(n8359) );
  AOI22_X1 U5849 ( .A1(wdata_a_i[6]), .A2(n7529), .B1(n4817), .B2(n9184), .ZN(
        n7528) );
  NOR2_X1 U5850 ( .A1(n1537), .A2(n4817), .ZN(n7529) );
  INV_X1 U5851 ( .A(n7530), .ZN(n8360) );
  AOI22_X1 U5852 ( .A1(wdata_a_i[5]), .A2(n7532), .B1(n4817), .B2(n9096), .ZN(
        n7530) );
  INV_X1 U5853 ( .A(n7531), .ZN(n8361) );
  AOI22_X1 U5854 ( .A1(wdata_a_i[4]), .A2(n7532), .B1(n4817), .B2(n4787), .ZN(
        n7531) );
  NOR2_X1 U5855 ( .A1(n1537), .A2(n4817), .ZN(n7532) );
  INV_X1 U5856 ( .A(n7533), .ZN(n8362) );
  AOI22_X1 U5857 ( .A1(wdata_a_i[3]), .A2(n7535), .B1(n4817), .B2(n9189), .ZN(
        n7533) );
  INV_X1 U5858 ( .A(n7534), .ZN(n8363) );
  AOI22_X1 U5859 ( .A1(wdata_a_i[2]), .A2(n7535), .B1(n4817), .B2(n9191), .ZN(
        n7534) );
  NOR2_X1 U5860 ( .A1(n1537), .A2(n4817), .ZN(n7535) );
  INV_X1 U5861 ( .A(n7536), .ZN(n8364) );
  AOI22_X1 U5862 ( .A1(wdata_a_i[1]), .A2(n7538), .B1(n4817), .B2(n4786), .ZN(
        n7536) );
  INV_X1 U5863 ( .A(n7537), .ZN(n8365) );
  AOI22_X1 U5864 ( .A1(wdata_a_i[0]), .A2(n7538), .B1(n4817), .B2(n9195), .ZN(
        n7537) );
  NOR2_X1 U5865 ( .A1(n1537), .A2(n4817), .ZN(n7538) );
  OR2_X1 U5866 ( .A1(n1539), .A2(n4817), .ZN(n8368) );
  NOR2_X1 U5867 ( .A1(n1597), .A2(n4807), .ZN(n7539) );
  MUX2_X1 U5868 ( .A(n4468), .B(n4803), .S(n4807), .Z(n8371) );
  MUX2_X1 U5869 ( .A(n4618), .B(wdata_b_i[28]), .S(n4807), .Z(n8372) );
  MUX2_X1 U5870 ( .A(n4394), .B(n8865), .S(n4807), .Z(n8373) );
  MUX2_X1 U5871 ( .A(n4459), .B(n9152), .S(n4807), .Z(n8374) );
  MUX2_X1 U5872 ( .A(n4614), .B(wdata_b_i[25]), .S(n4807), .Z(n8375) );
  MUX2_X1 U5873 ( .A(n4386), .B(n9155), .S(n4807), .Z(n8376) );
  NOR2_X1 U5874 ( .A1(n1597), .A2(n4807), .ZN(n7540) );
  MUX2_X1 U5875 ( .A(wdata_a_i[21]), .B(n9032), .S(n4807), .Z(n8379) );
  NOR2_X1 U5876 ( .A1(n1597), .A2(n4807), .ZN(n7541) );
  NOR2_X1 U5877 ( .A1(n1597), .A2(n4807), .ZN(n7542) );
  INV_X1 U5878 ( .A(n7543), .ZN(n8384) );
  AOI22_X1 U5879 ( .A1(wdata_a_i[16]), .A2(n7544), .B1(n4807), .B2(n8349), 
        .ZN(n7543) );
  NOR2_X1 U5880 ( .A1(n1597), .A2(n4807), .ZN(n7544) );
  MUX2_X1 U5881 ( .A(wdata_a_i[14]), .B(n9172), .S(n4807), .Z(n8386) );
  MUX2_X1 U5882 ( .A(wdata_a_i[13]), .B(n9174), .S(n4807), .Z(n8387) );
  MUX2_X1 U5883 ( .A(wdata_a_i[12]), .B(n9085), .S(n4807), .Z(n8388) );
  INV_X1 U5884 ( .A(n7545), .ZN(n8389) );
  AOI22_X1 U5885 ( .A1(wdata_a_i[11]), .A2(n7546), .B1(n4807), .B2(n4782), 
        .ZN(n7545) );
  NOR2_X1 U5886 ( .A1(n1597), .A2(n4807), .ZN(n7546) );
  INV_X1 U5887 ( .A(n7547), .ZN(n8391) );
  AOI22_X1 U5888 ( .A1(wdata_a_i[9]), .A2(n7549), .B1(n4807), .B2(n9091), .ZN(
        n7547) );
  INV_X1 U5889 ( .A(n7548), .ZN(n8392) );
  AOI22_X1 U5890 ( .A1(wdata_a_i[8]), .A2(n7549), .B1(n4807), .B2(n8898), .ZN(
        n7548) );
  NOR2_X1 U5891 ( .A1(n1597), .A2(n4807), .ZN(n7549) );
  INV_X1 U5892 ( .A(n7550), .ZN(n8393) );
  AOI22_X1 U5893 ( .A1(wdata_a_i[7]), .A2(n7552), .B1(n4807), .B2(n8848), .ZN(
        n7550) );
  INV_X1 U5894 ( .A(n7551), .ZN(n8394) );
  AOI22_X1 U5895 ( .A1(wdata_a_i[6]), .A2(n7552), .B1(n4807), .B2(n9184), .ZN(
        n7551) );
  NOR2_X1 U5896 ( .A1(n1597), .A2(n4807), .ZN(n7552) );
  INV_X1 U5897 ( .A(n7553), .ZN(n8395) );
  AOI22_X1 U5898 ( .A1(wdata_a_i[5]), .A2(n7555), .B1(n4807), .B2(n8902), .ZN(
        n7553) );
  INV_X1 U5899 ( .A(n7554), .ZN(n8396) );
  AOI22_X1 U5900 ( .A1(wdata_a_i[4]), .A2(n7555), .B1(n4807), .B2(n9098), .ZN(
        n7554) );
  NOR2_X1 U5901 ( .A1(n1597), .A2(n4807), .ZN(n7555) );
  INV_X1 U5902 ( .A(n7556), .ZN(n8397) );
  AOI22_X1 U5903 ( .A1(wdata_a_i[3]), .A2(n7558), .B1(n4807), .B2(n9189), .ZN(
        n7556) );
  INV_X1 U5904 ( .A(n7557), .ZN(n8398) );
  AOI22_X1 U5905 ( .A1(wdata_a_i[2]), .A2(n7558), .B1(n4807), .B2(n9191), .ZN(
        n7557) );
  NOR2_X1 U5906 ( .A1(n1597), .A2(n4807), .ZN(n7558) );
  INV_X1 U5907 ( .A(n7559), .ZN(n8399) );
  AOI22_X1 U5908 ( .A1(wdata_a_i[1]), .A2(n7561), .B1(n4807), .B2(n4786), .ZN(
        n7559) );
  INV_X1 U5909 ( .A(n7560), .ZN(n8400) );
  AOI22_X1 U5910 ( .A1(wdata_a_i[0]), .A2(n7561), .B1(n4807), .B2(n9195), .ZN(
        n7560) );
  NOR2_X1 U5911 ( .A1(n1597), .A2(n4807), .ZN(n7561) );
  OR2_X1 U5912 ( .A1(n4807), .A2(n1598), .ZN(n8403) );
  NOR2_X1 U5913 ( .A1(n2481), .A2(n4745), .ZN(n7562) );
  INV_X1 U5914 ( .A(n7563), .ZN(n8407) );
  AOI22_X1 U5915 ( .A1(wdata_a_i[28]), .A2(n7564), .B1(n4745), .B2(
        wdata_b_i[28]), .ZN(n7563) );
  NOR2_X1 U5916 ( .A1(n2481), .A2(n4745), .ZN(n7564) );
  INV_X1 U5917 ( .A(n7565), .ZN(n8408) );
  AOI22_X1 U5918 ( .A1(wdata_a_i[27]), .A2(n7567), .B1(n4745), .B2(n8865), 
        .ZN(n7565) );
  INV_X1 U5919 ( .A(n7566), .ZN(n8409) );
  AOI22_X1 U5920 ( .A1(wdata_a_i[26]), .A2(n7567), .B1(n4745), .B2(n9063), 
        .ZN(n7566) );
  NOR2_X1 U5921 ( .A1(n2481), .A2(n4745), .ZN(n7567) );
  INV_X1 U5922 ( .A(n7568), .ZN(n8410) );
  AOI22_X1 U5923 ( .A1(wdata_a_i[25]), .A2(n7570), .B1(n4745), .B2(
        wdata_b_i[25]), .ZN(n7568) );
  INV_X1 U5924 ( .A(n7569), .ZN(n8411) );
  AOI22_X1 U5925 ( .A1(wdata_a_i[24]), .A2(n7570), .B1(n4745), .B2(n8923), 
        .ZN(n7569) );
  NOR2_X1 U5926 ( .A1(n2481), .A2(n4745), .ZN(n7570) );
  NOR2_X1 U5927 ( .A1(n2481), .A2(n4745), .ZN(n7571) );
  NOR2_X1 U5928 ( .A1(n2481), .A2(n4745), .ZN(n7572) );
  NOR2_X1 U5929 ( .A1(n2481), .A2(n4745), .ZN(n7573) );
  INV_X1 U5930 ( .A(n7574), .ZN(n8419) );
  AOI22_X1 U5931 ( .A1(wdata_a_i[16]), .A2(n7575), .B1(n4745), .B2(n8349), 
        .ZN(n7574) );
  NOR2_X1 U5932 ( .A1(n2481), .A2(n4745), .ZN(n7575) );
  MUX2_X1 U5933 ( .A(wdata_a_i[14]), .B(n8887), .S(n4745), .Z(n8421) );
  MUX2_X1 U5934 ( .A(wdata_a_i[13]), .B(n9174), .S(n4745), .Z(n8422) );
  MUX2_X1 U5935 ( .A(wdata_a_i[12]), .B(n9085), .S(n4745), .Z(n8423) );
  MUX2_X1 U5936 ( .A(wdata_a_i[11]), .B(n9087), .S(n4745), .Z(n8424) );
  MUX2_X1 U5937 ( .A(wdata_a_i[10]), .B(n9089), .S(n4745), .Z(n8425) );
  MUX2_X1 U5938 ( .A(wdata_a_i[9]), .B(n4783), .S(n4745), .Z(n8426) );
  MUX2_X1 U5939 ( .A(wdata_a_i[8]), .B(n4774), .S(n4745), .Z(n8427) );
  MUX2_X1 U5940 ( .A(wdata_a_i[7]), .B(wdata_b_i[7]), .S(n4745), .Z(n8428) );
  MUX2_X1 U5941 ( .A(wdata_a_i[6]), .B(n4420), .S(n4745), .Z(n8429) );
  INV_X1 U5942 ( .A(n7576), .ZN(n8430) );
  AOI22_X1 U5943 ( .A1(wdata_a_i[5]), .A2(n7577), .B1(n8902), .B2(n4745), .ZN(
        n7576) );
  NOR2_X1 U5944 ( .A1(n2481), .A2(n4745), .ZN(n7577) );
  INV_X1 U5945 ( .A(n7578), .ZN(n8431) );
  AOI22_X1 U5946 ( .A1(wdata_a_i[4]), .A2(n7580), .B1(n4745), .B2(n9098), .ZN(
        n7578) );
  MUX2_X1 U5947 ( .A(wdata_a_i[3]), .B(n9100), .S(n4745), .Z(n8432) );
  INV_X1 U5948 ( .A(n7579), .ZN(n8433) );
  AOI22_X1 U5949 ( .A1(wdata_a_i[2]), .A2(n7580), .B1(n4745), .B2(n9102), .ZN(
        n7579) );
  NOR2_X1 U5950 ( .A1(n2481), .A2(n4745), .ZN(n7580) );
  INV_X1 U5951 ( .A(n7581), .ZN(n8434) );
  AOI22_X1 U5952 ( .A1(wdata_a_i[1]), .A2(n7583), .B1(n4745), .B2(n9104), .ZN(
        n7581) );
  INV_X1 U5953 ( .A(n7582), .ZN(n8435) );
  AOI22_X1 U5954 ( .A1(wdata_a_i[0]), .A2(n7583), .B1(n4745), .B2(n4791), .ZN(
        n7582) );
  NOR2_X1 U5955 ( .A1(n2481), .A2(n4745), .ZN(n7583) );
  NAND2_X1 U5956 ( .A1(n2481), .A2(n4747), .ZN(n8438) );
  NOR2_X1 U5957 ( .A1(n1561), .A2(n4810), .ZN(n7584) );
  MUX2_X1 U5958 ( .A(n4468), .B(n4796), .S(n4810), .Z(n8441) );
  MUX2_X1 U5959 ( .A(n4618), .B(wdata_b_i[28]), .S(n4810), .Z(n8442) );
  MUX2_X1 U5960 ( .A(wdata_a_i[27]), .B(n4732), .S(n4810), .Z(n8443) );
  MUX2_X1 U5961 ( .A(n4459), .B(n8867), .S(n4810), .Z(n8444) );
  MUX2_X1 U5962 ( .A(n4614), .B(wdata_b_i[25]), .S(n4810), .Z(n8445) );
  MUX2_X1 U5963 ( .A(n4386), .B(n8923), .S(n4810), .Z(n8446) );
  NOR2_X1 U5964 ( .A1(n1561), .A2(n4810), .ZN(n7585) );
  MUX2_X1 U5965 ( .A(wdata_a_i[21]), .B(n9032), .S(n4810), .Z(n8449) );
  NOR2_X1 U5966 ( .A1(n1561), .A2(n4810), .ZN(n7586) );
  NOR2_X1 U5967 ( .A1(n1561), .A2(n4810), .ZN(n7587) );
  INV_X1 U5968 ( .A(n7588), .ZN(n8454) );
  AOI22_X1 U5969 ( .A1(wdata_a_i[16]), .A2(n7590), .B1(n4810), .B2(n8883), 
        .ZN(n7588) );
  INV_X1 U5970 ( .A(n7589), .ZN(n8455) );
  AOI22_X1 U5971 ( .A1(wdata_a_i[15]), .A2(n7590), .B1(n4810), .B2(n8885), 
        .ZN(n7589) );
  NOR2_X1 U5972 ( .A1(n1561), .A2(n4810), .ZN(n7590) );
  MUX2_X1 U5973 ( .A(wdata_a_i[14]), .B(n8887), .S(n4810), .Z(n8456) );
  MUX2_X1 U5974 ( .A(wdata_a_i[13]), .B(wdata_b_i[13]), .S(n4810), .Z(n8457)
         );
  MUX2_X1 U5975 ( .A(wdata_a_i[12]), .B(n8890), .S(n4810), .Z(n8458) );
  INV_X1 U5976 ( .A(n7591), .ZN(n8459) );
  AOI22_X1 U5977 ( .A1(wdata_a_i[11]), .A2(n7592), .B1(n4810), .B2(n8892), 
        .ZN(n7591) );
  NOR2_X1 U5978 ( .A1(n1561), .A2(n4810), .ZN(n7592) );
  INV_X1 U5979 ( .A(n7593), .ZN(n8461) );
  AOI22_X1 U5980 ( .A1(wdata_a_i[9]), .A2(n7595), .B1(n4810), .B2(n8896), .ZN(
        n7593) );
  INV_X1 U5981 ( .A(n7594), .ZN(n8462) );
  AOI22_X1 U5982 ( .A1(wdata_a_i[8]), .A2(n7595), .B1(n4810), .B2(wdata_b_i[8]), .ZN(n7594) );
  NOR2_X1 U5983 ( .A1(n1561), .A2(n4810), .ZN(n7595) );
  INV_X1 U5984 ( .A(n7596), .ZN(n8463) );
  AOI22_X1 U5985 ( .A1(n4486), .A2(n7598), .B1(n4810), .B2(n8848), .ZN(n7596)
         );
  INV_X1 U5986 ( .A(n7597), .ZN(n8464) );
  AOI22_X1 U5987 ( .A1(wdata_a_i[6]), .A2(n7598), .B1(n4810), .B2(n4420), .ZN(
        n7597) );
  NOR2_X1 U5988 ( .A1(n1561), .A2(n4810), .ZN(n7598) );
  INV_X1 U5989 ( .A(n7599), .ZN(n8465) );
  AOI22_X1 U5990 ( .A1(wdata_a_i[5]), .A2(n7601), .B1(n4810), .B2(n9186), .ZN(
        n7599) );
  INV_X1 U5991 ( .A(n7600), .ZN(n8466) );
  AOI22_X1 U5992 ( .A1(wdata_a_i[4]), .A2(n7601), .B1(n4810), .B2(n8904), .ZN(
        n7600) );
  NOR2_X1 U5993 ( .A1(n1561), .A2(n4810), .ZN(n7601) );
  INV_X1 U5994 ( .A(n7602), .ZN(n8467) );
  AOI22_X1 U5995 ( .A1(wdata_a_i[3]), .A2(n7604), .B1(n4810), .B2(n8906), .ZN(
        n7602) );
  INV_X1 U5996 ( .A(n7603), .ZN(n8468) );
  AOI22_X1 U5997 ( .A1(wdata_a_i[2]), .A2(n7604), .B1(n4810), .B2(n8908), .ZN(
        n7603) );
  NOR2_X1 U5998 ( .A1(n1561), .A2(n4810), .ZN(n7604) );
  INV_X1 U5999 ( .A(n7605), .ZN(n8469) );
  AOI22_X1 U6000 ( .A1(wdata_a_i[1]), .A2(n7607), .B1(n4810), .B2(n8910), .ZN(
        n7605) );
  INV_X1 U6001 ( .A(n7606), .ZN(n8470) );
  AOI22_X1 U6002 ( .A1(wdata_a_i[0]), .A2(n7607), .B1(n4810), .B2(n9195), .ZN(
        n7606) );
  NOR2_X1 U6003 ( .A1(n1561), .A2(n4810), .ZN(n7607) );
  OR2_X1 U6004 ( .A1(n1563), .A2(n4810), .ZN(n8473) );
  NOR2_X1 U6005 ( .A1(n1555), .A2(n4808), .ZN(n7608) );
  MUX2_X1 U6006 ( .A(n4468), .B(n4796), .S(n4808), .Z(n8476) );
  MUX2_X1 U6007 ( .A(n4618), .B(wdata_b_i[28]), .S(n4808), .Z(n8477) );
  MUX2_X1 U6008 ( .A(wdata_a_i[27]), .B(n8865), .S(n4808), .Z(n8478) );
  MUX2_X1 U6009 ( .A(n4459), .B(n9152), .S(n4808), .Z(n8479) );
  MUX2_X1 U6010 ( .A(n4614), .B(wdata_b_i[25]), .S(n4808), .Z(n8480) );
  MUX2_X1 U6011 ( .A(wdata_a_i[24]), .B(n8923), .S(n4808), .Z(n8481) );
  NOR2_X1 U6012 ( .A1(n1555), .A2(n4808), .ZN(n7609) );
  NOR2_X1 U6013 ( .A1(n1555), .A2(n4808), .ZN(n7610) );
  NOR2_X1 U6014 ( .A1(n1555), .A2(n4808), .ZN(n7611) );
  MUX2_X1 U6015 ( .A(wdata_a_i[16]), .B(n4734), .S(n4808), .Z(n8489) );
  INV_X1 U6016 ( .A(n7612), .ZN(n8490) );
  AOI22_X1 U6017 ( .A1(wdata_a_i[15]), .A2(n7613), .B1(n4808), .B2(n9081), 
        .ZN(n7612) );
  NOR2_X1 U6018 ( .A1(n1555), .A2(n4808), .ZN(n7613) );
  MUX2_X1 U6019 ( .A(wdata_a_i[14]), .B(n8887), .S(n4808), .Z(n8491) );
  MUX2_X1 U6020 ( .A(wdata_a_i[13]), .B(wdata_b_i[13]), .S(n4808), .Z(n8492)
         );
  MUX2_X1 U6021 ( .A(wdata_a_i[12]), .B(n8890), .S(n4808), .Z(n8493) );
  INV_X1 U6022 ( .A(n7614), .ZN(n8494) );
  AOI22_X1 U6023 ( .A1(wdata_a_i[11]), .A2(n7615), .B1(n4808), .B2(n8892), 
        .ZN(n7614) );
  NOR2_X1 U6024 ( .A1(n1555), .A2(n4808), .ZN(n7615) );
  INV_X1 U6025 ( .A(n7616), .ZN(n8496) );
  AOI22_X1 U6026 ( .A1(wdata_a_i[9]), .A2(n7618), .B1(n4808), .B2(n9091), .ZN(
        n7616) );
  INV_X1 U6027 ( .A(n7617), .ZN(n8497) );
  AOI22_X1 U6028 ( .A1(wdata_a_i[8]), .A2(n7618), .B1(n4808), .B2(wdata_b_i[8]), .ZN(n7617) );
  NOR2_X1 U6029 ( .A1(n1555), .A2(n4808), .ZN(n7618) );
  INV_X1 U6030 ( .A(n7619), .ZN(n8498) );
  AOI22_X1 U6031 ( .A1(n4486), .A2(n7621), .B1(n4808), .B2(n9182), .ZN(n7619)
         );
  INV_X1 U6032 ( .A(n7620), .ZN(n8499) );
  AOI22_X1 U6033 ( .A1(wdata_a_i[6]), .A2(n7621), .B1(n4808), .B2(n4420), .ZN(
        n7620) );
  NOR2_X1 U6034 ( .A1(n1555), .A2(n4808), .ZN(n7621) );
  INV_X1 U6035 ( .A(n7622), .ZN(n8500) );
  AOI22_X1 U6036 ( .A1(wdata_a_i[5]), .A2(n7624), .B1(n4808), .B2(n9186), .ZN(
        n7622) );
  INV_X1 U6037 ( .A(n7623), .ZN(n8501) );
  AOI22_X1 U6038 ( .A1(wdata_a_i[4]), .A2(n7624), .B1(n4808), .B2(n8904), .ZN(
        n7623) );
  NOR2_X1 U6039 ( .A1(n1555), .A2(n4808), .ZN(n7624) );
  INV_X1 U6040 ( .A(n7625), .ZN(n8502) );
  AOI22_X1 U6041 ( .A1(wdata_a_i[3]), .A2(n7627), .B1(n4808), .B2(n8906), .ZN(
        n7625) );
  INV_X1 U6042 ( .A(n7626), .ZN(n8503) );
  AOI22_X1 U6043 ( .A1(wdata_a_i[2]), .A2(n7627), .B1(n4808), .B2(n8908), .ZN(
        n7626) );
  NOR2_X1 U6044 ( .A1(n1555), .A2(n4808), .ZN(n7627) );
  INV_X1 U6045 ( .A(n7628), .ZN(n8504) );
  AOI22_X1 U6046 ( .A1(wdata_a_i[1]), .A2(n7630), .B1(n4808), .B2(n8910), .ZN(
        n7628) );
  INV_X1 U6047 ( .A(n7629), .ZN(n8505) );
  AOI22_X1 U6048 ( .A1(wdata_a_i[0]), .A2(n7630), .B1(n4808), .B2(n4790), .ZN(
        n7629) );
  NOR2_X1 U6049 ( .A1(n1555), .A2(n4808), .ZN(n7630) );
  OR2_X1 U6050 ( .A1(n4808), .A2(n1556), .ZN(n8508) );
  NOR2_X1 U6051 ( .A1(n1566), .A2(n4811), .ZN(n7631) );
  MUX2_X1 U6052 ( .A(n4468), .B(n4796), .S(n4811), .Z(n8511) );
  MUX2_X1 U6053 ( .A(n4618), .B(wdata_b_i[28]), .S(n4811), .Z(n8512) );
  MUX2_X1 U6054 ( .A(wdata_a_i[27]), .B(n4732), .S(n4811), .Z(n8513) );
  MUX2_X1 U6055 ( .A(n4459), .B(n8867), .S(n4811), .Z(n8514) );
  MUX2_X1 U6056 ( .A(n4614), .B(wdata_b_i[25]), .S(n4811), .Z(n8515) );
  MUX2_X1 U6057 ( .A(wdata_a_i[24]), .B(n8923), .S(n4811), .Z(n8516) );
  NOR2_X1 U6058 ( .A1(n1566), .A2(n4811), .ZN(n7632) );
  MUX2_X1 U6059 ( .A(wdata_a_i[21]), .B(n9032), .S(n4811), .Z(n8519) );
  NOR2_X1 U6060 ( .A1(n1566), .A2(n4811), .ZN(n7633) );
  NOR2_X1 U6061 ( .A1(n1566), .A2(n4811), .ZN(n7634) );
  INV_X1 U6062 ( .A(n7635), .ZN(n8524) );
  AOI22_X1 U6063 ( .A1(wdata_a_i[16]), .A2(n7637), .B1(n4811), .B2(n8883), 
        .ZN(n7635) );
  INV_X1 U6064 ( .A(n7636), .ZN(n8525) );
  AOI22_X1 U6065 ( .A1(wdata_a_i[15]), .A2(n7637), .B1(n4811), .B2(n8885), 
        .ZN(n7636) );
  NOR2_X1 U6066 ( .A1(n1566), .A2(n4811), .ZN(n7637) );
  MUX2_X1 U6067 ( .A(wdata_a_i[14]), .B(n8887), .S(n4811), .Z(n8526) );
  MUX2_X1 U6068 ( .A(wdata_a_i[13]), .B(wdata_b_i[13]), .S(n4811), .Z(n8527)
         );
  MUX2_X1 U6069 ( .A(wdata_a_i[12]), .B(n8890), .S(n4811), .Z(n8528) );
  INV_X1 U6070 ( .A(n7638), .ZN(n8529) );
  AOI22_X1 U6071 ( .A1(wdata_a_i[11]), .A2(n7639), .B1(n4811), .B2(n8892), 
        .ZN(n7638) );
  NOR2_X1 U6072 ( .A1(n1566), .A2(n4811), .ZN(n7639) );
  INV_X1 U6073 ( .A(n7640), .ZN(n8531) );
  AOI22_X1 U6074 ( .A1(wdata_a_i[9]), .A2(n7642), .B1(n4811), .B2(n9091), .ZN(
        n7640) );
  INV_X1 U6075 ( .A(n7641), .ZN(n8532) );
  AOI22_X1 U6076 ( .A1(wdata_a_i[8]), .A2(n7642), .B1(n4811), .B2(wdata_b_i[8]), .ZN(n7641) );
  NOR2_X1 U6077 ( .A1(n1566), .A2(n4811), .ZN(n7642) );
  INV_X1 U6078 ( .A(n7643), .ZN(n8533) );
  AOI22_X1 U6079 ( .A1(n4486), .A2(n7645), .B1(n4811), .B2(n9182), .ZN(n7643)
         );
  INV_X1 U6080 ( .A(n7644), .ZN(n8534) );
  AOI22_X1 U6081 ( .A1(wdata_a_i[6]), .A2(n7645), .B1(n4811), .B2(n4420), .ZN(
        n7644) );
  NOR2_X1 U6082 ( .A1(n1566), .A2(n4811), .ZN(n7645) );
  INV_X1 U6083 ( .A(n7646), .ZN(n8535) );
  AOI22_X1 U6084 ( .A1(wdata_a_i[5]), .A2(n7648), .B1(n4811), .B2(n9186), .ZN(
        n7646) );
  INV_X1 U6085 ( .A(n7647), .ZN(n8536) );
  AOI22_X1 U6086 ( .A1(wdata_a_i[4]), .A2(n7648), .B1(n4811), .B2(n8904), .ZN(
        n7647) );
  NOR2_X1 U6087 ( .A1(n1566), .A2(n4811), .ZN(n7648) );
  INV_X1 U6088 ( .A(n7649), .ZN(n8537) );
  AOI22_X1 U6089 ( .A1(wdata_a_i[3]), .A2(n7651), .B1(n4811), .B2(n9100), .ZN(
        n7649) );
  INV_X1 U6090 ( .A(n7650), .ZN(n8538) );
  AOI22_X1 U6091 ( .A1(wdata_a_i[2]), .A2(n7651), .B1(n4811), .B2(n8908), .ZN(
        n7650) );
  NOR2_X1 U6092 ( .A1(n1566), .A2(n4811), .ZN(n7651) );
  INV_X1 U6093 ( .A(n7652), .ZN(n8539) );
  AOI22_X1 U6094 ( .A1(wdata_a_i[1]), .A2(n7654), .B1(n4811), .B2(n8910), .ZN(
        n7652) );
  INV_X1 U6095 ( .A(n7653), .ZN(n8540) );
  AOI22_X1 U6096 ( .A1(wdata_a_i[0]), .A2(n7654), .B1(n4811), .B2(n4790), .ZN(
        n7653) );
  NOR2_X1 U6097 ( .A1(n1566), .A2(n4811), .ZN(n7654) );
  OR2_X1 U6098 ( .A1(n1568), .A2(n4811), .ZN(n8543) );
  NOR2_X1 U6099 ( .A1(n1610), .A2(n4809), .ZN(n7655) );
  MUX2_X1 U6100 ( .A(n4468), .B(n4796), .S(n4809), .Z(n8546) );
  MUX2_X1 U6101 ( .A(n4618), .B(wdata_b_i[28]), .S(n4809), .Z(n8547) );
  MUX2_X1 U6102 ( .A(n4394), .B(n8865), .S(n4809), .Z(n8548) );
  MUX2_X1 U6103 ( .A(n4459), .B(n9152), .S(n4809), .Z(n8549) );
  MUX2_X1 U6104 ( .A(n4614), .B(wdata_b_i[25]), .S(n4809), .Z(n8550) );
  MUX2_X1 U6105 ( .A(wdata_a_i[24]), .B(n8923), .S(n4809), .Z(n8551) );
  NOR2_X1 U6106 ( .A1(n1610), .A2(n4809), .ZN(n7656) );
  NOR2_X1 U6107 ( .A1(n1610), .A2(n4809), .ZN(n7657) );
  NOR2_X1 U6108 ( .A1(n1610), .A2(n4809), .ZN(n7658) );
  MUX2_X1 U6109 ( .A(wdata_a_i[16]), .B(n4734), .S(n4809), .Z(n8559) );
  INV_X1 U6110 ( .A(n7659), .ZN(n8560) );
  AOI22_X1 U6111 ( .A1(wdata_a_i[15]), .A2(n7660), .B1(n4809), .B2(n9081), 
        .ZN(n7659) );
  NOR2_X1 U6112 ( .A1(n1610), .A2(n4809), .ZN(n7660) );
  MUX2_X1 U6113 ( .A(wdata_a_i[14]), .B(n8887), .S(n4809), .Z(n8561) );
  MUX2_X1 U6114 ( .A(wdata_a_i[13]), .B(wdata_b_i[13]), .S(n4809), .Z(n8562)
         );
  MUX2_X1 U6115 ( .A(wdata_a_i[12]), .B(n8890), .S(n4809), .Z(n8563) );
  INV_X1 U6116 ( .A(n7661), .ZN(n8564) );
  AOI22_X1 U6117 ( .A1(wdata_a_i[11]), .A2(n7662), .B1(n4809), .B2(n8892), 
        .ZN(n7661) );
  NOR2_X1 U6118 ( .A1(n1610), .A2(n4809), .ZN(n7662) );
  INV_X1 U6119 ( .A(n7663), .ZN(n8566) );
  AOI22_X1 U6120 ( .A1(wdata_a_i[9]), .A2(n7665), .B1(n4809), .B2(n9091), .ZN(
        n7663) );
  INV_X1 U6121 ( .A(n7664), .ZN(n8567) );
  AOI22_X1 U6122 ( .A1(wdata_a_i[8]), .A2(n7665), .B1(n4809), .B2(wdata_b_i[8]), .ZN(n7664) );
  NOR2_X1 U6123 ( .A1(n1610), .A2(n4809), .ZN(n7665) );
  INV_X1 U6124 ( .A(n7666), .ZN(n8568) );
  AOI22_X1 U6125 ( .A1(n4486), .A2(n7668), .B1(n4809), .B2(n9182), .ZN(n7666)
         );
  INV_X1 U6126 ( .A(n7667), .ZN(n8569) );
  AOI22_X1 U6127 ( .A1(wdata_a_i[6]), .A2(n7668), .B1(n4809), .B2(n4420), .ZN(
        n7667) );
  NOR2_X1 U6128 ( .A1(n1610), .A2(n4809), .ZN(n7668) );
  INV_X1 U6129 ( .A(n7669), .ZN(n8570) );
  AOI22_X1 U6130 ( .A1(wdata_a_i[5]), .A2(n7671), .B1(n4809), .B2(n9186), .ZN(
        n7669) );
  INV_X1 U6131 ( .A(n7670), .ZN(n8571) );
  AOI22_X1 U6132 ( .A1(wdata_a_i[4]), .A2(n7671), .B1(n4809), .B2(n4787), .ZN(
        n7670) );
  NOR2_X1 U6133 ( .A1(n1610), .A2(n4809), .ZN(n7671) );
  INV_X1 U6134 ( .A(n7672), .ZN(n8572) );
  AOI22_X1 U6135 ( .A1(wdata_a_i[3]), .A2(n7674), .B1(n4809), .B2(n8906), .ZN(
        n7672) );
  INV_X1 U6136 ( .A(n7673), .ZN(n8573) );
  AOI22_X1 U6137 ( .A1(wdata_a_i[2]), .A2(n7674), .B1(n4809), .B2(n8908), .ZN(
        n7673) );
  NOR2_X1 U6138 ( .A1(n1610), .A2(n4809), .ZN(n7674) );
  INV_X1 U6139 ( .A(n7675), .ZN(n8574) );
  AOI22_X1 U6140 ( .A1(wdata_a_i[1]), .A2(n7677), .B1(n4809), .B2(n8910), .ZN(
        n7675) );
  INV_X1 U6141 ( .A(n7676), .ZN(n8575) );
  AOI22_X1 U6142 ( .A1(wdata_a_i[0]), .A2(n7677), .B1(n4809), .B2(n4790), .ZN(
        n7676) );
  NOR2_X1 U6143 ( .A1(n1610), .A2(n4809), .ZN(n7677) );
  OR2_X1 U6144 ( .A1(n4809), .A2(n1611), .ZN(n8578) );
  NOR2_X1 U6145 ( .A1(n3849), .A2(n3851), .ZN(n7678) );
  INV_X1 U6146 ( .A(n7679), .ZN(n8581) );
  AOI22_X1 U6147 ( .A1(wdata_a_i[29]), .A2(n7681), .B1(n3851), .B2(n4796), 
        .ZN(n7679) );
  INV_X1 U6148 ( .A(n7680), .ZN(n8582) );
  AOI22_X1 U6149 ( .A1(n4618), .A2(n7681), .B1(n3851), .B2(wdata_b_i[28]), 
        .ZN(n7680) );
  NOR2_X1 U6150 ( .A1(n3849), .A2(n3851), .ZN(n7681) );
  INV_X1 U6151 ( .A(n7682), .ZN(n8583) );
  AOI22_X1 U6152 ( .A1(n4394), .A2(n7684), .B1(n3851), .B2(n9150), .ZN(n7682)
         );
  INV_X1 U6153 ( .A(n7683), .ZN(n8584) );
  AOI22_X1 U6154 ( .A1(n4459), .A2(n7684), .B1(n3851), .B2(n9063), .ZN(n7683)
         );
  NOR2_X1 U6155 ( .A1(n3849), .A2(n3851), .ZN(n7684) );
  INV_X1 U6156 ( .A(n7685), .ZN(n8585) );
  AOI22_X1 U6157 ( .A1(n4614), .A2(n7687), .B1(n3851), .B2(wdata_b_i[25]), 
        .ZN(n7685) );
  INV_X1 U6158 ( .A(n7686), .ZN(n8586) );
  AOI22_X1 U6159 ( .A1(wdata_a_i[24]), .A2(n7687), .B1(n3851), .B2(n8923), 
        .ZN(n7686) );
  NOR2_X1 U6160 ( .A1(n3849), .A2(n3851), .ZN(n7687) );
  NOR2_X1 U6161 ( .A1(n3849), .A2(n3851), .ZN(n7688) );
  NOR2_X1 U6162 ( .A1(n3849), .A2(n3851), .ZN(n7689) );
  NOR2_X1 U6163 ( .A1(n3849), .A2(n3851), .ZN(n7690) );
  INV_X1 U6164 ( .A(n7691), .ZN(n8594) );
  AOI22_X1 U6165 ( .A1(wdata_a_i[16]), .A2(n7692), .B1(n3851), .B2(n8883), 
        .ZN(n7691) );
  NOR2_X1 U6166 ( .A1(n3849), .A2(n3851), .ZN(n7692) );
  MUX2_X1 U6167 ( .A(wdata_a_i[15]), .B(n8885), .S(n3851), .Z(n8595) );
  INV_X1 U6168 ( .A(n7693), .ZN(n8596) );
  AOI22_X1 U6169 ( .A1(wdata_a_i[14]), .A2(n7695), .B1(n3851), .B2(n8887), 
        .ZN(n7693) );
  MUX2_X1 U6170 ( .A(wdata_a_i[13]), .B(wdata_b_i[13]), .S(n3851), .Z(n8597)
         );
  MUX2_X1 U6171 ( .A(wdata_a_i[12]), .B(n8890), .S(n3851), .Z(n8598) );
  MUX2_X1 U6172 ( .A(wdata_a_i[11]), .B(n4781), .S(n3851), .Z(n8599) );
  MUX2_X1 U6173 ( .A(wdata_a_i[10]), .B(n9089), .S(n3851), .Z(n8600) );
  MUX2_X1 U6174 ( .A(wdata_a_i[9]), .B(n4783), .S(n3851), .Z(n8601) );
  MUX2_X1 U6175 ( .A(wdata_a_i[8]), .B(wdata_b_i[8]), .S(n3851), .Z(n8602) );
  INV_X1 U6176 ( .A(n7694), .ZN(n8603) );
  AOI22_X1 U6177 ( .A1(n4486), .A2(n7695), .B1(n3851), .B2(n4780), .ZN(n7694)
         );
  NOR2_X1 U6178 ( .A1(n3849), .A2(n3851), .ZN(n7695) );
  MUX2_X1 U6179 ( .A(wdata_a_i[6]), .B(n4420), .S(n3851), .Z(n8604) );
  MUX2_X1 U6180 ( .A(wdata_a_i[5]), .B(n8902), .S(n3851), .Z(n8605) );
  INV_X1 U6181 ( .A(n7696), .ZN(n8606) );
  AOI22_X1 U6182 ( .A1(wdata_a_i[4]), .A2(n7698), .B1(n3851), .B2(n8904), .ZN(
        n7696) );
  INV_X1 U6183 ( .A(n7697), .ZN(n8607) );
  AOI22_X1 U6184 ( .A1(wdata_a_i[3]), .A2(n7698), .B1(n3851), .B2(n8906), .ZN(
        n7697) );
  NOR2_X1 U6185 ( .A1(n3849), .A2(n3851), .ZN(n7698) );
  MUX2_X1 U6186 ( .A(wdata_a_i[2]), .B(n8908), .S(n3851), .Z(n8608) );
  INV_X1 U6187 ( .A(n7699), .ZN(n8609) );
  AOI22_X1 U6188 ( .A1(wdata_a_i[1]), .A2(n7701), .B1(n3851), .B2(n8910), .ZN(
        n7699) );
  INV_X1 U6189 ( .A(n7700), .ZN(n8610) );
  AOI22_X1 U6190 ( .A1(wdata_a_i[0]), .A2(n7701), .B1(n3851), .B2(n9195), .ZN(
        n7700) );
  NOR2_X1 U6191 ( .A1(n3849), .A2(n3851), .ZN(n7701) );
  NAND2_X1 U6192 ( .A1(n3849), .A2(n4794), .ZN(n8613) );
  NOR2_X1 U6193 ( .A1(n1646), .A2(n1647), .ZN(n7702) );
  INV_X1 U6194 ( .A(n7703), .ZN(n8616) );
  AOI22_X1 U6195 ( .A1(wdata_a_i[29]), .A2(n7704), .B1(n1647), .B2(n4796), 
        .ZN(n7703) );
  NOR2_X1 U6196 ( .A1(n1646), .A2(n1647), .ZN(n7704) );
  INV_X1 U6197 ( .A(n7705), .ZN(n8617) );
  AOI22_X1 U6198 ( .A1(n4394), .A2(n7707), .B1(n1647), .B2(n9150), .ZN(n7705)
         );
  INV_X1 U6199 ( .A(n7706), .ZN(n8618) );
  AOI22_X1 U6200 ( .A1(n4459), .A2(n7707), .B1(n1647), .B2(n9063), .ZN(n7706)
         );
  NOR2_X1 U6201 ( .A1(n1646), .A2(n1647), .ZN(n7707) );
  INV_X1 U6202 ( .A(n7708), .ZN(n8619) );
  AOI22_X1 U6203 ( .A1(n4614), .A2(n7710), .B1(n1647), .B2(wdata_b_i[25]), 
        .ZN(n7708) );
  INV_X1 U6204 ( .A(n7709), .ZN(n8620) );
  AOI22_X1 U6205 ( .A1(wdata_a_i[24]), .A2(n7710), .B1(n1647), .B2(n8923), 
        .ZN(n7709) );
  NOR2_X1 U6206 ( .A1(n1646), .A2(n1647), .ZN(n7710) );
  NOR2_X1 U6207 ( .A1(n1646), .A2(n1647), .ZN(n7711) );
  NOR2_X1 U6208 ( .A1(n1646), .A2(n1647), .ZN(n7712) );
  NOR2_X1 U6209 ( .A1(n1646), .A2(n1647), .ZN(n7713) );
  INV_X1 U6210 ( .A(n7714), .ZN(n8628) );
  AOI22_X1 U6211 ( .A1(wdata_a_i[16]), .A2(n7715), .B1(n1647), .B2(n4734), 
        .ZN(n7714) );
  NOR2_X1 U6212 ( .A1(n1646), .A2(n1647), .ZN(n7715) );
  INV_X1 U6213 ( .A(n7716), .ZN(n8629) );
  AOI22_X1 U6214 ( .A1(wdata_a_i[15]), .A2(n7718), .B1(n1647), .B2(n8885), 
        .ZN(n7716) );
  INV_X1 U6215 ( .A(n7717), .ZN(n8630) );
  AOI22_X1 U6216 ( .A1(wdata_a_i[14]), .A2(n7718), .B1(n1647), .B2(n8887), 
        .ZN(n7717) );
  NOR2_X1 U6217 ( .A1(n1646), .A2(n1647), .ZN(n7718) );
  MUX2_X1 U6218 ( .A(wdata_a_i[13]), .B(wdata_b_i[13]), .S(n1647), .Z(n8631)
         );
  MUX2_X1 U6219 ( .A(wdata_a_i[12]), .B(n8890), .S(n1647), .Z(n8632) );
  MUX2_X1 U6220 ( .A(wdata_a_i[11]), .B(n4781), .S(n1647), .Z(n8633) );
  MUX2_X1 U6221 ( .A(wdata_a_i[10]), .B(n9089), .S(n1647), .Z(n8634) );
  MUX2_X1 U6222 ( .A(wdata_a_i[9]), .B(n4783), .S(n1647), .Z(n8635) );
  MUX2_X1 U6223 ( .A(wdata_a_i[8]), .B(wdata_b_i[8]), .S(n1647), .Z(n8636) );
  MUX2_X1 U6224 ( .A(n4486), .B(n4780), .S(n1647), .Z(n8637) );
  MUX2_X1 U6225 ( .A(wdata_a_i[6]), .B(n4420), .S(n1647), .Z(n8638) );
  MUX2_X1 U6226 ( .A(wdata_a_i[5]), .B(n8902), .S(n1647), .Z(n8639) );
  INV_X1 U6227 ( .A(n7719), .ZN(n8640) );
  AOI22_X1 U6228 ( .A1(wdata_a_i[4]), .A2(n7721), .B1(n1647), .B2(n4787), .ZN(
        n7719) );
  MUX2_X1 U6229 ( .A(wdata_a_i[3]), .B(n9100), .S(n1647), .Z(n8641) );
  INV_X1 U6230 ( .A(n7720), .ZN(n8642) );
  AOI22_X1 U6231 ( .A1(wdata_a_i[2]), .A2(n7721), .B1(n1647), .B2(n8908), .ZN(
        n7720) );
  NOR2_X1 U6232 ( .A1(n1646), .A2(n1647), .ZN(n7721) );
  INV_X1 U6233 ( .A(n7722), .ZN(n8643) );
  AOI22_X1 U6234 ( .A1(wdata_a_i[1]), .A2(n7724), .B1(n1647), .B2(n8910), .ZN(
        n7722) );
  INV_X1 U6235 ( .A(n7723), .ZN(n8644) );
  AOI22_X1 U6236 ( .A1(wdata_a_i[0]), .A2(n7724), .B1(n1647), .B2(n4791), .ZN(
        n7723) );
  NOR2_X1 U6237 ( .A1(n1646), .A2(n1647), .ZN(n7724) );
  OR2_X1 U6238 ( .A1(n1648), .A2(n1647), .ZN(n8647) );
  NOR2_X1 U6239 ( .A1(n3772), .A2(n3774), .ZN(n7725) );
  INV_X1 U6240 ( .A(n7726), .ZN(n8650) );
  AOI22_X1 U6241 ( .A1(n4468), .A2(n7728), .B1(n3774), .B2(n4796), .ZN(n7726)
         );
  INV_X1 U6242 ( .A(n7727), .ZN(n8651) );
  AOI22_X1 U6243 ( .A1(n4618), .A2(n7728), .B1(n3774), .B2(wdata_b_i[28]), 
        .ZN(n7727) );
  NOR2_X1 U6244 ( .A1(n3772), .A2(n3774), .ZN(n7728) );
  INV_X1 U6245 ( .A(n7729), .ZN(n8652) );
  AOI22_X1 U6246 ( .A1(n4394), .A2(n7731), .B1(n3774), .B2(n9150), .ZN(n7729)
         );
  INV_X1 U6247 ( .A(n7730), .ZN(n8653) );
  AOI22_X1 U6248 ( .A1(n4459), .A2(n7731), .B1(n3774), .B2(n9063), .ZN(n7730)
         );
  NOR2_X1 U6249 ( .A1(n3772), .A2(n3774), .ZN(n7731) );
  INV_X1 U6250 ( .A(n7732), .ZN(n8654) );
  AOI22_X1 U6251 ( .A1(n4614), .A2(n7734), .B1(n3774), .B2(wdata_b_i[25]), 
        .ZN(n7732) );
  INV_X1 U6252 ( .A(n7733), .ZN(n8655) );
  AOI22_X1 U6253 ( .A1(wdata_a_i[24]), .A2(n7734), .B1(n3774), .B2(n8923), 
        .ZN(n7733) );
  NOR2_X1 U6254 ( .A1(n3772), .A2(n3774), .ZN(n7734) );
  NOR2_X1 U6255 ( .A1(n3772), .A2(n3774), .ZN(n7735) );
  NOR2_X1 U6256 ( .A1(n3772), .A2(n3774), .ZN(n7736) );
  NOR2_X1 U6257 ( .A1(n3772), .A2(n3774), .ZN(n7737) );
  INV_X1 U6258 ( .A(n7738), .ZN(n8663) );
  AOI22_X1 U6259 ( .A1(wdata_a_i[16]), .A2(n7739), .B1(n3774), .B2(n4734), 
        .ZN(n7738) );
  NOR2_X1 U6260 ( .A1(n3772), .A2(n3774), .ZN(n7739) );
  MUX2_X1 U6261 ( .A(wdata_a_i[15]), .B(n9081), .S(n3774), .Z(n8664) );
  INV_X1 U6262 ( .A(n7740), .ZN(n8665) );
  AOI22_X1 U6263 ( .A1(wdata_a_i[14]), .A2(n7742), .B1(n3774), .B2(n8887), 
        .ZN(n7740) );
  MUX2_X1 U6264 ( .A(wdata_a_i[13]), .B(wdata_b_i[13]), .S(n3774), .Z(n8666)
         );
  MUX2_X1 U6265 ( .A(wdata_a_i[12]), .B(n8890), .S(n3774), .Z(n8667) );
  MUX2_X1 U6266 ( .A(wdata_a_i[11]), .B(n4781), .S(n3774), .Z(n8668) );
  MUX2_X1 U6267 ( .A(wdata_a_i[10]), .B(n9089), .S(n3774), .Z(n8669) );
  MUX2_X1 U6268 ( .A(wdata_a_i[9]), .B(n4783), .S(n3774), .Z(n8670) );
  MUX2_X1 U6269 ( .A(wdata_a_i[8]), .B(n8898), .S(n3774), .Z(n8671) );
  INV_X1 U6270 ( .A(n7741), .ZN(n8672) );
  AOI22_X1 U6271 ( .A1(n4486), .A2(n7742), .B1(n3774), .B2(n4779), .ZN(n7741)
         );
  NOR2_X1 U6272 ( .A1(n3772), .A2(n3774), .ZN(n7742) );
  MUX2_X1 U6273 ( .A(wdata_a_i[6]), .B(n4420), .S(n3774), .Z(n8673) );
  MUX2_X1 U6274 ( .A(wdata_a_i[5]), .B(n9096), .S(n3774), .Z(n8674) );
  INV_X1 U6275 ( .A(n7743), .ZN(n8675) );
  AOI22_X1 U6276 ( .A1(wdata_a_i[4]), .A2(n7745), .B1(n3774), .B2(n4787), .ZN(
        n7743) );
  INV_X1 U6277 ( .A(n7744), .ZN(n8676) );
  AOI22_X1 U6278 ( .A1(wdata_a_i[3]), .A2(n7745), .B1(n3774), .B2(n9100), .ZN(
        n7744) );
  NOR2_X1 U6279 ( .A1(n3772), .A2(n3774), .ZN(n7745) );
  MUX2_X1 U6280 ( .A(wdata_a_i[2]), .B(n8908), .S(n3774), .Z(n8677) );
  INV_X1 U6281 ( .A(n7746), .ZN(n8678) );
  AOI22_X1 U6282 ( .A1(wdata_a_i[1]), .A2(n7748), .B1(n3774), .B2(n8910), .ZN(
        n7746) );
  INV_X1 U6283 ( .A(n7747), .ZN(n8679) );
  AOI22_X1 U6284 ( .A1(wdata_a_i[0]), .A2(n7748), .B1(n3774), .B2(n4790), .ZN(
        n7747) );
  NOR2_X1 U6285 ( .A1(n3772), .A2(n3774), .ZN(n7748) );
  NAND2_X1 U6286 ( .A1(n3772), .A2(n4827), .ZN(n8682) );
  NOR2_X1 U6287 ( .A1(n1616), .A2(n1617), .ZN(n7749) );
  MUX2_X1 U6288 ( .A(n4468), .B(n4796), .S(n1617), .Z(n8685) );
  MUX2_X1 U6289 ( .A(n4618), .B(wdata_b_i[28]), .S(n1617), .Z(n8686) );
  MUX2_X1 U6290 ( .A(n4394), .B(n4732), .S(n1617), .Z(n8687) );
  MUX2_X1 U6291 ( .A(n4459), .B(n8867), .S(n1617), .Z(n8688) );
  MUX2_X1 U6292 ( .A(n4614), .B(wdata_b_i[25]), .S(n1617), .Z(n8689) );
  MUX2_X1 U6293 ( .A(n4386), .B(n8923), .S(n1617), .Z(n8690) );
  NOR2_X1 U6294 ( .A1(n1616), .A2(n1617), .ZN(n7750) );
  MUX2_X1 U6295 ( .A(wdata_a_i[21]), .B(n9032), .S(n1617), .Z(n8693) );
  NOR2_X1 U6296 ( .A1(n1616), .A2(n1617), .ZN(n7751) );
  NOR2_X1 U6297 ( .A1(n1616), .A2(n1617), .ZN(n7752) );
  INV_X1 U6298 ( .A(n7753), .ZN(n8698) );
  AOI22_X1 U6299 ( .A1(wdata_a_i[16]), .A2(n7755), .B1(n1617), .B2(n4734), 
        .ZN(n7753) );
  INV_X1 U6300 ( .A(n7754), .ZN(n8699) );
  AOI22_X1 U6301 ( .A1(wdata_a_i[15]), .A2(n7755), .B1(n1617), .B2(n9081), 
        .ZN(n7754) );
  NOR2_X1 U6302 ( .A1(n1616), .A2(n1617), .ZN(n7755) );
  MUX2_X1 U6303 ( .A(wdata_a_i[14]), .B(n8887), .S(n1617), .Z(n8700) );
  MUX2_X1 U6304 ( .A(wdata_a_i[13]), .B(wdata_b_i[13]), .S(n1617), .Z(n8701)
         );
  MUX2_X1 U6305 ( .A(wdata_a_i[12]), .B(n8890), .S(n1617), .Z(n8702) );
  INV_X1 U6306 ( .A(n7756), .ZN(n8703) );
  AOI22_X1 U6307 ( .A1(wdata_a_i[11]), .A2(n7757), .B1(n1617), .B2(n4781), 
        .ZN(n7756) );
  NOR2_X1 U6308 ( .A1(n1616), .A2(n1617), .ZN(n7757) );
  INV_X1 U6309 ( .A(n7758), .ZN(n8705) );
  AOI22_X1 U6310 ( .A1(wdata_a_i[9]), .A2(n7760), .B1(n1617), .B2(n9091), .ZN(
        n7758) );
  INV_X1 U6311 ( .A(n7759), .ZN(n8706) );
  AOI22_X1 U6312 ( .A1(wdata_a_i[8]), .A2(n7760), .B1(n1617), .B2(n4774), .ZN(
        n7759) );
  NOR2_X1 U6313 ( .A1(n1616), .A2(n1617), .ZN(n7760) );
  INV_X1 U6314 ( .A(n7761), .ZN(n8707) );
  AOI22_X1 U6315 ( .A1(n4486), .A2(n7763), .B1(n1617), .B2(n9182), .ZN(n7761)
         );
  INV_X1 U6316 ( .A(n7762), .ZN(n8708) );
  AOI22_X1 U6317 ( .A1(wdata_a_i[6]), .A2(n7763), .B1(n1617), .B2(n4420), .ZN(
        n7762) );
  NOR2_X1 U6318 ( .A1(n1616), .A2(n1617), .ZN(n7763) );
  INV_X1 U6319 ( .A(n7764), .ZN(n8709) );
  AOI22_X1 U6320 ( .A1(wdata_a_i[5]), .A2(n7766), .B1(n1617), .B2(n9186), .ZN(
        n7764) );
  INV_X1 U6321 ( .A(n7765), .ZN(n8710) );
  AOI22_X1 U6322 ( .A1(wdata_a_i[4]), .A2(n7766), .B1(n1617), .B2(n4787), .ZN(
        n7765) );
  NOR2_X1 U6323 ( .A1(n1616), .A2(n1617), .ZN(n7766) );
  INV_X1 U6324 ( .A(n7767), .ZN(n8711) );
  AOI22_X1 U6325 ( .A1(wdata_a_i[3]), .A2(n7769), .B1(n1617), .B2(n8906), .ZN(
        n7767) );
  INV_X1 U6326 ( .A(n7768), .ZN(n8712) );
  AOI22_X1 U6327 ( .A1(wdata_a_i[2]), .A2(n7769), .B1(n1617), .B2(n8908), .ZN(
        n7768) );
  NOR2_X1 U6328 ( .A1(n1616), .A2(n1617), .ZN(n7769) );
  INV_X1 U6329 ( .A(n7770), .ZN(n8713) );
  AOI22_X1 U6330 ( .A1(wdata_a_i[1]), .A2(n7772), .B1(n1617), .B2(n8910), .ZN(
        n7770) );
  INV_X1 U6331 ( .A(n7771), .ZN(n8714) );
  AOI22_X1 U6332 ( .A1(wdata_a_i[0]), .A2(n7772), .B1(n1617), .B2(n4791), .ZN(
        n7771) );
  NOR2_X1 U6333 ( .A1(n1616), .A2(n1617), .ZN(n7772) );
  OR2_X1 U6334 ( .A1(n1618), .A2(n1617), .ZN(n8717) );
  NOR2_X1 U6335 ( .A1(n1632), .A2(n1634), .ZN(n7773) );
  INV_X1 U6336 ( .A(n7774), .ZN(n8720) );
  AOI22_X1 U6337 ( .A1(n4468), .A2(n7776), .B1(n1634), .B2(n4796), .ZN(n7774)
         );
  INV_X1 U6338 ( .A(n7775), .ZN(n8721) );
  AOI22_X1 U6339 ( .A1(n4618), .A2(n7776), .B1(n1634), .B2(wdata_b_i[28]), 
        .ZN(n7775) );
  NOR2_X1 U6340 ( .A1(n1632), .A2(n1634), .ZN(n7776) );
  INV_X1 U6341 ( .A(n7777), .ZN(n8722) );
  AOI22_X1 U6342 ( .A1(n4394), .A2(n7779), .B1(n1634), .B2(n9150), .ZN(n7777)
         );
  INV_X1 U6343 ( .A(n7778), .ZN(n8723) );
  AOI22_X1 U6344 ( .A1(n4459), .A2(n7779), .B1(n1634), .B2(n9063), .ZN(n7778)
         );
  NOR2_X1 U6345 ( .A1(n1632), .A2(n1634), .ZN(n7779) );
  INV_X1 U6346 ( .A(n7780), .ZN(n8724) );
  AOI22_X1 U6347 ( .A1(n4614), .A2(n7782), .B1(n1634), .B2(wdata_b_i[25]), 
        .ZN(n7780) );
  INV_X1 U6348 ( .A(n7781), .ZN(n8725) );
  AOI22_X1 U6349 ( .A1(wdata_a_i[24]), .A2(n7782), .B1(n1634), .B2(n8923), 
        .ZN(n7781) );
  NOR2_X1 U6350 ( .A1(n1632), .A2(n1634), .ZN(n7782) );
  NOR2_X1 U6351 ( .A1(n1632), .A2(n1634), .ZN(n7783) );
  NOR2_X1 U6352 ( .A1(n1632), .A2(n1634), .ZN(n7784) );
  NOR2_X1 U6353 ( .A1(n1632), .A2(n1634), .ZN(n7785) );
  INV_X1 U6354 ( .A(n7786), .ZN(n8733) );
  AOI22_X1 U6355 ( .A1(wdata_a_i[16]), .A2(n7787), .B1(n1634), .B2(n4734), 
        .ZN(n7786) );
  NOR2_X1 U6356 ( .A1(n1632), .A2(n1634), .ZN(n7787) );
  INV_X1 U6357 ( .A(n7788), .ZN(n8734) );
  AOI22_X1 U6358 ( .A1(wdata_a_i[15]), .A2(n7790), .B1(n1634), .B2(n8885), 
        .ZN(n7788) );
  INV_X1 U6359 ( .A(n7789), .ZN(n8735) );
  AOI22_X1 U6360 ( .A1(wdata_a_i[14]), .A2(n7790), .B1(n1634), .B2(n8887), 
        .ZN(n7789) );
  NOR2_X1 U6361 ( .A1(n1632), .A2(n1634), .ZN(n7790) );
  MUX2_X1 U6362 ( .A(wdata_a_i[13]), .B(wdata_b_i[13]), .S(n1634), .Z(n8736)
         );
  MUX2_X1 U6363 ( .A(wdata_a_i[12]), .B(n8890), .S(n1634), .Z(n8737) );
  MUX2_X1 U6364 ( .A(wdata_a_i[11]), .B(n4781), .S(n1634), .Z(n8738) );
  MUX2_X1 U6365 ( .A(wdata_a_i[10]), .B(n9089), .S(n1634), .Z(n8739) );
  MUX2_X1 U6366 ( .A(wdata_a_i[9]), .B(n4783), .S(n1634), .Z(n8740) );
  MUX2_X1 U6367 ( .A(wdata_a_i[8]), .B(n8898), .S(n1634), .Z(n8741) );
  MUX2_X1 U6368 ( .A(n4486), .B(n4779), .S(n1634), .Z(n8742) );
  MUX2_X1 U6369 ( .A(wdata_a_i[6]), .B(n4420), .S(n1634), .Z(n8743) );
  MUX2_X1 U6370 ( .A(wdata_a_i[5]), .B(n9096), .S(n1634), .Z(n8744) );
  INV_X1 U6371 ( .A(n7791), .ZN(n8745) );
  AOI22_X1 U6372 ( .A1(wdata_a_i[4]), .A2(n7793), .B1(n1634), .B2(n4787), .ZN(
        n7791) );
  MUX2_X1 U6373 ( .A(wdata_a_i[3]), .B(n8906), .S(n1634), .Z(n8746) );
  INV_X1 U6374 ( .A(n7792), .ZN(n8747) );
  AOI22_X1 U6375 ( .A1(wdata_a_i[2]), .A2(n7793), .B1(n1634), .B2(n8908), .ZN(
        n7792) );
  NOR2_X1 U6376 ( .A1(n1632), .A2(n1634), .ZN(n7793) );
  INV_X1 U6377 ( .A(n7794), .ZN(n8748) );
  AOI22_X1 U6378 ( .A1(wdata_a_i[1]), .A2(n7796), .B1(n1634), .B2(n8910), .ZN(
        n7794) );
  INV_X1 U6379 ( .A(n7795), .ZN(n8749) );
  AOI22_X1 U6380 ( .A1(wdata_a_i[0]), .A2(n7796), .B1(n1634), .B2(n4790), .ZN(
        n7795) );
  NOR2_X1 U6381 ( .A1(n1632), .A2(n1634), .ZN(n7796) );
  NAND2_X1 U6382 ( .A1(n1632), .A2(n7797), .ZN(n8752) );
  INV_X1 U6383 ( .A(n1634), .ZN(n7797) );
  NOR2_X1 U6384 ( .A1(n1639), .A2(n1640), .ZN(n7798) );
  MUX2_X1 U6385 ( .A(n4468), .B(n4796), .S(n1640), .Z(n8755) );
  MUX2_X1 U6386 ( .A(n4618), .B(wdata_b_i[28]), .S(n1640), .Z(n8756) );
  MUX2_X1 U6387 ( .A(n4394), .B(n8865), .S(n1640), .Z(n8757) );
  MUX2_X1 U6388 ( .A(n4459), .B(n9152), .S(n1640), .Z(n8758) );
  MUX2_X1 U6389 ( .A(n4614), .B(wdata_b_i[25]), .S(n1640), .Z(n8759) );
  MUX2_X1 U6390 ( .A(wdata_a_i[24]), .B(n8923), .S(n1640), .Z(n8760) );
  NOR2_X1 U6391 ( .A1(n1639), .A2(n1640), .ZN(n7799) );
  MUX2_X1 U6392 ( .A(wdata_a_i[21]), .B(n9032), .S(n1640), .Z(n8763) );
  NOR2_X1 U6393 ( .A1(n1639), .A2(n1640), .ZN(n7800) );
  NOR2_X1 U6394 ( .A1(n1639), .A2(n1640), .ZN(n7801) );
  INV_X1 U6395 ( .A(n7802), .ZN(n8768) );
  AOI22_X1 U6396 ( .A1(wdata_a_i[16]), .A2(n7804), .B1(n1640), .B2(n4734), 
        .ZN(n7802) );
  INV_X1 U6397 ( .A(n7803), .ZN(n8769) );
  AOI22_X1 U6398 ( .A1(wdata_a_i[15]), .A2(n7804), .B1(n1640), .B2(n9081), 
        .ZN(n7803) );
  NOR2_X1 U6399 ( .A1(n1639), .A2(n1640), .ZN(n7804) );
  MUX2_X1 U6400 ( .A(wdata_a_i[14]), .B(n8887), .S(n1640), .Z(n8770) );
  MUX2_X1 U6401 ( .A(wdata_a_i[13]), .B(wdata_b_i[13]), .S(n1640), .Z(n8771)
         );
  MUX2_X1 U6402 ( .A(wdata_a_i[12]), .B(n8890), .S(n1640), .Z(n8772) );
  INV_X1 U6403 ( .A(n7805), .ZN(n8773) );
  AOI22_X1 U6404 ( .A1(wdata_a_i[11]), .A2(n7806), .B1(n1640), .B2(n4781), 
        .ZN(n7805) );
  NOR2_X1 U6405 ( .A1(n1639), .A2(n1640), .ZN(n7806) );
  INV_X1 U6406 ( .A(n7807), .ZN(n8775) );
  AOI22_X1 U6407 ( .A1(wdata_a_i[9]), .A2(n7809), .B1(n1640), .B2(n8896), .ZN(
        n7807) );
  INV_X1 U6408 ( .A(n7808), .ZN(n8776) );
  AOI22_X1 U6409 ( .A1(wdata_a_i[8]), .A2(n7809), .B1(n1640), .B2(n4774), .ZN(
        n7808) );
  NOR2_X1 U6410 ( .A1(n1639), .A2(n1640), .ZN(n7809) );
  INV_X1 U6411 ( .A(n7810), .ZN(n8777) );
  AOI22_X1 U6412 ( .A1(n4486), .A2(n7812), .B1(n1640), .B2(n9182), .ZN(n7810)
         );
  INV_X1 U6413 ( .A(n7811), .ZN(n8778) );
  AOI22_X1 U6414 ( .A1(wdata_a_i[6]), .A2(n7812), .B1(n1640), .B2(n4420), .ZN(
        n7811) );
  NOR2_X1 U6415 ( .A1(n1639), .A2(n1640), .ZN(n7812) );
  INV_X1 U6416 ( .A(n7813), .ZN(n8779) );
  AOI22_X1 U6417 ( .A1(wdata_a_i[5]), .A2(n7815), .B1(n1640), .B2(n9186), .ZN(
        n7813) );
  INV_X1 U6418 ( .A(n7814), .ZN(n8780) );
  AOI22_X1 U6419 ( .A1(wdata_a_i[4]), .A2(n7815), .B1(n1640), .B2(n4787), .ZN(
        n7814) );
  NOR2_X1 U6420 ( .A1(n1639), .A2(n1640), .ZN(n7815) );
  INV_X1 U6421 ( .A(n7816), .ZN(n8781) );
  AOI22_X1 U6422 ( .A1(wdata_a_i[3]), .A2(n7818), .B1(n1640), .B2(n8906), .ZN(
        n7816) );
  INV_X1 U6423 ( .A(n7817), .ZN(n8782) );
  AOI22_X1 U6424 ( .A1(wdata_a_i[2]), .A2(n7818), .B1(n1640), .B2(n8908), .ZN(
        n7817) );
  NOR2_X1 U6425 ( .A1(n1639), .A2(n1640), .ZN(n7818) );
  INV_X1 U6426 ( .A(n7819), .ZN(n8783) );
  AOI22_X1 U6427 ( .A1(wdata_a_i[1]), .A2(n7821), .B1(n1640), .B2(n8910), .ZN(
        n7819) );
  INV_X1 U6428 ( .A(n7820), .ZN(n8784) );
  AOI22_X1 U6429 ( .A1(wdata_a_i[0]), .A2(n7821), .B1(n1640), .B2(n4791), .ZN(
        n7820) );
  NOR2_X1 U6430 ( .A1(n1639), .A2(n1640), .ZN(n7821) );
  OR2_X1 U6431 ( .A1(n1641), .A2(n1640), .ZN(n8787) );
  NOR2_X1 U6432 ( .A1(n2535), .A2(n4821), .ZN(n7822) );
  INV_X1 U6433 ( .A(n7823), .ZN(n8791) );
  AOI22_X1 U6434 ( .A1(wdata_a_i[28]), .A2(n7824), .B1(n4821), .B2(
        wdata_b_i[28]), .ZN(n7823) );
  NOR2_X1 U6435 ( .A1(n2535), .A2(n4821), .ZN(n7824) );
  INV_X1 U6436 ( .A(n7825), .ZN(n8792) );
  AOI22_X1 U6437 ( .A1(wdata_a_i[27]), .A2(n7827), .B1(n4821), .B2(n4732), 
        .ZN(n7825) );
  INV_X1 U6438 ( .A(n7826), .ZN(n8793) );
  AOI22_X1 U6439 ( .A1(wdata_a_i[26]), .A2(n7827), .B1(n4821), .B2(n9063), 
        .ZN(n7826) );
  NOR2_X1 U6440 ( .A1(n2535), .A2(n4821), .ZN(n7827) );
  INV_X1 U6441 ( .A(n7828), .ZN(n8794) );
  AOI22_X1 U6442 ( .A1(wdata_a_i[25]), .A2(n7830), .B1(n4821), .B2(
        wdata_b_i[25]), .ZN(n7828) );
  INV_X1 U6443 ( .A(n7829), .ZN(n8795) );
  AOI22_X1 U6444 ( .A1(wdata_a_i[24]), .A2(n7830), .B1(n4821), .B2(n9155), 
        .ZN(n7829) );
  NOR2_X1 U6445 ( .A1(n2535), .A2(n4821), .ZN(n7830) );
  NOR2_X1 U6446 ( .A1(n2535), .A2(n4821), .ZN(n7831) );
  NOR2_X1 U6447 ( .A1(n2535), .A2(n4821), .ZN(n7832) );
  NOR2_X1 U6448 ( .A1(n2535), .A2(n4821), .ZN(n7833) );
  INV_X1 U6449 ( .A(n7834), .ZN(n8803) );
  AOI22_X1 U6450 ( .A1(wdata_a_i[16]), .A2(n7835), .B1(n4821), .B2(n8349), 
        .ZN(n7834) );
  NOR2_X1 U6451 ( .A1(n2535), .A2(n4821), .ZN(n7835) );
  MUX2_X1 U6452 ( .A(wdata_a_i[14]), .B(n9172), .S(n4821), .Z(n8805) );
  MUX2_X1 U6453 ( .A(wdata_a_i[13]), .B(n9174), .S(n4821), .Z(n8806) );
  MUX2_X1 U6454 ( .A(wdata_a_i[12]), .B(n9085), .S(n4821), .Z(n8807) );
  MUX2_X1 U6455 ( .A(wdata_a_i[11]), .B(n9087), .S(n4821), .Z(n8808) );
  MUX2_X1 U6456 ( .A(wdata_a_i[10]), .B(n9089), .S(n4821), .Z(n8809) );
  MUX2_X1 U6457 ( .A(wdata_a_i[9]), .B(n4783), .S(n4821), .Z(n8810) );
  MUX2_X1 U6458 ( .A(wdata_a_i[8]), .B(n4774), .S(n4821), .Z(n8811) );
  MUX2_X1 U6459 ( .A(wdata_a_i[7]), .B(wdata_b_i[7]), .S(n4821), .Z(n8812) );
  MUX2_X1 U6460 ( .A(wdata_a_i[6]), .B(n4420), .S(n4821), .Z(n8813) );
  INV_X1 U6461 ( .A(n7836), .ZN(n8814) );
  AOI22_X1 U6462 ( .A1(wdata_a_i[5]), .A2(n7837), .B1(n4821), .B2(n9096), .ZN(
        n7836) );
  NOR2_X1 U6463 ( .A1(n2535), .A2(n4821), .ZN(n7837) );
  INV_X1 U6464 ( .A(n7838), .ZN(n8815) );
  AOI22_X1 U6465 ( .A1(wdata_a_i[4]), .A2(n7840), .B1(n4821), .B2(n9098), .ZN(
        n7838) );
  MUX2_X1 U6466 ( .A(wdata_a_i[3]), .B(n9100), .S(n4821), .Z(n8816) );
  INV_X1 U6467 ( .A(n7839), .ZN(n8817) );
  AOI22_X1 U6468 ( .A1(wdata_a_i[2]), .A2(n7840), .B1(n4821), .B2(n9102), .ZN(
        n7839) );
  NOR2_X1 U6469 ( .A1(n2535), .A2(n4821), .ZN(n7840) );
  INV_X1 U6470 ( .A(n7841), .ZN(n8818) );
  AOI22_X1 U6471 ( .A1(wdata_a_i[1]), .A2(n7843), .B1(n4821), .B2(n9104), .ZN(
        n7841) );
  INV_X1 U6472 ( .A(n7842), .ZN(n8819) );
  AOI22_X1 U6473 ( .A1(wdata_a_i[0]), .A2(n7843), .B1(n4821), .B2(n4790), .ZN(
        n7842) );
  NOR2_X1 U6474 ( .A1(n2535), .A2(n4821), .ZN(n7843) );
  NAND2_X1 U6475 ( .A1(n2535), .A2(n4764), .ZN(n8822) );
  NOR2_X1 U6476 ( .A1(n1627), .A2(n1629), .ZN(n7844) );
  INV_X1 U6477 ( .A(n7845), .ZN(n8825) );
  AOI22_X1 U6478 ( .A1(n4468), .A2(n7847), .B1(n1629), .B2(n4796), .ZN(n7845)
         );
  INV_X1 U6479 ( .A(n7846), .ZN(n8826) );
  AOI22_X1 U6480 ( .A1(n4618), .A2(n7847), .B1(n1629), .B2(wdata_b_i[28]), 
        .ZN(n7846) );
  NOR2_X1 U6481 ( .A1(n1627), .A2(n1629), .ZN(n7847) );
  INV_X1 U6482 ( .A(n7848), .ZN(n8827) );
  AOI22_X1 U6483 ( .A1(n4394), .A2(n7850), .B1(n1629), .B2(n9150), .ZN(n7848)
         );
  INV_X1 U6484 ( .A(n7849), .ZN(n8828) );
  AOI22_X1 U6485 ( .A1(n4459), .A2(n7850), .B1(n1629), .B2(n9063), .ZN(n7849)
         );
  NOR2_X1 U6486 ( .A1(n1627), .A2(n1629), .ZN(n7850) );
  INV_X1 U6487 ( .A(n7851), .ZN(n8829) );
  AOI22_X1 U6488 ( .A1(n4614), .A2(n7853), .B1(n1629), .B2(wdata_b_i[25]), 
        .ZN(n7851) );
  INV_X1 U6489 ( .A(n7852), .ZN(n8830) );
  AOI22_X1 U6490 ( .A1(n4386), .A2(n7853), .B1(n1629), .B2(n8923), .ZN(n7852)
         );
  NOR2_X1 U6491 ( .A1(n1627), .A2(n1629), .ZN(n7853) );
  NOR2_X1 U6492 ( .A1(n1627), .A2(n1629), .ZN(n7854) );
  NOR2_X1 U6493 ( .A1(n1627), .A2(n1629), .ZN(n7855) );
  NOR2_X1 U6494 ( .A1(n1627), .A2(n1629), .ZN(n7856) );
  INV_X1 U6495 ( .A(n7857), .ZN(n8838) );
  AOI22_X1 U6496 ( .A1(wdata_a_i[16]), .A2(n7858), .B1(n1629), .B2(n8883), 
        .ZN(n7857) );
  NOR2_X1 U6497 ( .A1(n1627), .A2(n1629), .ZN(n7858) );
  INV_X1 U6498 ( .A(n7859), .ZN(n8839) );
  AOI22_X1 U6499 ( .A1(wdata_a_i[15]), .A2(n7861), .B1(n1629), .B2(n8885), 
        .ZN(n7859) );
  INV_X1 U6500 ( .A(n7860), .ZN(n8840) );
  AOI22_X1 U6501 ( .A1(wdata_a_i[14]), .A2(n7861), .B1(n1629), .B2(n8887), 
        .ZN(n7860) );
  NOR2_X1 U6502 ( .A1(n1627), .A2(n1629), .ZN(n7861) );
  MUX2_X1 U6503 ( .A(wdata_a_i[13]), .B(wdata_b_i[13]), .S(n1629), .Z(n8841)
         );
  MUX2_X1 U6504 ( .A(wdata_a_i[12]), .B(n8890), .S(n1629), .Z(n8842) );
  MUX2_X1 U6505 ( .A(wdata_a_i[11]), .B(n4781), .S(n1629), .Z(n8843) );
  MUX2_X1 U6506 ( .A(wdata_a_i[10]), .B(n9089), .S(n1629), .Z(n8844) );
  MUX2_X1 U6507 ( .A(wdata_a_i[9]), .B(n4783), .S(n1629), .Z(n8845) );
  MUX2_X1 U6508 ( .A(wdata_a_i[8]), .B(n8898), .S(n1629), .Z(n8846) );
  MUX2_X1 U6509 ( .A(n4486), .B(n8848), .S(n1629), .Z(n8847) );
  MUX2_X1 U6510 ( .A(wdata_a_i[6]), .B(n4420), .S(n1629), .Z(n8849) );
  MUX2_X1 U6511 ( .A(wdata_a_i[5]), .B(n8902), .S(n1629), .Z(n8850) );
  INV_X1 U6512 ( .A(n7862), .ZN(n8851) );
  AOI22_X1 U6513 ( .A1(wdata_a_i[4]), .A2(n7864), .B1(n1629), .B2(n4787), .ZN(
        n7862) );
  MUX2_X1 U6514 ( .A(wdata_a_i[3]), .B(n9100), .S(n1629), .Z(n8852) );
  INV_X1 U6515 ( .A(n7863), .ZN(n8853) );
  AOI22_X1 U6516 ( .A1(wdata_a_i[2]), .A2(n7864), .B1(n1629), .B2(n8908), .ZN(
        n7863) );
  NOR2_X1 U6517 ( .A1(n1627), .A2(n1629), .ZN(n7864) );
  INV_X1 U6518 ( .A(n7865), .ZN(n8854) );
  AOI22_X1 U6519 ( .A1(wdata_a_i[1]), .A2(n7867), .B1(n1629), .B2(n8910), .ZN(
        n7865) );
  INV_X1 U6520 ( .A(n7866), .ZN(n8855) );
  AOI22_X1 U6521 ( .A1(wdata_a_i[0]), .A2(n7867), .B1(n1629), .B2(n4790), .ZN(
        n7866) );
  NOR2_X1 U6522 ( .A1(n1627), .A2(n1629), .ZN(n7867) );
  NAND2_X1 U6523 ( .A1(n1627), .A2(n7868), .ZN(n8858) );
  INV_X1 U6524 ( .A(n1629), .ZN(n7868) );
  OAI22_X1 U6525 ( .A1(n1623), .A2(n7869), .B1(n4474), .B2(n4744), .ZN(n8859)
         );
  NAND2_X1 U6526 ( .A1(n4477), .A2(n4744), .ZN(n7869) );
  OAI22_X1 U6527 ( .A1(n1623), .A2(n7870), .B1(n4470), .B2(n4744), .ZN(n8860)
         );
  NAND2_X1 U6528 ( .A1(n4623), .A2(n4744), .ZN(n7870) );
  OAI22_X1 U6529 ( .A1(n1623), .A2(n7871), .B1(n4467), .B2(n4744), .ZN(n8862)
         );
  NAND2_X1 U6530 ( .A1(n4468), .A2(n4744), .ZN(n7871) );
  OAI22_X1 U6531 ( .A1(n1623), .A2(n7872), .B1(n4017), .B2(n4744), .ZN(n8863)
         );
  NAND2_X1 U6532 ( .A1(n4618), .A2(n4744), .ZN(n7872) );
  OAI22_X1 U6533 ( .A1(n1623), .A2(n7873), .B1(n4795), .B2(n4744), .ZN(n8864)
         );
  NAND2_X1 U6534 ( .A1(n4394), .A2(n4744), .ZN(n7873) );
  INV_X1 U6535 ( .A(n4461), .ZN(n8865) );
  OAI22_X1 U6536 ( .A1(n1623), .A2(n7874), .B1(n4458), .B2(n4744), .ZN(n8866)
         );
  NAND2_X1 U6537 ( .A1(n4459), .A2(n4744), .ZN(n7874) );
  INV_X1 U6538 ( .A(n4458), .ZN(n8867) );
  OAI22_X1 U6539 ( .A1(n1623), .A2(n7875), .B1(n4011), .B2(n4744), .ZN(n8868)
         );
  NAND2_X1 U6540 ( .A1(n4614), .A2(n4744), .ZN(n7875) );
  INV_X1 U6541 ( .A(n7876), .ZN(n8869) );
  AOI22_X1 U6542 ( .A1(wdata_a_i[24]), .A2(n7877), .B1(n1624), .B2(n8923), 
        .ZN(n7876) );
  NOR2_X1 U6543 ( .A1(n1623), .A2(n1624), .ZN(n7877) );
  OAI22_X1 U6544 ( .A1(n1623), .A2(n7878), .B1(n4385), .B2(n4744), .ZN(n8870)
         );
  NAND2_X1 U6545 ( .A1(wdata_a_i[23]), .A2(n4744), .ZN(n7878) );
  OAI22_X1 U6546 ( .A1(n1623), .A2(n7879), .B1(n4004), .B2(n4744), .ZN(n8872)
         );
  NAND2_X1 U6547 ( .A1(wdata_a_i[22]), .A2(n4744), .ZN(n7879) );
  OAI22_X1 U6548 ( .A1(n1623), .A2(n7880), .B1(n4002), .B2(n4744), .ZN(n8874)
         );
  NAND2_X1 U6549 ( .A1(wdata_a_i[20]), .A2(n4744), .ZN(n7880) );
  OAI22_X1 U6550 ( .A1(n1623), .A2(n7881), .B1(n4040), .B2(n4744), .ZN(n8876)
         );
  NAND2_X1 U6551 ( .A1(wdata_a_i[19]), .A2(n4744), .ZN(n7881) );
  OAI22_X1 U6552 ( .A1(n1623), .A2(n7882), .B1(n4444), .B2(n4744), .ZN(n8878)
         );
  NAND2_X1 U6553 ( .A1(wdata_a_i[18]), .A2(n4744), .ZN(n7882) );
  OAI22_X1 U6554 ( .A1(n1623), .A2(n7883), .B1(n4374), .B2(n4744), .ZN(n8880)
         );
  NAND2_X1 U6555 ( .A1(wdata_a_i[17]), .A2(n4744), .ZN(n7883) );
  OAI22_X1 U6556 ( .A1(n1623), .A2(n7884), .B1(n4441), .B2(n4744), .ZN(n8882)
         );
  NAND2_X1 U6557 ( .A1(wdata_a_i[16]), .A2(n4744), .ZN(n7884) );
  OAI22_X1 U6558 ( .A1(n1623), .A2(n7885), .B1(n4439), .B2(n4744), .ZN(n8884)
         );
  NAND2_X1 U6559 ( .A1(wdata_a_i[15]), .A2(n4744), .ZN(n7885) );
  MUX2_X1 U6560 ( .A(wdata_a_i[14]), .B(n8887), .S(n1624), .Z(n8886) );
  MUX2_X1 U6561 ( .A(wdata_a_i[13]), .B(n9174), .S(n1624), .Z(n8888) );
  MUX2_X1 U6562 ( .A(wdata_a_i[12]), .B(n8890), .S(n1624), .Z(n8889) );
  INV_X1 U6563 ( .A(n4432), .ZN(n8890) );
  MUX2_X1 U6564 ( .A(wdata_a_i[11]), .B(n4781), .S(n1624), .Z(n8891) );
  MUX2_X1 U6565 ( .A(wdata_a_i[10]), .B(n9089), .S(n1624), .Z(n8893) );
  MUX2_X1 U6566 ( .A(wdata_a_i[9]), .B(n4783), .S(n1624), .Z(n8895) );
  INV_X1 U6567 ( .A(n4426), .ZN(n8896) );
  MUX2_X1 U6568 ( .A(wdata_a_i[8]), .B(n8898), .S(n1624), .Z(n8897) );
  MUX2_X1 U6569 ( .A(n4486), .B(wdata_b_i[7]), .S(n1624), .Z(n8899) );
  MUX2_X1 U6570 ( .A(wdata_a_i[6]), .B(n4420), .S(n1624), .Z(n8900) );
  OAI22_X1 U6571 ( .A1(n1623), .A2(n7886), .B1(n4418), .B2(n4744), .ZN(n8901)
         );
  NAND2_X1 U6572 ( .A1(wdata_a_i[5]), .A2(n4744), .ZN(n7886) );
  INV_X1 U6573 ( .A(n4418), .ZN(n8902) );
  OAI22_X1 U6574 ( .A1(n1623), .A2(n7887), .B1(n4416), .B2(n4744), .ZN(n8903)
         );
  NAND2_X1 U6575 ( .A1(wdata_a_i[4]), .A2(n4744), .ZN(n7887) );
  MUX2_X1 U6576 ( .A(wdata_a_i[3]), .B(n9100), .S(n1624), .Z(n8905) );
  OAI22_X1 U6577 ( .A1(n1623), .A2(n7888), .B1(n4412), .B2(n4744), .ZN(n8907)
         );
  NAND2_X1 U6578 ( .A1(wdata_a_i[2]), .A2(n4744), .ZN(n7888) );
  INV_X1 U6579 ( .A(n4412), .ZN(n8908) );
  OAI22_X1 U6580 ( .A1(n1623), .A2(n7889), .B1(n4410), .B2(n4744), .ZN(n8909)
         );
  NAND2_X1 U6581 ( .A1(wdata_a_i[1]), .A2(n4744), .ZN(n7889) );
  INV_X1 U6582 ( .A(n7890), .ZN(n8911) );
  AOI22_X1 U6583 ( .A1(wdata_a_i[0]), .A2(n7891), .B1(n1624), .B2(n9195), .ZN(
        n7890) );
  NOR2_X1 U6584 ( .A1(n1623), .A2(n1624), .ZN(n7891) );
  OR2_X1 U6585 ( .A1(n1625), .A2(n1624), .ZN(n8914) );
  NOR2_X1 U6586 ( .A1(n2469), .A2(n4823), .ZN(n7892) );
  NOR2_X1 U6587 ( .A1(n2469), .A2(n4823), .ZN(n7893) );
  INV_X1 U6588 ( .A(n7894), .ZN(n8918) );
  AOI22_X1 U6589 ( .A1(n4618), .A2(n7896), .B1(n4823), .B2(wdata_b_i[28]), 
        .ZN(n7894) );
  INV_X1 U6590 ( .A(n7895), .ZN(n8919) );
  AOI22_X1 U6591 ( .A1(wdata_a_i[27]), .A2(n7896), .B1(n4823), .B2(n8865), 
        .ZN(n7895) );
  NOR2_X1 U6592 ( .A1(n2469), .A2(n4823), .ZN(n7896) );
  INV_X1 U6593 ( .A(n7897), .ZN(n8920) );
  AOI22_X1 U6594 ( .A1(wdata_a_i[26]), .A2(n7899), .B1(n4823), .B2(n9152), 
        .ZN(n7897) );
  INV_X1 U6595 ( .A(n7898), .ZN(n8921) );
  AOI22_X1 U6596 ( .A1(n4614), .A2(n7899), .B1(n4823), .B2(wdata_b_i[25]), 
        .ZN(n7898) );
  NOR2_X1 U6597 ( .A1(n2469), .A2(n4823), .ZN(n7899) );
  OAI22_X1 U6598 ( .A1(n2469), .A2(n7900), .B1(n4047), .B2(n4750), .ZN(n8922)
         );
  NAND2_X1 U6599 ( .A1(wdata_a_i[24]), .A2(n4750), .ZN(n7900) );
  NOR2_X1 U6600 ( .A1(n2469), .A2(n4823), .ZN(n7901) );
  NOR2_X1 U6601 ( .A1(n2469), .A2(n4823), .ZN(n7902) );
  NOR2_X1 U6602 ( .A1(n2469), .A2(n4823), .ZN(n7903) );
  INV_X1 U6603 ( .A(n7904), .ZN(n8931) );
  AOI22_X1 U6604 ( .A1(wdata_a_i[16]), .A2(n7905), .B1(n4823), .B2(n8349), 
        .ZN(n7904) );
  NOR2_X1 U6605 ( .A1(n2469), .A2(n4823), .ZN(n7905) );
  MUX2_X1 U6606 ( .A(wdata_a_i[14]), .B(n9172), .S(n4823), .Z(n8933) );
  MUX2_X1 U6607 ( .A(wdata_a_i[13]), .B(n9174), .S(n4823), .Z(n8934) );
  MUX2_X1 U6608 ( .A(wdata_a_i[12]), .B(n9085), .S(n4823), .Z(n8935) );
  MUX2_X1 U6609 ( .A(wdata_a_i[11]), .B(n9087), .S(n4823), .Z(n8936) );
  MUX2_X1 U6610 ( .A(wdata_a_i[10]), .B(n9089), .S(n4823), .Z(n8937) );
  MUX2_X1 U6611 ( .A(wdata_a_i[9]), .B(n4783), .S(n4823), .Z(n8938) );
  MUX2_X1 U6612 ( .A(wdata_a_i[8]), .B(n4774), .S(n4823), .Z(n8939) );
  MUX2_X1 U6613 ( .A(wdata_a_i[7]), .B(wdata_b_i[7]), .S(n4823), .Z(n8940) );
  MUX2_X1 U6614 ( .A(wdata_a_i[6]), .B(n4420), .S(n4823), .Z(n8941) );
  INV_X1 U6615 ( .A(n7906), .ZN(n8942) );
  AOI22_X1 U6616 ( .A1(wdata_a_i[5]), .A2(n7907), .B1(n4823), .B2(n8902), .ZN(
        n7906) );
  NOR2_X1 U6617 ( .A1(n2469), .A2(n4823), .ZN(n7907) );
  INV_X1 U6618 ( .A(n7908), .ZN(n8943) );
  AOI22_X1 U6619 ( .A1(wdata_a_i[4]), .A2(n7910), .B1(n4823), .B2(n9098), .ZN(
        n7908) );
  MUX2_X1 U6620 ( .A(wdata_a_i[3]), .B(n9100), .S(n4823), .Z(n8944) );
  INV_X1 U6621 ( .A(n7909), .ZN(n8945) );
  AOI22_X1 U6622 ( .A1(wdata_a_i[2]), .A2(n7910), .B1(n4823), .B2(n9102), .ZN(
        n7909) );
  NOR2_X1 U6623 ( .A1(n2469), .A2(n4823), .ZN(n7910) );
  INV_X1 U6624 ( .A(n7911), .ZN(n8946) );
  AOI22_X1 U6625 ( .A1(wdata_a_i[1]), .A2(n7913), .B1(n4823), .B2(n9104), .ZN(
        n7911) );
  INV_X1 U6626 ( .A(n7912), .ZN(n8947) );
  AOI22_X1 U6627 ( .A1(wdata_a_i[0]), .A2(n7913), .B1(n4823), .B2(n4791), .ZN(
        n7912) );
  NOR2_X1 U6628 ( .A1(n2469), .A2(n4823), .ZN(n7913) );
  NAND2_X1 U6629 ( .A1(n2469), .A2(n4750), .ZN(n8950) );
  NOR2_X1 U6630 ( .A1(n2528), .A2(n4814), .ZN(n7914) );
  MUX2_X1 U6631 ( .A(wdata_a_i[29]), .B(n4803), .S(n4814), .Z(n8953) );
  MUX2_X1 U6632 ( .A(wdata_a_i[28]), .B(wdata_b_i[28]), .S(n4814), .Z(n8954)
         );
  MUX2_X1 U6633 ( .A(wdata_a_i[27]), .B(n8865), .S(n4814), .Z(n8955) );
  MUX2_X1 U6634 ( .A(wdata_a_i[26]), .B(n9152), .S(n4814), .Z(n8956) );
  MUX2_X1 U6635 ( .A(wdata_a_i[25]), .B(wdata_b_i[25]), .S(n4814), .Z(n8957)
         );
  MUX2_X1 U6636 ( .A(wdata_a_i[24]), .B(n9155), .S(n4814), .Z(n8958) );
  NOR2_X1 U6637 ( .A1(n2528), .A2(n4814), .ZN(n7915) );
  MUX2_X1 U6638 ( .A(wdata_a_i[20]), .B(n9072), .S(n4814), .Z(n8962) );
  NOR2_X1 U6639 ( .A1(n2528), .A2(n4814), .ZN(n7916) );
  NOR2_X1 U6640 ( .A1(n2528), .A2(n4814), .ZN(n7917) );
  INV_X1 U6641 ( .A(n7918), .ZN(n8966) );
  AOI22_X1 U6642 ( .A1(wdata_a_i[16]), .A2(n7919), .B1(n4814), .B2(n8349), 
        .ZN(n7918) );
  NOR2_X1 U6643 ( .A1(n2528), .A2(n4814), .ZN(n7919) );
  MUX2_X1 U6644 ( .A(wdata_a_i[14]), .B(n9172), .S(n4814), .Z(n8968) );
  MUX2_X1 U6645 ( .A(wdata_a_i[13]), .B(n9174), .S(n4814), .Z(n8969) );
  MUX2_X1 U6646 ( .A(wdata_a_i[12]), .B(n9085), .S(n4814), .Z(n8970) );
  INV_X1 U6647 ( .A(n7920), .ZN(n8971) );
  AOI22_X1 U6648 ( .A1(wdata_a_i[11]), .A2(n7921), .B1(n4814), .B2(n9087), 
        .ZN(n7920) );
  NOR2_X1 U6649 ( .A1(n2528), .A2(n4814), .ZN(n7921) );
  INV_X1 U6650 ( .A(n7922), .ZN(n8973) );
  AOI22_X1 U6651 ( .A1(wdata_a_i[9]), .A2(n7924), .B1(n4814), .B2(n9091), .ZN(
        n7922) );
  INV_X1 U6652 ( .A(n7923), .ZN(n8974) );
  AOI22_X1 U6653 ( .A1(wdata_a_i[8]), .A2(n7924), .B1(n4814), .B2(n4774), .ZN(
        n7923) );
  NOR2_X1 U6654 ( .A1(n2528), .A2(n4814), .ZN(n7924) );
  INV_X1 U6655 ( .A(n7925), .ZN(n8975) );
  AOI22_X1 U6656 ( .A1(wdata_a_i[7]), .A2(n7927), .B1(n4814), .B2(n8848), .ZN(
        n7925) );
  INV_X1 U6657 ( .A(n7926), .ZN(n8976) );
  AOI22_X1 U6658 ( .A1(wdata_a_i[6]), .A2(n7927), .B1(n4814), .B2(n4420), .ZN(
        n7926) );
  NOR2_X1 U6659 ( .A1(n2528), .A2(n4814), .ZN(n7927) );
  INV_X1 U6660 ( .A(n7928), .ZN(n8977) );
  AOI22_X1 U6661 ( .A1(wdata_a_i[5]), .A2(n7930), .B1(n4814), .B2(n9096), .ZN(
        n7928) );
  INV_X1 U6662 ( .A(n7929), .ZN(n8978) );
  AOI22_X1 U6663 ( .A1(wdata_a_i[4]), .A2(n7930), .B1(n4814), .B2(n9098), .ZN(
        n7929) );
  NOR2_X1 U6664 ( .A1(n2528), .A2(n4814), .ZN(n7930) );
  INV_X1 U6665 ( .A(n7931), .ZN(n8979) );
  AOI22_X1 U6666 ( .A1(wdata_a_i[3]), .A2(n7933), .B1(n4814), .B2(n8906), .ZN(
        n7931) );
  INV_X1 U6667 ( .A(n7932), .ZN(n8980) );
  AOI22_X1 U6668 ( .A1(wdata_a_i[2]), .A2(n7933), .B1(n4814), .B2(n9102), .ZN(
        n7932) );
  NOR2_X1 U6669 ( .A1(n2528), .A2(n4814), .ZN(n7933) );
  INV_X1 U6670 ( .A(n7934), .ZN(n8981) );
  AOI22_X1 U6671 ( .A1(wdata_a_i[1]), .A2(n7936), .B1(n4814), .B2(n9104), .ZN(
        n7934) );
  INV_X1 U6672 ( .A(n7935), .ZN(n8982) );
  AOI22_X1 U6673 ( .A1(wdata_a_i[0]), .A2(n7936), .B1(n4814), .B2(n4790), .ZN(
        n7935) );
  NOR2_X1 U6674 ( .A1(n2528), .A2(n4814), .ZN(n7936) );
  OR2_X1 U6675 ( .A1(n2530), .A2(n4814), .ZN(n8985) );
  NOR2_X1 U6676 ( .A1(n2542), .A2(n4826), .ZN(n7937) );
  INV_X1 U6677 ( .A(n7938), .ZN(n8989) );
  AOI22_X1 U6678 ( .A1(wdata_a_i[28]), .A2(n7939), .B1(n4826), .B2(
        wdata_b_i[28]), .ZN(n7938) );
  NOR2_X1 U6679 ( .A1(n2542), .A2(n4826), .ZN(n7939) );
  INV_X1 U6680 ( .A(n7940), .ZN(n8990) );
  AOI22_X1 U6681 ( .A1(wdata_a_i[27]), .A2(n7942), .B1(n4826), .B2(n4732), 
        .ZN(n7940) );
  INV_X1 U6682 ( .A(n7941), .ZN(n8991) );
  AOI22_X1 U6683 ( .A1(wdata_a_i[26]), .A2(n7942), .B1(n4826), .B2(n8867), 
        .ZN(n7941) );
  NOR2_X1 U6684 ( .A1(n2542), .A2(n4826), .ZN(n7942) );
  INV_X1 U6685 ( .A(n7943), .ZN(n8992) );
  AOI22_X1 U6686 ( .A1(wdata_a_i[25]), .A2(n7945), .B1(n4826), .B2(
        wdata_b_i[25]), .ZN(n7943) );
  INV_X1 U6687 ( .A(n7944), .ZN(n8993) );
  AOI22_X1 U6688 ( .A1(wdata_a_i[24]), .A2(n7945), .B1(n4826), .B2(n9155), 
        .ZN(n7944) );
  NOR2_X1 U6689 ( .A1(n2542), .A2(n4826), .ZN(n7945) );
  NOR2_X1 U6690 ( .A1(n2542), .A2(n4826), .ZN(n7946) );
  NOR2_X1 U6691 ( .A1(n2542), .A2(n4826), .ZN(n7947) );
  NOR2_X1 U6692 ( .A1(n2542), .A2(n4826), .ZN(n7948) );
  INV_X1 U6693 ( .A(n7949), .ZN(n9001) );
  AOI22_X1 U6694 ( .A1(wdata_a_i[16]), .A2(n7950), .B1(n4826), .B2(n8349), 
        .ZN(n7949) );
  NOR2_X1 U6695 ( .A1(n2542), .A2(n4826), .ZN(n7950) );
  MUX2_X1 U6696 ( .A(wdata_a_i[14]), .B(n9172), .S(n4826), .Z(n9003) );
  MUX2_X1 U6697 ( .A(wdata_a_i[13]), .B(n9174), .S(n4826), .Z(n9004) );
  MUX2_X1 U6698 ( .A(wdata_a_i[12]), .B(n9085), .S(n4826), .Z(n9005) );
  MUX2_X1 U6699 ( .A(wdata_a_i[11]), .B(n9087), .S(n4826), .Z(n9006) );
  MUX2_X1 U6700 ( .A(wdata_a_i[10]), .B(n9089), .S(n4826), .Z(n9007) );
  MUX2_X1 U6701 ( .A(wdata_a_i[9]), .B(n4783), .S(n4826), .Z(n9008) );
  MUX2_X1 U6702 ( .A(wdata_a_i[8]), .B(n4774), .S(n4826), .Z(n9009) );
  MUX2_X1 U6703 ( .A(wdata_a_i[7]), .B(wdata_b_i[7]), .S(n4826), .Z(n9010) );
  MUX2_X1 U6704 ( .A(wdata_a_i[6]), .B(n4420), .S(n4826), .Z(n9011) );
  INV_X1 U6705 ( .A(n7951), .ZN(n9012) );
  AOI22_X1 U6706 ( .A1(wdata_a_i[5]), .A2(n7952), .B1(n4826), .B2(n9096), .ZN(
        n7951) );
  NOR2_X1 U6707 ( .A1(n2542), .A2(n4826), .ZN(n7952) );
  INV_X1 U6708 ( .A(n7953), .ZN(n9013) );
  AOI22_X1 U6709 ( .A1(wdata_a_i[4]), .A2(n7955), .B1(n4826), .B2(n9098), .ZN(
        n7953) );
  MUX2_X1 U6710 ( .A(wdata_a_i[3]), .B(n8906), .S(n4826), .Z(n9014) );
  INV_X1 U6711 ( .A(n7954), .ZN(n9015) );
  AOI22_X1 U6712 ( .A1(wdata_a_i[2]), .A2(n7955), .B1(n4826), .B2(n9102), .ZN(
        n7954) );
  NOR2_X1 U6713 ( .A1(n2542), .A2(n4826), .ZN(n7955) );
  INV_X1 U6714 ( .A(n7956), .ZN(n9016) );
  AOI22_X1 U6715 ( .A1(wdata_a_i[1]), .A2(n7958), .B1(n4826), .B2(n9104), .ZN(
        n7956) );
  INV_X1 U6716 ( .A(n7957), .ZN(n9017) );
  AOI22_X1 U6717 ( .A1(wdata_a_i[0]), .A2(n7958), .B1(n4826), .B2(n4791), .ZN(
        n7957) );
  NOR2_X1 U6718 ( .A1(n2542), .A2(n4826), .ZN(n7958) );
  NAND2_X1 U6719 ( .A1(n2542), .A2(n4753), .ZN(n9020) );
  NOR2_X1 U6720 ( .A1(n2550), .A2(n4813), .ZN(n7959) );
  MUX2_X1 U6721 ( .A(wdata_a_i[29]), .B(n4803), .S(n4813), .Z(n9023) );
  MUX2_X1 U6722 ( .A(wdata_a_i[28]), .B(wdata_b_i[28]), .S(n4813), .Z(n9024)
         );
  MUX2_X1 U6723 ( .A(wdata_a_i[27]), .B(n4732), .S(n4813), .Z(n9025) );
  MUX2_X1 U6724 ( .A(wdata_a_i[26]), .B(n8867), .S(n4813), .Z(n9026) );
  MUX2_X1 U6725 ( .A(wdata_a_i[25]), .B(wdata_b_i[25]), .S(n4813), .Z(n9027)
         );
  MUX2_X1 U6726 ( .A(wdata_a_i[24]), .B(wdata_b_i[24]), .S(n4813), .Z(n9028)
         );
  NOR2_X1 U6727 ( .A1(n2550), .A2(n4813), .ZN(n7960) );
  OAI22_X1 U6728 ( .A1(n2550), .A2(n7961), .B1(n4449), .B2(n4760), .ZN(n9031)
         );
  NAND2_X1 U6729 ( .A1(wdata_a_i[21]), .A2(n4760), .ZN(n7961) );
  INV_X1 U6730 ( .A(n4449), .ZN(n9032) );
  MUX2_X1 U6731 ( .A(wdata_a_i[20]), .B(n9072), .S(n4813), .Z(n9033) );
  NOR2_X1 U6732 ( .A1(n2550), .A2(n4813), .ZN(n7962) );
  NOR2_X1 U6733 ( .A1(n2550), .A2(n4813), .ZN(n7963) );
  INV_X1 U6734 ( .A(n7964), .ZN(n9037) );
  AOI22_X1 U6735 ( .A1(wdata_a_i[16]), .A2(n7965), .B1(n4813), .B2(n8349), 
        .ZN(n7964) );
  NOR2_X1 U6736 ( .A1(n2550), .A2(n4813), .ZN(n7965) );
  MUX2_X1 U6737 ( .A(wdata_a_i[14]), .B(n9172), .S(n4813), .Z(n9039) );
  MUX2_X1 U6738 ( .A(wdata_a_i[13]), .B(n9174), .S(n4813), .Z(n9040) );
  MUX2_X1 U6739 ( .A(wdata_a_i[12]), .B(n9085), .S(n4813), .Z(n9041) );
  INV_X1 U6740 ( .A(n7966), .ZN(n9042) );
  AOI22_X1 U6741 ( .A1(wdata_a_i[11]), .A2(n7967), .B1(n4813), .B2(n9087), 
        .ZN(n7966) );
  NOR2_X1 U6742 ( .A1(n2550), .A2(n4813), .ZN(n7967) );
  INV_X1 U6743 ( .A(n7968), .ZN(n9044) );
  AOI22_X1 U6744 ( .A1(wdata_a_i[9]), .A2(n7970), .B1(n4813), .B2(n4783), .ZN(
        n7968) );
  INV_X1 U6745 ( .A(n7969), .ZN(n9045) );
  AOI22_X1 U6746 ( .A1(wdata_a_i[8]), .A2(n7970), .B1(n4813), .B2(n4774), .ZN(
        n7969) );
  NOR2_X1 U6747 ( .A1(n2550), .A2(n4813), .ZN(n7970) );
  INV_X1 U6748 ( .A(n7971), .ZN(n9046) );
  AOI22_X1 U6749 ( .A1(n4486), .A2(n7973), .B1(n4813), .B2(n9182), .ZN(n7971)
         );
  INV_X1 U6750 ( .A(n7972), .ZN(n9047) );
  AOI22_X1 U6751 ( .A1(wdata_a_i[6]), .A2(n7973), .B1(n4813), .B2(n4420), .ZN(
        n7972) );
  NOR2_X1 U6752 ( .A1(n2550), .A2(n4813), .ZN(n7973) );
  INV_X1 U6753 ( .A(n7974), .ZN(n9048) );
  AOI22_X1 U6754 ( .A1(wdata_a_i[5]), .A2(n7976), .B1(n4813), .B2(n8902), .ZN(
        n7974) );
  INV_X1 U6755 ( .A(n7975), .ZN(n9049) );
  AOI22_X1 U6756 ( .A1(wdata_a_i[4]), .A2(n7976), .B1(n4813), .B2(n9098), .ZN(
        n7975) );
  NOR2_X1 U6757 ( .A1(n2550), .A2(n4813), .ZN(n7976) );
  INV_X1 U6758 ( .A(n7977), .ZN(n9050) );
  AOI22_X1 U6759 ( .A1(wdata_a_i[3]), .A2(n7979), .B1(n4813), .B2(n9100), .ZN(
        n7977) );
  INV_X1 U6760 ( .A(n7978), .ZN(n9051) );
  AOI22_X1 U6761 ( .A1(wdata_a_i[2]), .A2(n7979), .B1(n4813), .B2(n9102), .ZN(
        n7978) );
  NOR2_X1 U6762 ( .A1(n2550), .A2(n4813), .ZN(n7979) );
  INV_X1 U6763 ( .A(n7980), .ZN(n9052) );
  AOI22_X1 U6764 ( .A1(wdata_a_i[1]), .A2(n7982), .B1(n4813), .B2(n9104), .ZN(
        n7980) );
  INV_X1 U6765 ( .A(n7981), .ZN(n9053) );
  AOI22_X1 U6766 ( .A1(wdata_a_i[0]), .A2(n7982), .B1(n4813), .B2(n4790), .ZN(
        n7981) );
  NOR2_X1 U6767 ( .A1(n2550), .A2(n4813), .ZN(n7982) );
  OR2_X1 U6768 ( .A1(n4813), .A2(n2551), .ZN(n9056) );
  OAI22_X1 U6769 ( .A1(n2474), .A2(n7983), .B1(n4474), .B2(n7984), .ZN(n9057)
         );
  NAND2_X1 U6770 ( .A1(n4477), .A2(n7984), .ZN(n7983) );
  INV_X1 U6771 ( .A(n4824), .ZN(n7984) );
  OAI22_X1 U6772 ( .A1(n2474), .A2(n7985), .B1(n4470), .B2(n7984), .ZN(n9058)
         );
  NAND2_X1 U6773 ( .A1(n4472), .A2(n7984), .ZN(n7985) );
  NOR2_X1 U6774 ( .A1(n2474), .A2(n4824), .ZN(n7986) );
  INV_X1 U6775 ( .A(n7987), .ZN(n9060) );
  AOI22_X1 U6776 ( .A1(n4618), .A2(n7991), .B1(n4824), .B2(wdata_b_i[28]), 
        .ZN(n7987) );
  OAI22_X1 U6777 ( .A1(n2474), .A2(n7988), .B1(n4795), .B2(n4754), .ZN(n9061)
         );
  NAND2_X1 U6778 ( .A1(n4394), .A2(n7984), .ZN(n7988) );
  OAI22_X1 U6779 ( .A1(n2474), .A2(n7989), .B1(n4458), .B2(n4754), .ZN(n9062)
         );
  NAND2_X1 U6780 ( .A1(n4459), .A2(n7984), .ZN(n7989) );
  INV_X1 U6781 ( .A(n4458), .ZN(n9063) );
  INV_X1 U6782 ( .A(n7990), .ZN(n9064) );
  AOI22_X1 U6783 ( .A1(n4614), .A2(n7991), .B1(n4824), .B2(wdata_b_i[25]), 
        .ZN(n7990) );
  NOR2_X1 U6784 ( .A1(n2474), .A2(n4824), .ZN(n7991) );
  OAI22_X1 U6785 ( .A1(n2474), .A2(n7992), .B1(n4047), .B2(n4754), .ZN(n9065)
         );
  NAND2_X1 U6786 ( .A1(n4386), .A2(n4754), .ZN(n7992) );
  OAI22_X1 U6787 ( .A1(n2474), .A2(n7993), .B1(n4385), .B2(n4754), .ZN(n9066)
         );
  NAND2_X1 U6788 ( .A1(wdata_a_i[23]), .A2(n4754), .ZN(n7993) );
  OAI22_X1 U6789 ( .A1(n2474), .A2(n7994), .B1(n4004), .B2(n7984), .ZN(n9067)
         );
  NAND2_X1 U6790 ( .A1(wdata_a_i[22]), .A2(n4754), .ZN(n7994) );
  OAI22_X1 U6791 ( .A1(n2474), .A2(n7995), .B1(n4449), .B2(n4754), .ZN(n9069)
         );
  NAND2_X1 U6792 ( .A1(wdata_a_i[21]), .A2(n4754), .ZN(n7995) );
  OAI22_X1 U6793 ( .A1(n2474), .A2(n7996), .B1(n4002), .B2(n7984), .ZN(n9071)
         );
  NAND2_X1 U6794 ( .A1(wdata_a_i[20]), .A2(n4754), .ZN(n7996) );
  OAI22_X1 U6795 ( .A1(n2474), .A2(n7997), .B1(n4040), .B2(n4754), .ZN(n9073)
         );
  NAND2_X1 U6796 ( .A1(wdata_a_i[19]), .A2(n7984), .ZN(n7997) );
  OAI22_X1 U6797 ( .A1(n2474), .A2(n7998), .B1(n4444), .B2(n4754), .ZN(n9075)
         );
  NAND2_X1 U6798 ( .A1(wdata_a_i[18]), .A2(n4754), .ZN(n7998) );
  OAI22_X1 U6799 ( .A1(n2474), .A2(n7999), .B1(n4374), .B2(n4754), .ZN(n9077)
         );
  NAND2_X1 U6800 ( .A1(wdata_a_i[17]), .A2(n4754), .ZN(n7999) );
  INV_X1 U6801 ( .A(n4037), .ZN(n9078) );
  INV_X1 U6802 ( .A(n8000), .ZN(n9079) );
  AOI22_X1 U6803 ( .A1(wdata_a_i[16]), .A2(n8007), .B1(n4824), .B2(n8349), 
        .ZN(n8000) );
  OAI22_X1 U6804 ( .A1(n2474), .A2(n8001), .B1(n4439), .B2(n4754), .ZN(n9080)
         );
  NAND2_X1 U6805 ( .A1(wdata_a_i[15]), .A2(n7984), .ZN(n8001) );
  MUX2_X1 U6806 ( .A(wdata_a_i[14]), .B(n9172), .S(n4824), .Z(n9082) );
  MUX2_X1 U6807 ( .A(wdata_a_i[13]), .B(n9174), .S(n4824), .Z(n9083) );
  MUX2_X1 U6808 ( .A(wdata_a_i[12]), .B(n9085), .S(n4824), .Z(n9084) );
  MUX2_X1 U6809 ( .A(wdata_a_i[11]), .B(n9087), .S(n4824), .Z(n9086) );
  INV_X1 U6810 ( .A(n4430), .ZN(n9087) );
  MUX2_X1 U6811 ( .A(wdata_a_i[10]), .B(n9089), .S(n4824), .Z(n9088) );
  INV_X1 U6812 ( .A(n4798), .ZN(n9089) );
  MUX2_X1 U6813 ( .A(wdata_a_i[9]), .B(n4783), .S(n4824), .Z(n9090) );
  MUX2_X1 U6814 ( .A(wdata_a_i[8]), .B(n4774), .S(n4824), .Z(n9092) );
  MUX2_X1 U6815 ( .A(wdata_a_i[7]), .B(wdata_b_i[7]), .S(n4824), .Z(n9093) );
  MUX2_X1 U6816 ( .A(wdata_a_i[6]), .B(n4420), .S(n4824), .Z(n9094) );
  OAI22_X1 U6817 ( .A1(n2474), .A2(n8002), .B1(n4418), .B2(n7984), .ZN(n9095)
         );
  NAND2_X1 U6818 ( .A1(wdata_a_i[5]), .A2(n7984), .ZN(n8002) );
  INV_X1 U6819 ( .A(n4418), .ZN(n9096) );
  OAI22_X1 U6820 ( .A1(n2474), .A2(n8003), .B1(n4416), .B2(n4754), .ZN(n9097)
         );
  NAND2_X1 U6821 ( .A1(wdata_a_i[4]), .A2(n4754), .ZN(n8003) );
  INV_X1 U6822 ( .A(n4416), .ZN(n9098) );
  MUX2_X1 U6823 ( .A(wdata_a_i[3]), .B(n8906), .S(n4824), .Z(n9099) );
  INV_X1 U6824 ( .A(n4414), .ZN(n9100) );
  OAI22_X1 U6825 ( .A1(n2474), .A2(n8004), .B1(n4412), .B2(n4754), .ZN(n9101)
         );
  NAND2_X1 U6826 ( .A1(wdata_a_i[2]), .A2(n7984), .ZN(n8004) );
  INV_X1 U6827 ( .A(n4412), .ZN(n9102) );
  OAI22_X1 U6828 ( .A1(n2474), .A2(n8005), .B1(n4410), .B2(n4754), .ZN(n9103)
         );
  NAND2_X1 U6829 ( .A1(wdata_a_i[1]), .A2(n4754), .ZN(n8005) );
  INV_X1 U6830 ( .A(n4410), .ZN(n9104) );
  INV_X1 U6831 ( .A(n8006), .ZN(n9105) );
  AOI22_X1 U6832 ( .A1(wdata_a_i[0]), .A2(n8007), .B1(n4824), .B2(n9195), .ZN(
        n8006) );
  NOR2_X1 U6833 ( .A1(n2474), .A2(n4824), .ZN(n8007) );
  NAND2_X1 U6834 ( .A1(n2474), .A2(n4754), .ZN(n9108) );
  NOR2_X1 U6835 ( .A1(n1604), .A2(n4818), .ZN(n8008) );
  MUX2_X1 U6836 ( .A(n4468), .B(n4803), .S(n4818), .Z(n9111) );
  MUX2_X1 U6837 ( .A(n4618), .B(wdata_b_i[28]), .S(n4818), .Z(n9112) );
  MUX2_X1 U6838 ( .A(n4394), .B(n4732), .S(n4818), .Z(n9113) );
  MUX2_X1 U6839 ( .A(n4459), .B(n8867), .S(n4818), .Z(n9114) );
  MUX2_X1 U6840 ( .A(n4614), .B(wdata_b_i[25]), .S(n4818), .Z(n9115) );
  MUX2_X1 U6841 ( .A(n4386), .B(n9155), .S(n4818), .Z(n9116) );
  NOR2_X1 U6842 ( .A1(n1604), .A2(n4818), .ZN(n8009) );
  NOR2_X1 U6843 ( .A1(n1604), .A2(n4818), .ZN(n8010) );
  NOR2_X1 U6844 ( .A1(n1604), .A2(n4818), .ZN(n8011) );
  MUX2_X1 U6845 ( .A(wdata_a_i[16]), .B(n8349), .S(n4818), .Z(n9124) );
  NOR2_X1 U6846 ( .A1(n1604), .A2(n4818), .ZN(n8012) );
  MUX2_X1 U6847 ( .A(wdata_a_i[14]), .B(n9172), .S(n4818), .Z(n9126) );
  MUX2_X1 U6848 ( .A(wdata_a_i[13]), .B(n9174), .S(n4818), .Z(n9127) );
  MUX2_X1 U6849 ( .A(wdata_a_i[12]), .B(n9085), .S(n4818), .Z(n9128) );
  INV_X1 U6850 ( .A(n8013), .ZN(n9129) );
  AOI22_X1 U6851 ( .A1(wdata_a_i[11]), .A2(n8014), .B1(n4818), .B2(n4782), 
        .ZN(n8013) );
  NOR2_X1 U6852 ( .A1(n1604), .A2(n4818), .ZN(n8014) );
  INV_X1 U6853 ( .A(n8015), .ZN(n9131) );
  AOI22_X1 U6854 ( .A1(wdata_a_i[9]), .A2(n8017), .B1(n4818), .B2(n9091), .ZN(
        n8015) );
  INV_X1 U6855 ( .A(n8016), .ZN(n9132) );
  AOI22_X1 U6856 ( .A1(wdata_a_i[8]), .A2(n8017), .B1(n4818), .B2(n8898), .ZN(
        n8016) );
  NOR2_X1 U6857 ( .A1(n1604), .A2(n4818), .ZN(n8017) );
  INV_X1 U6858 ( .A(n8018), .ZN(n9133) );
  AOI22_X1 U6859 ( .A1(n4486), .A2(n8020), .B1(n4818), .B2(n4780), .ZN(n8018)
         );
  INV_X1 U6860 ( .A(n8019), .ZN(n9134) );
  AOI22_X1 U6861 ( .A1(wdata_a_i[6]), .A2(n8020), .B1(n4818), .B2(n9184), .ZN(
        n8019) );
  NOR2_X1 U6862 ( .A1(n1604), .A2(n4818), .ZN(n8020) );
  INV_X1 U6863 ( .A(n8021), .ZN(n9135) );
  AOI22_X1 U6864 ( .A1(wdata_a_i[5]), .A2(n8023), .B1(n4818), .B2(n9096), .ZN(
        n8021) );
  INV_X1 U6865 ( .A(n8022), .ZN(n9136) );
  AOI22_X1 U6866 ( .A1(wdata_a_i[4]), .A2(n8023), .B1(n4818), .B2(n4787), .ZN(
        n8022) );
  NOR2_X1 U6867 ( .A1(n1604), .A2(n4818), .ZN(n8023) );
  INV_X1 U6868 ( .A(n8024), .ZN(n9137) );
  AOI22_X1 U6869 ( .A1(wdata_a_i[3]), .A2(n8026), .B1(n4818), .B2(n9100), .ZN(
        n8024) );
  INV_X1 U6870 ( .A(n8025), .ZN(n9138) );
  AOI22_X1 U6871 ( .A1(wdata_a_i[2]), .A2(n8026), .B1(n4818), .B2(n9191), .ZN(
        n8025) );
  NOR2_X1 U6872 ( .A1(n1604), .A2(n4818), .ZN(n8026) );
  INV_X1 U6873 ( .A(n8027), .ZN(n9139) );
  AOI22_X1 U6874 ( .A1(wdata_a_i[1]), .A2(n8029), .B1(n4818), .B2(n4786), .ZN(
        n8027) );
  INV_X1 U6875 ( .A(n8028), .ZN(n9140) );
  AOI22_X1 U6876 ( .A1(wdata_a_i[0]), .A2(n8029), .B1(n4818), .B2(n4791), .ZN(
        n8028) );
  NOR2_X1 U6877 ( .A1(n1604), .A2(n4818), .ZN(n8029) );
  OR2_X1 U6878 ( .A1(n1606), .A2(n4818), .ZN(n9143) );
  OAI22_X1 U6879 ( .A1(n1550), .A2(n8030), .B1(n4474), .B2(n8031), .ZN(n9144)
         );
  NAND2_X1 U6880 ( .A1(n4477), .A2(n8031), .ZN(n8030) );
  INV_X1 U6881 ( .A(n4825), .ZN(n8031) );
  OAI22_X1 U6882 ( .A1(n1550), .A2(n8032), .B1(n4470), .B2(n4748), .ZN(n9145)
         );
  NAND2_X1 U6883 ( .A1(n4472), .A2(n4748), .ZN(n8032) );
  MUX2_X1 U6884 ( .A(n4468), .B(n4803), .S(n4825), .Z(n9147) );
  MUX2_X1 U6885 ( .A(wdata_a_i[28]), .B(wdata_b_i[28]), .S(n4825), .Z(n9148)
         );
  MUX2_X1 U6886 ( .A(n4394), .B(n8865), .S(n4825), .Z(n9149) );
  INV_X1 U6887 ( .A(n4461), .ZN(n9150) );
  MUX2_X1 U6888 ( .A(wdata_a_i[26]), .B(n9152), .S(n4825), .Z(n9151) );
  INV_X1 U6889 ( .A(n4458), .ZN(n9152) );
  MUX2_X1 U6890 ( .A(wdata_a_i[25]), .B(wdata_b_i[25]), .S(n4825), .Z(n9153)
         );
  MUX2_X1 U6891 ( .A(n4386), .B(n9155), .S(n4825), .Z(n9154) );
  OAI22_X1 U6892 ( .A1(n1550), .A2(n8033), .B1(n4385), .B2(n8031), .ZN(n9156)
         );
  NAND2_X1 U6893 ( .A1(wdata_a_i[23]), .A2(n4748), .ZN(n8033) );
  OAI22_X1 U6894 ( .A1(n1550), .A2(n8034), .B1(n4382), .B2(n8031), .ZN(n9158)
         );
  NAND2_X1 U6895 ( .A1(wdata_a_i[22]), .A2(n4748), .ZN(n8034) );
  OAI22_X1 U6896 ( .A1(n1550), .A2(n8035), .B1(n4449), .B2(n8031), .ZN(n9160)
         );
  NAND2_X1 U6897 ( .A1(wdata_a_i[21]), .A2(n4748), .ZN(n8035) );
  OAI22_X1 U6898 ( .A1(n1550), .A2(n8036), .B1(n4002), .B2(n8031), .ZN(n9161)
         );
  NAND2_X1 U6899 ( .A1(wdata_a_i[20]), .A2(n4748), .ZN(n8036) );
  OAI22_X1 U6900 ( .A1(n1550), .A2(n8037), .B1(n4040), .B2(n8031), .ZN(n9163)
         );
  NAND2_X1 U6901 ( .A1(wdata_a_i[19]), .A2(n8031), .ZN(n8037) );
  OAI22_X1 U6902 ( .A1(n1550), .A2(n8038), .B1(n4444), .B2(n4748), .ZN(n9165)
         );
  NAND2_X1 U6903 ( .A1(wdata_a_i[18]), .A2(n4748), .ZN(n8038) );
  OAI22_X1 U6904 ( .A1(n1550), .A2(n8039), .B1(n4374), .B2(n4748), .ZN(n9167)
         );
  NAND2_X1 U6905 ( .A1(wdata_a_i[17]), .A2(n4748), .ZN(n8039) );
  MUX2_X1 U6906 ( .A(wdata_a_i[16]), .B(n8349), .S(n4825), .Z(n9169) );
  OAI22_X1 U6907 ( .A1(n1550), .A2(n8040), .B1(n4439), .B2(n4748), .ZN(n9170)
         );
  NAND2_X1 U6908 ( .A1(wdata_a_i[15]), .A2(n4748), .ZN(n8040) );
  MUX2_X1 U6909 ( .A(wdata_a_i[14]), .B(n9172), .S(n4825), .Z(n9171) );
  MUX2_X1 U6910 ( .A(wdata_a_i[13]), .B(n9174), .S(n4825), .Z(n9173) );
  MUX2_X1 U6911 ( .A(wdata_a_i[12]), .B(n9085), .S(n4825), .Z(n9175) );
  OAI22_X1 U6912 ( .A1(n1550), .A2(n8041), .B1(n4430), .B2(n4748), .ZN(n9176)
         );
  NAND2_X1 U6913 ( .A1(wdata_a_i[11]), .A2(n4748), .ZN(n8041) );
  OAI22_X1 U6914 ( .A1(n1550), .A2(n8042), .B1(n4798), .B2(n4748), .ZN(n9177)
         );
  NAND2_X1 U6915 ( .A1(wdata_a_i[10]), .A2(n8031), .ZN(n8042) );
  OAI22_X1 U6916 ( .A1(n1550), .A2(n8043), .B1(n4426), .B2(n8031), .ZN(n9179)
         );
  NAND2_X1 U6917 ( .A1(wdata_a_i[9]), .A2(n4748), .ZN(n8043) );
  OAI22_X1 U6918 ( .A1(n1550), .A2(n8044), .B1(n4424), .B2(n8031), .ZN(n9180)
         );
  NAND2_X1 U6919 ( .A1(wdata_a_i[8]), .A2(n8031), .ZN(n8044) );
  OAI22_X1 U6920 ( .A1(n1550), .A2(n8045), .B1(n4422), .B2(n8031), .ZN(n9181)
         );
  NAND2_X1 U6921 ( .A1(n4486), .A2(n4748), .ZN(n8045) );
  OAI22_X1 U6922 ( .A1(n1550), .A2(n8046), .B1(n4785), .B2(n8031), .ZN(n9183)
         );
  NAND2_X1 U6923 ( .A1(wdata_a_i[6]), .A2(n8031), .ZN(n8046) );
  OAI22_X1 U6924 ( .A1(n1550), .A2(n8047), .B1(n4418), .B2(n4748), .ZN(n9185)
         );
  NAND2_X1 U6925 ( .A1(wdata_a_i[5]), .A2(n8031), .ZN(n8047) );
  INV_X1 U6926 ( .A(n4418), .ZN(n9186) );
  OAI22_X1 U6927 ( .A1(n1550), .A2(n8048), .B1(n4416), .B2(n8031), .ZN(n9187)
         );
  NAND2_X1 U6928 ( .A1(wdata_a_i[4]), .A2(n8031), .ZN(n8048) );
  OAI22_X1 U6929 ( .A1(n1550), .A2(n8049), .B1(n4414), .B2(n8031), .ZN(n9188)
         );
  NAND2_X1 U6930 ( .A1(wdata_a_i[3]), .A2(n8031), .ZN(n8049) );
  INV_X1 U6931 ( .A(n4414), .ZN(n9189) );
  OAI22_X1 U6932 ( .A1(n1550), .A2(n8050), .B1(n4412), .B2(n8031), .ZN(n9190)
         );
  NAND2_X1 U6933 ( .A1(wdata_a_i[2]), .A2(n4748), .ZN(n8050) );
  OAI22_X1 U6934 ( .A1(n1550), .A2(n8051), .B1(n4410), .B2(n4748), .ZN(n9192)
         );
  NAND2_X1 U6935 ( .A1(wdata_a_i[1]), .A2(n4748), .ZN(n8051) );
  OAI22_X1 U6936 ( .A1(n1550), .A2(n8052), .B1(n4408), .B2(n8031), .ZN(n9194)
         );
  NAND2_X1 U6937 ( .A1(wdata_a_i[0]), .A2(n4748), .ZN(n8052) );
  OR2_X1 U6938 ( .A1(n4825), .A2(n1551), .ZN(n9198) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_prefetch_L0_buffer_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_prefetch_L0_buffer_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_prefetch_L0_buffer_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module riscv_L0_buffer_RDATA_IN_WIDTH128 ( clk, rst_n, prefetch_i, 
        prefetch_addr_i, branch_i, branch_addr_i, hwlp_i, hwlp_addr_i, 
        fetch_gnt_o, fetch_valid_o, valid_o, rdata_o, addr_o, instr_req_o, 
        instr_addr_o, instr_gnt_i, instr_rvalid_i, instr_rdata_i, busy_o );
  input [31:0] prefetch_addr_i;
  input [31:0] branch_addr_i;
  input [31:0] hwlp_addr_i;
  output [127:0] rdata_o;
  output [31:0] addr_o;
  output [31:0] instr_addr_o;
  input [127:0] instr_rdata_i;
  input clk, rst_n, prefetch_i, branch_i, hwlp_i, instr_gnt_i, instr_rvalid_i;
  output fetch_gnt_o, fetch_valid_o, valid_o, instr_req_o, busy_o;
  wire   instr_gnt_i, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n274, n275, n276, n277, n279, n280,
         n281, n283, n284, n288, n289, n290, n31, n34, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n60, n62, n64, n65, n66, n67, n68, n69, n70,
         n71, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n207, n208, n209, n210, n211, n212, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n256, n291, n292, n293, n294, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n306, n307, n308, n309, n310, n311, n313,
         n314, n315, n316, n317, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n367, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n383, n384, n385, n386, n387, n388, n709, n711, n712,
         n713, n714, n716, n717, n718, n719, n720;
  wire   [2:0] CS;
  wire   [112:0] L0_buffer;
  assign fetch_gnt_o = instr_gnt_i;

  INV_X1 U296 ( .A(rst_n) );
  CLKBUF_X1 U3 ( .A(n298), .Z(n31) );
  NOR2_X1 U27 ( .A1(n298), .A2(n96), .ZN(n97) );
  AND2_X2 U29 ( .A1(branch_i), .A2(n79), .ZN(n103) );
  OAI21_X1 U30 ( .B1(instr_rvalid_i), .B2(n351), .A(n333), .ZN(rdata_o[97]) );
  OAI21_X1 U31 ( .B1(instr_rvalid_i), .B2(n353), .A(n78), .ZN(rdata_o[113]) );
  NAND3_X1 U32 ( .A1(n147), .A2(n145), .A3(n146), .ZN(instr_addr_o[29]) );
  NAND3_X1 U33 ( .A1(n65), .A2(n117), .A3(n118), .ZN(instr_addr_o[11]) );
  NAND3_X1 U36 ( .A1(n49), .A2(n133), .A3(n132), .ZN(instr_addr_o[16]) );
  NAND2_X1 U37 ( .A1(branch_addr_i[16]), .A2(n103), .ZN(n49) );
  NAND3_X1 U39 ( .A1(n64), .A2(n164), .A3(n165), .ZN(instr_addr_o[13]) );
  AOI21_X1 U40 ( .B1(prefetch_addr_i[15]), .B2(n307), .A(n50), .ZN(n123) );
  NAND2_X1 U41 ( .A1(n52), .A2(n51), .ZN(n50) );
  NAND2_X1 U42 ( .A1(n314), .A2(hwlp_addr_i[15]), .ZN(n51) );
  NAND2_X1 U43 ( .A1(n163), .A2(n18), .ZN(n52) );
  NAND2_X1 U45 ( .A1(n98), .A2(n53), .ZN(instr_addr_o[20]) );
  AOI21_X1 U46 ( .B1(prefetch_addr_i[20]), .B2(n307), .A(n97), .ZN(n53) );
  AND2_X1 U47 ( .A1(n100), .A2(n99), .ZN(n101) );
  NAND3_X1 U49 ( .A1(n90), .A2(n88), .A3(n89), .ZN(instr_addr_o[21]) );
  AND2_X1 U52 ( .A1(n101), .A2(n102), .ZN(n54) );
  NOR2_X1 U55 ( .A1(branch_i), .A2(n81), .ZN(n106) );
  AOI21_X1 U56 ( .B1(n162), .B2(prefetch_addr_i[10]), .A(n74), .ZN(n73) );
  AND2_X1 U57 ( .A1(n156), .A2(n157), .ZN(n62) );
  AND2_X1 U58 ( .A1(n113), .A2(n112), .ZN(n71) );
  AND2_X1 U59 ( .A1(n108), .A2(n109), .ZN(n110) );
  CLKBUF_X1 U61 ( .A(instr_addr_o[19]), .Z(n236) );
  CLKBUF_X1 U62 ( .A(instr_addr_o[18]), .Z(n233) );
  CLKBUF_X1 U63 ( .A(instr_addr_o[17]), .Z(n230) );
  CLKBUF_X1 U64 ( .A(instr_addr_o[15]), .Z(n224) );
  CLKBUF_X1 U65 ( .A(instr_addr_o[10]), .Z(n212) );
  CLKBUF_X1 U67 ( .A(instr_addr_o[5]), .Z(n201) );
  NOR2_X1 U68 ( .A1(n298), .A2(n139), .ZN(n57) );
  INV_X1 U69 ( .A(instr_addr_o[20]), .ZN(n240) );
  NAND2_X1 U70 ( .A1(prefetch_addr_i[31]), .A2(n307), .ZN(n58) );
  AND3_X1 U72 ( .A1(n69), .A2(n154), .A3(n155), .ZN(n60) );
  NAND2_X1 U73 ( .A1(n158), .A2(n62), .ZN(instr_addr_o[26]) );
  NAND2_X1 U75 ( .A1(branch_addr_i[13]), .A2(n103), .ZN(n64) );
  AND2_X1 U76 ( .A1(n115), .A2(n114), .ZN(n116) );
  NAND2_X1 U77 ( .A1(n140), .A2(n141), .ZN(instr_addr_o[6]) );
  NAND2_X2 U78 ( .A1(n85), .A2(n86), .ZN(instr_addr_o[23]) );
  NAND2_X1 U79 ( .A1(branch_addr_i[11]), .A2(n103), .ZN(n65) );
  NAND3_X1 U80 ( .A1(n136), .A2(n137), .A3(n135), .ZN(instr_addr_o[5]) );
  NAND2_X1 U81 ( .A1(n66), .A2(n116), .ZN(instr_addr_o[14]) );
  NAND2_X1 U82 ( .A1(branch_addr_i[14]), .A2(n153), .ZN(n66) );
  NAND2_X1 U83 ( .A1(n67), .A2(n73), .ZN(instr_addr_o[10]) );
  NAND2_X1 U84 ( .A1(branch_addr_i[10]), .A2(n153), .ZN(n67) );
  NAND2_X1 U85 ( .A1(n68), .A2(n110), .ZN(instr_addr_o[8]) );
  NAND2_X1 U86 ( .A1(branch_addr_i[8]), .A2(n103), .ZN(n68) );
  NAND2_X1 U87 ( .A1(prefetch_addr_i[12]), .A2(n162), .ZN(n70) );
  INV_X1 U89 ( .A(n134), .ZN(n74) );
  NAND2_X1 U90 ( .A1(prefetch_addr_i[18]), .A2(n307), .ZN(n75) );
  INV_X1 U93 ( .A(n379), .ZN(n216) );
  NAND3_X1 U94 ( .A1(n76), .A2(n160), .A3(n161), .ZN(instr_addr_o[25]) );
  NAND2_X1 U95 ( .A1(branch_addr_i[25]), .A2(n159), .ZN(n76) );
  INV_X1 U96 ( .A(instr_addr_o[8]), .ZN(n210) );
  INV_X1 U97 ( .A(n380), .ZN(n291) );
  NAND2_X1 U99 ( .A1(instr_rvalid_i), .A2(instr_rdata_i[112]), .ZN(n77) );
  NAND2_X1 U100 ( .A1(instr_rvalid_i), .A2(instr_rdata_i[113]), .ZN(n78) );
  INV_X1 U101 ( .A(n375), .ZN(n223) );
  AND2_X1 U102 ( .A1(n84), .A2(n83), .ZN(n85) );
  AOI21_X1 U103 ( .B1(n162), .B2(prefetch_addr_i[7]), .A(n120), .ZN(n121) );
  AOI21_X1 U104 ( .B1(prefetch_addr_i[6]), .B2(n307), .A(n57), .ZN(n140) );
  OR2_X1 U105 ( .A1(CS[1]), .A2(CS[0]), .ZN(n190) );
  NAND2_X1 U106 ( .A1(n190), .A2(CS[2]), .ZN(n79) );
  NAND2_X1 U107 ( .A1(branch_addr_i[23]), .A2(n153), .ZN(n86) );
  INV_X1 U108 ( .A(hwlp_i), .ZN(n80) );
  OR2_X1 U109 ( .A1(n336), .A2(CS[0]), .ZN(n178) );
  NAND3_X1 U110 ( .A1(n80), .A2(n337), .A3(n178), .ZN(n81) );
  NAND2_X1 U111 ( .A1(prefetch_addr_i[23]), .A2(n307), .ZN(n84) );
  NAND2_X1 U112 ( .A1(hwlp_i), .A2(n337), .ZN(n95) );
  NOR2_X1 U113 ( .A1(branch_i), .A2(n95), .ZN(n87) );
  NOR2_X1 U114 ( .A1(hwlp_i), .A2(CS[2]), .ZN(n82) );
  NOR2_X1 U115 ( .A1(CS[2]), .A2(CS[1]), .ZN(n180) );
  INV_X1 U116 ( .A(n180), .ZN(n176) );
  OAI211_X1 U117 ( .C1(n82), .C2(n336), .A(n176), .B(n338), .ZN(n94) );
  NOR2_X1 U118 ( .A1(branch_i), .A2(n94), .ZN(n304) );
  AOI22_X1 U119 ( .A1(n314), .A2(hwlp_addr_i[23]), .B1(n166), .B2(n10), .ZN(
        n83) );
  NAND2_X1 U120 ( .A1(branch_addr_i[21]), .A2(n153), .ZN(n90) );
  NAND2_X1 U121 ( .A1(prefetch_addr_i[21]), .A2(n307), .ZN(n89) );
  AOI22_X1 U123 ( .A1(n308), .A2(hwlp_addr_i[21]), .B1(n166), .B2(n12), .ZN(
        n88) );
  NAND2_X1 U124 ( .A1(branch_addr_i[27]), .A2(n159), .ZN(n93) );
  AOI22_X1 U125 ( .A1(n308), .A2(hwlp_addr_i[27]), .B1(n166), .B2(n6), .ZN(n92) );
  NAND2_X1 U126 ( .A1(prefetch_addr_i[27]), .A2(n307), .ZN(n91) );
  NAND3_X1 U127 ( .A1(n93), .A2(n92), .A3(n91), .ZN(instr_addr_o[27]) );
  NAND2_X1 U128 ( .A1(branch_addr_i[20]), .A2(n153), .ZN(n98) );
  INV_X1 U129 ( .A(n94), .ZN(n138) );
  INV_X1 U130 ( .A(n95), .ZN(n182) );
  AOI22_X1 U131 ( .A1(n138), .A2(n13), .B1(n182), .B2(hwlp_addr_i[20]), .ZN(
        n96) );
  NAND2_X1 U133 ( .A1(prefetch_addr_i[30]), .A2(n307), .ZN(n100) );
  AOI22_X1 U134 ( .A1(n314), .A2(hwlp_addr_i[30]), .B1(n166), .B2(n3), .ZN(n99) );
  NAND2_X1 U135 ( .A1(prefetch_addr_i[17]), .A2(n307), .ZN(n105) );
  AOI22_X1 U136 ( .A1(n308), .A2(hwlp_addr_i[17]), .B1(n163), .B2(n16), .ZN(
        n104) );
  AOI22_X1 U137 ( .A1(n314), .A2(hwlp_addr_i[8]), .B1(n163), .B2(n25), .ZN(
        n109) );
  INV_X1 U138 ( .A(n106), .ZN(n107) );
  NAND2_X1 U139 ( .A1(prefetch_addr_i[8]), .A2(n162), .ZN(n108) );
  INV_X1 U140 ( .A(n298), .ZN(n111) );
  NAND3_X1 U141 ( .A1(n111), .A2(n21), .A3(n138), .ZN(n113) );
  NAND3_X1 U142 ( .A1(n111), .A2(n182), .A3(hwlp_addr_i[12]), .ZN(n112) );
  AOI22_X1 U143 ( .A1(n308), .A2(hwlp_addr_i[14]), .B1(n163), .B2(n19), .ZN(
        n115) );
  NAND2_X1 U144 ( .A1(prefetch_addr_i[14]), .A2(n162), .ZN(n114) );
  AOI22_X1 U145 ( .A1(n308), .A2(hwlp_addr_i[11]), .B1(n163), .B2(n22), .ZN(
        n118) );
  NAND2_X1 U146 ( .A1(prefetch_addr_i[11]), .A2(n162), .ZN(n117) );
  NAND2_X1 U147 ( .A1(branch_addr_i[7]), .A2(n153), .ZN(n122) );
  AOI22_X1 U148 ( .A1(n138), .A2(n26), .B1(n182), .B2(hwlp_addr_i[7]), .ZN(
        n119) );
  NOR2_X1 U149 ( .A1(n298), .A2(n119), .ZN(n120) );
  NAND2_X1 U150 ( .A1(n122), .A2(n121), .ZN(instr_addr_o[7]) );
  NAND2_X1 U151 ( .A1(branch_addr_i[15]), .A2(n159), .ZN(n124) );
  NAND2_X1 U152 ( .A1(n124), .A2(n123), .ZN(instr_addr_o[15]) );
  AOI22_X1 U153 ( .A1(n308), .A2(hwlp_addr_i[18]), .B1(n163), .B2(n15), .ZN(
        n125) );
  NAND2_X1 U154 ( .A1(branch_addr_i[4]), .A2(n153), .ZN(n128) );
  NAND2_X1 U155 ( .A1(prefetch_addr_i[4]), .A2(n162), .ZN(n127) );
  AOI22_X1 U156 ( .A1(n308), .A2(hwlp_addr_i[4]), .B1(n163), .B2(n29), .ZN(
        n126) );
  AOI22_X1 U157 ( .A1(n308), .A2(hwlp_addr_i[22]), .B1(n166), .B2(n11), .ZN(
        n130) );
  NAND2_X1 U158 ( .A1(prefetch_addr_i[22]), .A2(n307), .ZN(n129) );
  NAND2_X1 U159 ( .A1(prefetch_addr_i[16]), .A2(n307), .ZN(n133) );
  AOI22_X1 U160 ( .A1(n314), .A2(hwlp_addr_i[16]), .B1(n163), .B2(n17), .ZN(
        n132) );
  AOI22_X1 U161 ( .A1(n87), .A2(hwlp_addr_i[10]), .B1(n304), .B2(n23), .ZN(
        n134) );
  NAND2_X1 U162 ( .A1(branch_addr_i[5]), .A2(n153), .ZN(n137) );
  NAND2_X1 U163 ( .A1(prefetch_addr_i[5]), .A2(n162), .ZN(n136) );
  AOI22_X1 U164 ( .A1(n314), .A2(hwlp_addr_i[5]), .B1(n163), .B2(n28), .ZN(
        n135) );
  NAND2_X1 U165 ( .A1(branch_addr_i[6]), .A2(n103), .ZN(n141) );
  AOI22_X1 U166 ( .A1(n138), .A2(n27), .B1(n182), .B2(hwlp_addr_i[6]), .ZN(
        n139) );
  AOI22_X1 U167 ( .A1(n308), .A2(hwlp_addr_i[19]), .B1(n166), .B2(n14), .ZN(
        n143) );
  NAND2_X1 U168 ( .A1(prefetch_addr_i[19]), .A2(n162), .ZN(n142) );
  NAND2_X1 U169 ( .A1(branch_addr_i[29]), .A2(n153), .ZN(n147) );
  AOI22_X1 U170 ( .A1(n308), .A2(hwlp_addr_i[29]), .B1(n166), .B2(n4), .ZN(
        n146) );
  NAND2_X1 U171 ( .A1(prefetch_addr_i[29]), .A2(n307), .ZN(n145) );
  NAND2_X1 U172 ( .A1(prefetch_addr_i[28]), .A2(n307), .ZN(n149) );
  AOI22_X1 U173 ( .A1(n314), .A2(hwlp_addr_i[28]), .B1(n166), .B2(n5), .ZN(
        n148) );
  NAND2_X1 U174 ( .A1(branch_addr_i[24]), .A2(n103), .ZN(n152) );
  AOI22_X1 U175 ( .A1(n314), .A2(hwlp_addr_i[24]), .B1(n166), .B2(n9), .ZN(
        n151) );
  NAND2_X1 U176 ( .A1(prefetch_addr_i[24]), .A2(n307), .ZN(n150) );
  NAND3_X1 U177 ( .A1(n152), .A2(n151), .A3(n150), .ZN(instr_addr_o[24]) );
  NAND2_X1 U178 ( .A1(prefetch_addr_i[9]), .A2(n162), .ZN(n155) );
  NAND2_X1 U180 ( .A1(branch_addr_i[26]), .A2(n153), .ZN(n158) );
  AOI22_X1 U181 ( .A1(n308), .A2(hwlp_addr_i[26]), .B1(n166), .B2(n7), .ZN(
        n157) );
  NAND2_X1 U182 ( .A1(prefetch_addr_i[26]), .A2(n307), .ZN(n156) );
  NAND2_X1 U183 ( .A1(prefetch_addr_i[25]), .A2(n307), .ZN(n161) );
  AOI22_X1 U184 ( .A1(n314), .A2(hwlp_addr_i[25]), .B1(n166), .B2(n8), .ZN(
        n160) );
  OR2_X1 U185 ( .A1(n338), .A2(CS[2]), .ZN(n189) );
  NOR2_X1 U186 ( .A1(n189), .A2(n336), .ZN(n196) );
  NAND2_X1 U188 ( .A1(prefetch_addr_i[13]), .A2(n162), .ZN(n165) );
  AOI22_X1 U189 ( .A1(n308), .A2(hwlp_addr_i[13]), .B1(n163), .B2(n20), .ZN(
        n164) );
  AOI22_X1 U190 ( .A1(n314), .A2(hwlp_addr_i[31]), .B1(n166), .B2(n2), .ZN(
        n167) );
  OR2_X1 U191 ( .A1(n31), .A2(hwlp_i), .ZN(n168) );
  NOR2_X1 U192 ( .A1(prefetch_i), .A2(n168), .ZN(n221) );
  NAND2_X1 U193 ( .A1(n221), .A2(n180), .ZN(busy_o) );
  INV_X1 U194 ( .A(n196), .ZN(n169) );
  NAND3_X1 U195 ( .A1(n336), .A2(n338), .A3(CS[2]), .ZN(n299) );
  OAI21_X1 U196 ( .B1(n31), .B2(n169), .A(n299), .ZN(n170) );
  NAND2_X1 U197 ( .A1(n170), .A2(n188), .ZN(n198) );
  NAND2_X1 U198 ( .A1(busy_o), .A2(n198), .ZN(n193) );
  NAND2_X1 U199 ( .A1(CS[0]), .A2(CS[1]), .ZN(n171) );
  NAND2_X1 U200 ( .A1(n337), .A2(n171), .ZN(n172) );
  NOR2_X1 U201 ( .A1(n193), .A2(n172), .ZN(n192) );
  NAND2_X1 U202 ( .A1(n34), .A2(n337), .ZN(n177) );
  OAI21_X1 U203 ( .B1(n367), .B2(n177), .A(n299), .ZN(n173) );
  INV_X1 U204 ( .A(n173), .ZN(n174) );
  OAI22_X1 U205 ( .A1(n193), .A2(n174), .B1(n336), .B2(n198), .ZN(n175) );
  OR2_X1 U206 ( .A1(n192), .A2(n175), .ZN(n289) );
  NAND2_X1 U207 ( .A1(n177), .A2(n176), .ZN(n181) );
  INV_X1 U209 ( .A(n178), .ZN(n179) );
  AOI22_X1 U210 ( .A1(hwlp_i), .A2(n180), .B1(n179), .B2(n337), .ZN(n186) );
  NAND2_X1 U211 ( .A1(n31), .A2(n181), .ZN(n185) );
  INV_X1 U212 ( .A(n299), .ZN(n183) );
  OAI21_X1 U213 ( .B1(n183), .B2(n182), .A(n34), .ZN(n184) );
  OAI22_X1 U215 ( .A1(n193), .A2(n190), .B1(n189), .B2(n188), .ZN(n191) );
  OAI21_X1 U216 ( .B1(n192), .B2(n191), .A(instr_gnt_i), .ZN(n195) );
  AOI22_X1 U217 ( .A1(n193), .A2(CS[0]), .B1(n367), .B2(fetch_valid_o), .ZN(
        n194) );
  NAND2_X1 U218 ( .A1(n195), .A2(n194), .ZN(n288) );
  NAND3_X1 U219 ( .A1(n31), .A2(n196), .A3(n188), .ZN(n197) );
  OAI21_X1 U220 ( .B1(n198), .B2(n337), .A(n197), .ZN(n290) );
  INV_X1 U221 ( .A(instr_addr_o[4]), .ZN(n200) );
  NAND2_X1 U222 ( .A1(n367), .A2(n29), .ZN(n199) );
  OAI21_X1 U223 ( .B1(n367), .B2(n200), .A(n199), .ZN(n284) );
  INV_X1 U224 ( .A(n201), .ZN(n203) );
  NAND2_X1 U225 ( .A1(n367), .A2(n28), .ZN(n202) );
  OAI21_X1 U226 ( .B1(n367), .B2(n203), .A(n202), .ZN(n283) );
  INV_X1 U230 ( .A(instr_addr_o[7]), .ZN(n208) );
  NAND2_X1 U231 ( .A1(n367), .A2(n26), .ZN(n207) );
  OAI21_X1 U232 ( .B1(n367), .B2(n208), .A(n207), .ZN(n281) );
  NAND2_X1 U233 ( .A1(n367), .A2(n25), .ZN(n209) );
  OAI21_X1 U234 ( .B1(n367), .B2(n210), .A(n209), .ZN(n280) );
  NAND2_X1 U235 ( .A1(n367), .A2(n24), .ZN(n211) );
  OAI21_X1 U236 ( .B1(n367), .B2(n60), .A(n211), .ZN(n279) );
  NAND2_X1 U240 ( .A1(n367), .A2(n22), .ZN(n215) );
  OAI21_X1 U241 ( .B1(n367), .B2(n216), .A(n215), .ZN(n277) );
  INV_X1 U242 ( .A(n377), .ZN(n218) );
  NAND2_X1 U243 ( .A1(n367), .A2(n21), .ZN(n217) );
  OAI21_X1 U244 ( .B1(n367), .B2(n218), .A(n217), .ZN(n276) );
  INV_X1 U245 ( .A(instr_addr_o[13]), .ZN(n220) );
  NAND2_X1 U246 ( .A1(n367), .A2(n20), .ZN(n219) );
  OAI21_X1 U247 ( .B1(n367), .B2(n220), .A(n219), .ZN(n275) );
  NAND2_X1 U248 ( .A1(n367), .A2(n19), .ZN(n222) );
  OAI21_X1 U249 ( .B1(n367), .B2(n223), .A(n222), .ZN(n274) );
  INV_X1 U253 ( .A(n56), .ZN(n229) );
  NAND2_X1 U254 ( .A1(n367), .A2(n17), .ZN(n228) );
  OAI21_X1 U255 ( .B1(n221), .B2(n229), .A(n228), .ZN(n272) );
  INV_X1 U256 ( .A(n230), .ZN(n232) );
  NAND2_X1 U257 ( .A1(n367), .A2(n16), .ZN(n231) );
  OAI21_X1 U258 ( .B1(n367), .B2(n232), .A(n231), .ZN(n271) );
  INV_X1 U259 ( .A(n233), .ZN(n235) );
  NAND2_X1 U260 ( .A1(n367), .A2(n15), .ZN(n234) );
  OAI21_X1 U261 ( .B1(n367), .B2(n235), .A(n234), .ZN(n270) );
  INV_X1 U262 ( .A(n236), .ZN(n238) );
  NAND2_X1 U263 ( .A1(n367), .A2(n14), .ZN(n237) );
  OAI21_X1 U264 ( .B1(n221), .B2(n238), .A(n237), .ZN(n269) );
  NAND2_X1 U265 ( .A1(n367), .A2(n13), .ZN(n239) );
  OAI21_X1 U266 ( .B1(n367), .B2(n240), .A(n239), .ZN(n268) );
  INV_X1 U267 ( .A(instr_addr_o[21]), .ZN(n242) );
  NAND2_X1 U268 ( .A1(n367), .A2(n12), .ZN(n241) );
  OAI21_X1 U269 ( .B1(n367), .B2(n242), .A(n241), .ZN(n267) );
  INV_X1 U270 ( .A(n376), .ZN(n244) );
  NAND2_X1 U271 ( .A1(n367), .A2(n11), .ZN(n243) );
  OAI21_X1 U272 ( .B1(n367), .B2(n244), .A(n243), .ZN(n266) );
  INV_X1 U273 ( .A(instr_addr_o[23]), .ZN(n246) );
  NAND2_X1 U274 ( .A1(n367), .A2(n10), .ZN(n245) );
  OAI21_X1 U275 ( .B1(n367), .B2(n246), .A(n245), .ZN(n265) );
  INV_X1 U276 ( .A(instr_addr_o[24]), .ZN(n248) );
  NAND2_X1 U277 ( .A1(n367), .A2(n9), .ZN(n247) );
  OAI21_X1 U278 ( .B1(n367), .B2(n248), .A(n247), .ZN(n264) );
  INV_X1 U279 ( .A(instr_addr_o[25]), .ZN(n250) );
  NAND2_X1 U280 ( .A1(n367), .A2(n8), .ZN(n249) );
  OAI21_X1 U281 ( .B1(n367), .B2(n250), .A(n249), .ZN(n263) );
  INV_X1 U282 ( .A(n55), .ZN(n252) );
  NAND2_X1 U283 ( .A1(n367), .A2(n7), .ZN(n251) );
  OAI21_X1 U284 ( .B1(n367), .B2(n252), .A(n251), .ZN(n262) );
  INV_X1 U285 ( .A(instr_addr_o[27]), .ZN(n254) );
  NAND2_X1 U286 ( .A1(n367), .A2(n6), .ZN(n253) );
  OAI21_X1 U287 ( .B1(n367), .B2(n254), .A(n253), .ZN(n261) );
  NAND2_X1 U288 ( .A1(n367), .A2(n5), .ZN(n256) );
  OAI21_X1 U289 ( .B1(n367), .B2(n291), .A(n256), .ZN(n260) );
  INV_X1 U290 ( .A(instr_addr_o[29]), .ZN(n293) );
  NAND2_X1 U291 ( .A1(n367), .A2(n4), .ZN(n292) );
  OAI21_X1 U292 ( .B1(n367), .B2(n293), .A(n292), .ZN(n259) );
  NAND2_X1 U293 ( .A1(n367), .A2(n3), .ZN(n294) );
  OAI21_X1 U294 ( .B1(n367), .B2(n54), .A(n294), .ZN(n258) );
  INV_X1 U295 ( .A(instr_addr_o[31]), .ZN(n297) );
  NAND2_X1 U297 ( .A1(n367), .A2(n2), .ZN(n296) );
  OAI21_X1 U298 ( .B1(n367), .B2(n297), .A(n296), .ZN(n257) );
  NAND2_X1 U299 ( .A1(n31), .A2(n337), .ZN(n300) );
  NAND2_X1 U300 ( .A1(n300), .A2(n299), .ZN(n315) );
  NAND2_X1 U301 ( .A1(prefetch_addr_i[1]), .A2(n307), .ZN(n302) );
  NAND2_X1 U302 ( .A1(n314), .A2(hwlp_addr_i[1]), .ZN(n301) );
  NAND2_X1 U303 ( .A1(n302), .A2(n301), .ZN(n303) );
  AOI21_X1 U304 ( .B1(branch_addr_i[1]), .B2(n315), .A(n303), .ZN(n306) );
  NAND2_X1 U308 ( .A1(prefetch_addr_i[2]), .A2(n307), .ZN(n310) );
  NAND2_X1 U309 ( .A1(n308), .A2(hwlp_addr_i[2]), .ZN(n309) );
  NAND2_X1 U310 ( .A1(n310), .A2(n309), .ZN(n311) );
  AOI21_X1 U311 ( .B1(branch_addr_i[2]), .B2(n315), .A(n311), .ZN(n313) );
  AOI22_X1 U314 ( .A1(prefetch_addr_i[3]), .A2(n307), .B1(n314), .B2(
        hwlp_addr_i[3]), .ZN(n317) );
  NAND2_X1 U315 ( .A1(branch_addr_i[3]), .A2(n315), .ZN(n316) );
  NAND2_X1 U319 ( .A1(n34), .A2(instr_rdata_i[0]), .ZN(n321) );
  OAI21_X1 U320 ( .B1(n34), .B2(n339), .A(n321), .ZN(rdata_o[0]) );
  NAND2_X1 U321 ( .A1(n34), .A2(instr_rdata_i[1]), .ZN(n322) );
  OAI21_X1 U322 ( .B1(n371), .B2(n340), .A(n322), .ZN(rdata_o[1]) );
  NAND2_X1 U323 ( .A1(n34), .A2(instr_rdata_i[16]), .ZN(n323) );
  OAI21_X1 U324 ( .B1(n371), .B2(n341), .A(n323), .ZN(rdata_o[16]) );
  NAND2_X1 U325 ( .A1(n371), .A2(instr_rdata_i[17]), .ZN(n324) );
  OAI21_X1 U326 ( .B1(n371), .B2(n342), .A(n324), .ZN(rdata_o[17]) );
  NAND2_X1 U327 ( .A1(n34), .A2(instr_rdata_i[32]), .ZN(n325) );
  OAI21_X1 U328 ( .B1(n371), .B2(n343), .A(n325), .ZN(rdata_o[32]) );
  NAND2_X1 U329 ( .A1(n34), .A2(instr_rdata_i[33]), .ZN(n326) );
  OAI21_X1 U330 ( .B1(n371), .B2(n344), .A(n326), .ZN(rdata_o[33]) );
  MUX2_X1 U331 ( .A(L0_buffer[42]), .B(instr_rdata_i[48]), .S(n371), .Z(
        rdata_o[48]) );
  NAND2_X1 U332 ( .A1(n34), .A2(instr_rdata_i[49]), .ZN(n327) );
  OAI21_X1 U333 ( .B1(n34), .B2(n345), .A(n327), .ZN(rdata_o[49]) );
  NAND2_X1 U334 ( .A1(n34), .A2(instr_rdata_i[64]), .ZN(n328) );
  OAI21_X1 U335 ( .B1(n34), .B2(n346), .A(n328), .ZN(rdata_o[64]) );
  NAND2_X1 U336 ( .A1(n34), .A2(instr_rdata_i[65]), .ZN(n329) );
  OAI21_X1 U337 ( .B1(n34), .B2(n347), .A(n329), .ZN(rdata_o[65]) );
  NAND2_X1 U338 ( .A1(instr_rvalid_i), .A2(instr_rdata_i[80]), .ZN(n330) );
  OAI21_X1 U339 ( .B1(instr_rvalid_i), .B2(n348), .A(n330), .ZN(rdata_o[80])
         );
  NAND2_X1 U340 ( .A1(instr_rvalid_i), .A2(instr_rdata_i[81]), .ZN(n331) );
  OAI21_X1 U341 ( .B1(instr_rvalid_i), .B2(n349), .A(n331), .ZN(rdata_o[81])
         );
  NAND2_X1 U342 ( .A1(instr_rvalid_i), .A2(instr_rdata_i[96]), .ZN(n332) );
  OAI21_X1 U343 ( .B1(instr_rvalid_i), .B2(n350), .A(n332), .ZN(rdata_o[96])
         );
  NAND2_X1 U344 ( .A1(instr_rvalid_i), .A2(instr_rdata_i[97]), .ZN(n333) );
  MUX2_X1 U345 ( .A(L0_buffer[112]), .B(instr_rdata_i[127]), .S(n34), .Z(
        rdata_o[127]) );
  MUX2_X1 U346 ( .A(L0_buffer[111]), .B(instr_rdata_i[126]), .S(n371), .Z(
        rdata_o[126]) );
  MUX2_X1 U347 ( .A(L0_buffer[110]), .B(instr_rdata_i[125]), .S(n34), .Z(
        rdata_o[125]) );
  MUX2_X1 U348 ( .A(L0_buffer[109]), .B(instr_rdata_i[124]), .S(n34), .Z(
        rdata_o[124]) );
  MUX2_X1 U349 ( .A(L0_buffer[108]), .B(instr_rdata_i[123]), .S(n371), .Z(
        rdata_o[123]) );
  MUX2_X1 U350 ( .A(L0_buffer[107]), .B(instr_rdata_i[122]), .S(n34), .Z(
        rdata_o[122]) );
  MUX2_X1 U351 ( .A(L0_buffer[106]), .B(instr_rdata_i[121]), .S(n34), .Z(
        rdata_o[121]) );
  MUX2_X1 U352 ( .A(L0_buffer[105]), .B(instr_rdata_i[120]), .S(n34), .Z(
        rdata_o[120]) );
  MUX2_X1 U353 ( .A(L0_buffer[104]), .B(instr_rdata_i[119]), .S(n34), .Z(
        rdata_o[119]) );
  MUX2_X1 U354 ( .A(L0_buffer[103]), .B(instr_rdata_i[118]), .S(n34), .Z(
        rdata_o[118]) );
  MUX2_X1 U355 ( .A(L0_buffer[102]), .B(instr_rdata_i[117]), .S(n34), .Z(
        rdata_o[117]) );
  MUX2_X1 U356 ( .A(L0_buffer[101]), .B(instr_rdata_i[116]), .S(n34), .Z(
        rdata_o[116]) );
  MUX2_X1 U357 ( .A(L0_buffer[100]), .B(instr_rdata_i[115]), .S(n371), .Z(
        rdata_o[115]) );
  MUX2_X1 U358 ( .A(L0_buffer[99]), .B(instr_rdata_i[114]), .S(n34), .Z(
        rdata_o[114]) );
  MUX2_X1 U359 ( .A(L0_buffer[98]), .B(instr_rdata_i[111]), .S(n34), .Z(
        rdata_o[111]) );
  MUX2_X1 U360 ( .A(L0_buffer[97]), .B(instr_rdata_i[110]), .S(n34), .Z(
        rdata_o[110]) );
  MUX2_X1 U361 ( .A(L0_buffer[96]), .B(instr_rdata_i[109]), .S(n34), .Z(
        rdata_o[109]) );
  MUX2_X1 U362 ( .A(L0_buffer[95]), .B(instr_rdata_i[108]), .S(n34), .Z(
        rdata_o[108]) );
  MUX2_X1 U363 ( .A(L0_buffer[94]), .B(instr_rdata_i[107]), .S(n34), .Z(
        rdata_o[107]) );
  MUX2_X1 U364 ( .A(L0_buffer[93]), .B(instr_rdata_i[106]), .S(n34), .Z(
        rdata_o[106]) );
  MUX2_X1 U365 ( .A(L0_buffer[92]), .B(instr_rdata_i[105]), .S(n34), .Z(
        rdata_o[105]) );
  MUX2_X1 U366 ( .A(L0_buffer[91]), .B(instr_rdata_i[104]), .S(n34), .Z(
        rdata_o[104]) );
  MUX2_X1 U367 ( .A(L0_buffer[90]), .B(instr_rdata_i[103]), .S(n34), .Z(
        rdata_o[103]) );
  MUX2_X1 U368 ( .A(L0_buffer[89]), .B(instr_rdata_i[102]), .S(n371), .Z(
        rdata_o[102]) );
  MUX2_X1 U369 ( .A(L0_buffer[88]), .B(instr_rdata_i[101]), .S(n34), .Z(
        rdata_o[101]) );
  MUX2_X1 U370 ( .A(L0_buffer[87]), .B(instr_rdata_i[100]), .S(n34), .Z(
        rdata_o[100]) );
  MUX2_X1 U371 ( .A(L0_buffer[86]), .B(instr_rdata_i[99]), .S(n34), .Z(
        rdata_o[99]) );
  MUX2_X1 U372 ( .A(L0_buffer[85]), .B(instr_rdata_i[98]), .S(n34), .Z(
        rdata_o[98]) );
  MUX2_X1 U373 ( .A(L0_buffer[84]), .B(instr_rdata_i[95]), .S(n34), .Z(
        rdata_o[95]) );
  MUX2_X1 U374 ( .A(L0_buffer[83]), .B(instr_rdata_i[94]), .S(n34), .Z(
        rdata_o[94]) );
  MUX2_X1 U375 ( .A(L0_buffer[82]), .B(instr_rdata_i[93]), .S(n371), .Z(
        rdata_o[93]) );
  MUX2_X1 U376 ( .A(L0_buffer[81]), .B(instr_rdata_i[92]), .S(n34), .Z(
        rdata_o[92]) );
  MUX2_X1 U377 ( .A(L0_buffer[80]), .B(instr_rdata_i[91]), .S(n34), .Z(
        rdata_o[91]) );
  MUX2_X1 U378 ( .A(L0_buffer[79]), .B(instr_rdata_i[90]), .S(n371), .Z(
        rdata_o[90]) );
  MUX2_X1 U379 ( .A(L0_buffer[78]), .B(instr_rdata_i[89]), .S(n34), .Z(
        rdata_o[89]) );
  MUX2_X1 U380 ( .A(L0_buffer[77]), .B(instr_rdata_i[88]), .S(n34), .Z(
        rdata_o[88]) );
  MUX2_X1 U381 ( .A(L0_buffer[76]), .B(instr_rdata_i[87]), .S(n371), .Z(
        rdata_o[87]) );
  MUX2_X1 U382 ( .A(L0_buffer[75]), .B(instr_rdata_i[86]), .S(n34), .Z(
        rdata_o[86]) );
  MUX2_X1 U383 ( .A(L0_buffer[74]), .B(instr_rdata_i[85]), .S(n34), .Z(
        rdata_o[85]) );
  MUX2_X1 U384 ( .A(L0_buffer[73]), .B(instr_rdata_i[84]), .S(n34), .Z(
        rdata_o[84]) );
  MUX2_X1 U385 ( .A(L0_buffer[72]), .B(instr_rdata_i[83]), .S(n34), .Z(
        rdata_o[83]) );
  MUX2_X1 U386 ( .A(L0_buffer[71]), .B(instr_rdata_i[82]), .S(n34), .Z(
        rdata_o[82]) );
  MUX2_X1 U387 ( .A(L0_buffer[70]), .B(instr_rdata_i[79]), .S(n34), .Z(
        rdata_o[79]) );
  MUX2_X1 U388 ( .A(L0_buffer[69]), .B(instr_rdata_i[78]), .S(n34), .Z(
        rdata_o[78]) );
  MUX2_X1 U389 ( .A(L0_buffer[68]), .B(instr_rdata_i[77]), .S(n34), .Z(
        rdata_o[77]) );
  MUX2_X1 U390 ( .A(L0_buffer[67]), .B(instr_rdata_i[76]), .S(n34), .Z(
        rdata_o[76]) );
  MUX2_X1 U391 ( .A(L0_buffer[66]), .B(instr_rdata_i[75]), .S(n34), .Z(
        rdata_o[75]) );
  MUX2_X1 U392 ( .A(L0_buffer[65]), .B(instr_rdata_i[74]), .S(n34), .Z(
        rdata_o[74]) );
  MUX2_X1 U393 ( .A(L0_buffer[64]), .B(instr_rdata_i[73]), .S(n34), .Z(
        rdata_o[73]) );
  MUX2_X1 U394 ( .A(L0_buffer[63]), .B(instr_rdata_i[72]), .S(n34), .Z(
        rdata_o[72]) );
  MUX2_X1 U395 ( .A(L0_buffer[62]), .B(instr_rdata_i[71]), .S(n34), .Z(
        rdata_o[71]) );
  MUX2_X1 U396 ( .A(L0_buffer[61]), .B(instr_rdata_i[70]), .S(n34), .Z(
        rdata_o[70]) );
  MUX2_X1 U397 ( .A(L0_buffer[60]), .B(instr_rdata_i[69]), .S(n34), .Z(
        rdata_o[69]) );
  MUX2_X1 U398 ( .A(L0_buffer[59]), .B(instr_rdata_i[68]), .S(n34), .Z(
        rdata_o[68]) );
  MUX2_X1 U399 ( .A(L0_buffer[58]), .B(instr_rdata_i[67]), .S(n34), .Z(
        rdata_o[67]) );
  MUX2_X1 U400 ( .A(L0_buffer[57]), .B(instr_rdata_i[66]), .S(n34), .Z(
        rdata_o[66]) );
  MUX2_X1 U401 ( .A(L0_buffer[56]), .B(instr_rdata_i[63]), .S(n34), .Z(
        rdata_o[63]) );
  MUX2_X1 U402 ( .A(L0_buffer[55]), .B(instr_rdata_i[62]), .S(n34), .Z(
        rdata_o[62]) );
  MUX2_X1 U403 ( .A(L0_buffer[54]), .B(instr_rdata_i[61]), .S(n34), .Z(
        rdata_o[61]) );
  MUX2_X1 U404 ( .A(L0_buffer[53]), .B(instr_rdata_i[60]), .S(n34), .Z(
        rdata_o[60]) );
  MUX2_X1 U405 ( .A(L0_buffer[52]), .B(instr_rdata_i[59]), .S(n34), .Z(
        rdata_o[59]) );
  MUX2_X1 U406 ( .A(L0_buffer[51]), .B(instr_rdata_i[58]), .S(n34), .Z(
        rdata_o[58]) );
  MUX2_X1 U407 ( .A(L0_buffer[50]), .B(instr_rdata_i[57]), .S(n34), .Z(
        rdata_o[57]) );
  MUX2_X1 U408 ( .A(L0_buffer[49]), .B(instr_rdata_i[56]), .S(n34), .Z(
        rdata_o[56]) );
  MUX2_X1 U410 ( .A(L0_buffer[48]), .B(instr_rdata_i[55]), .S(n34), .Z(
        rdata_o[55]) );
  MUX2_X1 U411 ( .A(L0_buffer[47]), .B(instr_rdata_i[54]), .S(n34), .Z(
        rdata_o[54]) );
  MUX2_X1 U412 ( .A(L0_buffer[46]), .B(instr_rdata_i[53]), .S(n34), .Z(
        rdata_o[53]) );
  MUX2_X1 U413 ( .A(L0_buffer[45]), .B(instr_rdata_i[52]), .S(n34), .Z(
        rdata_o[52]) );
  MUX2_X1 U414 ( .A(L0_buffer[44]), .B(instr_rdata_i[51]), .S(n34), .Z(
        rdata_o[51]) );
  MUX2_X1 U415 ( .A(L0_buffer[43]), .B(instr_rdata_i[50]), .S(n34), .Z(
        rdata_o[50]) );
  MUX2_X1 U416 ( .A(L0_buffer[41]), .B(instr_rdata_i[47]), .S(n34), .Z(
        rdata_o[47]) );
  MUX2_X1 U417 ( .A(L0_buffer[40]), .B(instr_rdata_i[46]), .S(n34), .Z(
        rdata_o[46]) );
  MUX2_X1 U418 ( .A(L0_buffer[39]), .B(instr_rdata_i[45]), .S(n34), .Z(
        rdata_o[45]) );
  MUX2_X1 U419 ( .A(L0_buffer[38]), .B(instr_rdata_i[44]), .S(n34), .Z(
        rdata_o[44]) );
  MUX2_X1 U420 ( .A(L0_buffer[37]), .B(instr_rdata_i[43]), .S(n34), .Z(
        rdata_o[43]) );
  MUX2_X1 U421 ( .A(L0_buffer[36]), .B(instr_rdata_i[42]), .S(n34), .Z(
        rdata_o[42]) );
  MUX2_X1 U422 ( .A(L0_buffer[35]), .B(instr_rdata_i[41]), .S(n34), .Z(
        rdata_o[41]) );
  MUX2_X1 U423 ( .A(L0_buffer[34]), .B(instr_rdata_i[40]), .S(n34), .Z(
        rdata_o[40]) );
  MUX2_X1 U424 ( .A(L0_buffer[33]), .B(instr_rdata_i[39]), .S(n34), .Z(
        rdata_o[39]) );
  MUX2_X1 U425 ( .A(L0_buffer[32]), .B(instr_rdata_i[38]), .S(n34), .Z(
        rdata_o[38]) );
  MUX2_X1 U426 ( .A(L0_buffer[31]), .B(instr_rdata_i[37]), .S(n34), .Z(
        rdata_o[37]) );
  MUX2_X1 U427 ( .A(L0_buffer[30]), .B(instr_rdata_i[36]), .S(n34), .Z(
        rdata_o[36]) );
  MUX2_X1 U428 ( .A(L0_buffer[29]), .B(instr_rdata_i[35]), .S(n371), .Z(
        rdata_o[35]) );
  MUX2_X1 U429 ( .A(L0_buffer[28]), .B(instr_rdata_i[34]), .S(n371), .Z(
        rdata_o[34]) );
  MUX2_X1 U430 ( .A(L0_buffer[27]), .B(instr_rdata_i[31]), .S(n371), .Z(
        rdata_o[31]) );
  MUX2_X1 U431 ( .A(L0_buffer[26]), .B(instr_rdata_i[30]), .S(n371), .Z(
        rdata_o[30]) );
  MUX2_X1 U432 ( .A(L0_buffer[25]), .B(instr_rdata_i[29]), .S(n34), .Z(
        rdata_o[29]) );
  MUX2_X1 U433 ( .A(L0_buffer[24]), .B(instr_rdata_i[28]), .S(n371), .Z(
        rdata_o[28]) );
  MUX2_X1 U434 ( .A(L0_buffer[23]), .B(instr_rdata_i[27]), .S(n34), .Z(
        rdata_o[27]) );
  MUX2_X1 U435 ( .A(L0_buffer[22]), .B(instr_rdata_i[26]), .S(n371), .Z(
        rdata_o[26]) );
  MUX2_X1 U436 ( .A(L0_buffer[21]), .B(instr_rdata_i[25]), .S(n371), .Z(
        rdata_o[25]) );
  MUX2_X1 U437 ( .A(L0_buffer[20]), .B(instr_rdata_i[24]), .S(n371), .Z(
        rdata_o[24]) );
  MUX2_X1 U438 ( .A(L0_buffer[19]), .B(instr_rdata_i[23]), .S(n34), .Z(
        rdata_o[23]) );
  MUX2_X1 U439 ( .A(L0_buffer[18]), .B(instr_rdata_i[22]), .S(n371), .Z(
        rdata_o[22]) );
  MUX2_X1 U440 ( .A(L0_buffer[17]), .B(instr_rdata_i[21]), .S(n34), .Z(
        rdata_o[21]) );
  MUX2_X1 U441 ( .A(L0_buffer[16]), .B(instr_rdata_i[20]), .S(n34), .Z(
        rdata_o[20]) );
  MUX2_X1 U442 ( .A(L0_buffer[15]), .B(instr_rdata_i[19]), .S(n371), .Z(
        rdata_o[19]) );
  MUX2_X1 U443 ( .A(L0_buffer[14]), .B(instr_rdata_i[18]), .S(n34), .Z(
        rdata_o[18]) );
  MUX2_X1 U444 ( .A(L0_buffer[13]), .B(instr_rdata_i[15]), .S(n34), .Z(
        rdata_o[15]) );
  MUX2_X1 U445 ( .A(L0_buffer[12]), .B(instr_rdata_i[14]), .S(n34), .Z(
        rdata_o[14]) );
  MUX2_X1 U446 ( .A(L0_buffer[11]), .B(instr_rdata_i[13]), .S(n34), .Z(
        rdata_o[13]) );
  MUX2_X1 U447 ( .A(L0_buffer[10]), .B(instr_rdata_i[12]), .S(n34), .Z(
        rdata_o[12]) );
  MUX2_X1 U448 ( .A(L0_buffer[9]), .B(instr_rdata_i[11]), .S(n34), .Z(
        rdata_o[11]) );
  MUX2_X1 U449 ( .A(L0_buffer[8]), .B(instr_rdata_i[10]), .S(n371), .Z(
        rdata_o[10]) );
  MUX2_X1 U450 ( .A(L0_buffer[7]), .B(instr_rdata_i[9]), .S(n371), .Z(
        rdata_o[9]) );
  MUX2_X1 U451 ( .A(L0_buffer[6]), .B(instr_rdata_i[8]), .S(n34), .Z(
        rdata_o[8]) );
  MUX2_X1 U452 ( .A(L0_buffer[5]), .B(instr_rdata_i[7]), .S(n371), .Z(
        rdata_o[7]) );
  MUX2_X1 U453 ( .A(L0_buffer[4]), .B(instr_rdata_i[6]), .S(n371), .Z(
        rdata_o[6]) );
  MUX2_X1 U454 ( .A(L0_buffer[3]), .B(instr_rdata_i[5]), .S(n34), .Z(
        rdata_o[5]) );
  MUX2_X1 U455 ( .A(L0_buffer[2]), .B(instr_rdata_i[4]), .S(n34), .Z(
        rdata_o[4]) );
  MUX2_X1 U456 ( .A(L0_buffer[1]), .B(instr_rdata_i[3]), .S(n34), .Z(
        rdata_o[3]) );
  MUX2_X1 U457 ( .A(L0_buffer[0]), .B(instr_rdata_i[2]), .S(n34), .Z(
        rdata_o[2]) );
  SDFFR_X1 CS_reg_2_ ( .D(n290), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(rst_n), 
        .Q(CS[2]), .QN(n337) );
  SDFFR_X1 addr_q_reg_3_ ( .D(n387), .SI(1'b0), .SE(1'b0), .CK(n714), .RN(
        rst_n), .Q(addr_o[3]) );
  SDFFR_X1 addr_q_reg_1_ ( .D(n712), .SI(1'b0), .SE(1'b0), .CK(n714), .RN(
        rst_n), .Q(addr_o[1]) );
  SDFFR_X1 addr_q_reg_2_ ( .D(n713), .SI(1'b0), .SE(1'b0), .CK(n714), .RN(
        rst_n), .Q(addr_o[2]) );
  SDFFR_X1 addr_q_reg_4_ ( .D(n284), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n29) );
  SDFFR_X1 addr_q_reg_5_ ( .D(n283), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n28) );
  SDFFR_X1 addr_q_reg_6_ ( .D(instr_addr_o[6]), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(rst_n), .Q(n27) );
  SDFFR_X1 addr_q_reg_7_ ( .D(n281), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n26) );
  SDFFR_X1 addr_q_reg_8_ ( .D(n280), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n25) );
  SDFFR_X1 addr_q_reg_9_ ( .D(n279), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n24) );
  SDFFR_X1 addr_q_reg_10_ ( .D(n212), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n23) );
  SDFFR_X1 addr_q_reg_11_ ( .D(n277), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n22) );
  SDFFR_X1 addr_q_reg_12_ ( .D(n276), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n21) );
  SDFFR_X1 addr_q_reg_13_ ( .D(n275), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n20) );
  SDFFR_X1 addr_q_reg_14_ ( .D(n274), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n19) );
  SDFFR_X1 addr_q_reg_15_ ( .D(n224), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n18) );
  SDFFR_X1 addr_q_reg_16_ ( .D(n272), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n17) );
  SDFFR_X1 addr_q_reg_17_ ( .D(n271), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n16) );
  SDFFR_X1 addr_q_reg_18_ ( .D(n270), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n15) );
  SDFFR_X1 addr_q_reg_19_ ( .D(n269), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n14) );
  SDFFR_X1 addr_q_reg_20_ ( .D(n268), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n13) );
  SDFFR_X1 addr_q_reg_21_ ( .D(n267), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n12) );
  SDFFR_X1 addr_q_reg_22_ ( .D(n266), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n11) );
  SDFFR_X1 addr_q_reg_23_ ( .D(n265), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n10) );
  SDFFR_X1 addr_q_reg_24_ ( .D(n264), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n9) );
  SDFFR_X1 addr_q_reg_25_ ( .D(n263), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n8) );
  SDFFR_X1 addr_q_reg_26_ ( .D(n262), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n7) );
  SDFFR_X1 addr_q_reg_27_ ( .D(n261), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n6) );
  SDFFR_X1 addr_q_reg_28_ ( .D(n260), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n5) );
  SDFFR_X1 addr_q_reg_29_ ( .D(n259), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n4) );
  SDFFR_X1 addr_q_reg_30_ ( .D(n258), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n3) );
  SDFFR_X1 addr_q_reg_31_ ( .D(n257), .SI(1'b0), .SE(1'b0), .CK(n709), .RN(
        rst_n), .Q(n2) );
  SDFFR_X1 L0_buffer_reg_3__31_ ( .D(instr_rdata_i[127]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[112]) );
  SDFFR_X1 L0_buffer_reg_3__30_ ( .D(instr_rdata_i[126]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[111]) );
  SDFFR_X1 L0_buffer_reg_3__29_ ( .D(instr_rdata_i[125]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[110]) );
  SDFFR_X1 L0_buffer_reg_3__28_ ( .D(instr_rdata_i[124]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[109]) );
  SDFFR_X1 L0_buffer_reg_3__27_ ( .D(instr_rdata_i[123]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[108]) );
  SDFFR_X1 L0_buffer_reg_3__26_ ( .D(instr_rdata_i[122]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[107]) );
  SDFFR_X1 L0_buffer_reg_3__25_ ( .D(instr_rdata_i[121]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[106]) );
  SDFFR_X1 L0_buffer_reg_3__24_ ( .D(instr_rdata_i[120]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[105]) );
  SDFFR_X1 L0_buffer_reg_3__23_ ( .D(instr_rdata_i[119]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[104]) );
  SDFFR_X1 L0_buffer_reg_3__22_ ( .D(instr_rdata_i[118]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[103]) );
  SDFFR_X1 L0_buffer_reg_3__21_ ( .D(instr_rdata_i[117]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[102]) );
  SDFFR_X1 L0_buffer_reg_3__20_ ( .D(instr_rdata_i[116]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[101]) );
  SDFFR_X1 L0_buffer_reg_3__19_ ( .D(instr_rdata_i[115]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[100]) );
  SDFFR_X1 L0_buffer_reg_3__18_ ( .D(instr_rdata_i[114]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[99]) );
  SDFFR_X1 L0_buffer_reg_3__17_ ( .D(instr_rdata_i[113]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .QN(n353) );
  SDFFR_X1 L0_buffer_reg_3__16_ ( .D(instr_rdata_i[112]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .QN(n352) );
  SDFFR_X1 L0_buffer_reg_3__15_ ( .D(instr_rdata_i[111]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[98]) );
  SDFFR_X1 L0_buffer_reg_3__14_ ( .D(instr_rdata_i[110]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[97]) );
  SDFFR_X1 L0_buffer_reg_3__13_ ( .D(instr_rdata_i[109]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[96]) );
  SDFFR_X1 L0_buffer_reg_3__12_ ( .D(instr_rdata_i[108]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[95]) );
  SDFFR_X1 L0_buffer_reg_3__11_ ( .D(instr_rdata_i[107]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[94]) );
  SDFFR_X1 L0_buffer_reg_3__10_ ( .D(instr_rdata_i[106]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[93]) );
  SDFFR_X1 L0_buffer_reg_3__9_ ( .D(instr_rdata_i[105]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[92]) );
  SDFFR_X1 L0_buffer_reg_3__8_ ( .D(instr_rdata_i[104]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[91]) );
  SDFFR_X1 L0_buffer_reg_3__7_ ( .D(instr_rdata_i[103]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[90]) );
  SDFFR_X1 L0_buffer_reg_3__6_ ( .D(instr_rdata_i[102]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[89]) );
  SDFFR_X1 L0_buffer_reg_3__5_ ( .D(instr_rdata_i[101]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[88]) );
  SDFFR_X1 L0_buffer_reg_3__4_ ( .D(instr_rdata_i[100]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[87]) );
  SDFFR_X1 L0_buffer_reg_3__3_ ( .D(instr_rdata_i[99]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[86]) );
  SDFFR_X1 L0_buffer_reg_3__2_ ( .D(instr_rdata_i[98]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[85]) );
  SDFFR_X1 L0_buffer_reg_3__1_ ( .D(instr_rdata_i[97]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .QN(n351) );
  SDFFR_X1 L0_buffer_reg_3__0_ ( .D(instr_rdata_i[96]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .QN(n350) );
  SDFFR_X1 L0_buffer_reg_2__31_ ( .D(instr_rdata_i[95]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[84]) );
  SDFFR_X1 L0_buffer_reg_2__30_ ( .D(instr_rdata_i[94]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[83]) );
  SDFFR_X1 L0_buffer_reg_2__29_ ( .D(instr_rdata_i[93]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[82]) );
  SDFFR_X1 L0_buffer_reg_2__28_ ( .D(instr_rdata_i[92]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[81]) );
  SDFFR_X1 L0_buffer_reg_2__27_ ( .D(instr_rdata_i[91]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[80]) );
  SDFFR_X1 L0_buffer_reg_2__26_ ( .D(instr_rdata_i[90]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[79]) );
  SDFFR_X1 L0_buffer_reg_2__25_ ( .D(instr_rdata_i[89]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[78]) );
  SDFFR_X1 L0_buffer_reg_2__24_ ( .D(instr_rdata_i[88]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[77]) );
  SDFFR_X1 L0_buffer_reg_2__23_ ( .D(instr_rdata_i[87]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[76]) );
  SDFFR_X1 L0_buffer_reg_2__22_ ( .D(instr_rdata_i[86]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[75]) );
  SDFFR_X1 L0_buffer_reg_2__21_ ( .D(instr_rdata_i[85]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[74]) );
  SDFFR_X1 L0_buffer_reg_2__20_ ( .D(instr_rdata_i[84]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[73]) );
  SDFFR_X1 L0_buffer_reg_2__19_ ( .D(instr_rdata_i[83]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[72]) );
  SDFFR_X1 L0_buffer_reg_2__18_ ( .D(instr_rdata_i[82]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[71]) );
  SDFFR_X1 L0_buffer_reg_2__17_ ( .D(instr_rdata_i[81]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .QN(n349) );
  SDFFR_X1 L0_buffer_reg_2__16_ ( .D(instr_rdata_i[80]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .QN(n348) );
  SDFFR_X1 L0_buffer_reg_2__15_ ( .D(instr_rdata_i[79]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[70]) );
  SDFFR_X1 L0_buffer_reg_2__14_ ( .D(instr_rdata_i[78]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[69]) );
  SDFFR_X1 L0_buffer_reg_2__13_ ( .D(instr_rdata_i[77]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[68]) );
  SDFFR_X1 L0_buffer_reg_2__12_ ( .D(instr_rdata_i[76]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[67]) );
  SDFFR_X1 L0_buffer_reg_2__11_ ( .D(instr_rdata_i[75]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[66]) );
  SDFFR_X1 L0_buffer_reg_2__10_ ( .D(instr_rdata_i[74]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[65]) );
  SDFFR_X1 L0_buffer_reg_2__9_ ( .D(instr_rdata_i[73]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[64]) );
  SDFFR_X1 L0_buffer_reg_2__8_ ( .D(instr_rdata_i[72]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[63]) );
  SDFFR_X1 L0_buffer_reg_2__7_ ( .D(instr_rdata_i[71]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[62]) );
  SDFFR_X1 L0_buffer_reg_2__6_ ( .D(instr_rdata_i[70]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[61]) );
  SDFFR_X1 L0_buffer_reg_2__5_ ( .D(instr_rdata_i[69]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[60]) );
  SDFFR_X1 L0_buffer_reg_2__4_ ( .D(instr_rdata_i[68]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[59]) );
  SDFFR_X1 L0_buffer_reg_2__3_ ( .D(instr_rdata_i[67]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[58]) );
  SDFFR_X1 L0_buffer_reg_2__2_ ( .D(instr_rdata_i[66]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[57]) );
  SDFFR_X1 L0_buffer_reg_2__1_ ( .D(n716), .SI(1'b0), .SE(1'b0), .CK(n720), 
        .RN(rst_n), .QN(n347) );
  SDFFR_X1 L0_buffer_reg_2__0_ ( .D(instr_rdata_i[64]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .QN(n346) );
  SDFFR_X1 L0_buffer_reg_1__31_ ( .D(instr_rdata_i[63]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[56]) );
  SDFFR_X1 L0_buffer_reg_1__30_ ( .D(instr_rdata_i[62]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[55]) );
  SDFFR_X1 L0_buffer_reg_1__29_ ( .D(instr_rdata_i[61]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[54]) );
  SDFFR_X1 L0_buffer_reg_1__28_ ( .D(instr_rdata_i[60]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[53]) );
  SDFFR_X1 L0_buffer_reg_1__27_ ( .D(instr_rdata_i[59]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[52]) );
  SDFFR_X1 L0_buffer_reg_1__26_ ( .D(instr_rdata_i[58]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[51]) );
  SDFFR_X1 L0_buffer_reg_1__25_ ( .D(instr_rdata_i[57]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[50]) );
  SDFFR_X1 L0_buffer_reg_1__24_ ( .D(instr_rdata_i[56]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[49]) );
  SDFFR_X1 L0_buffer_reg_1__23_ ( .D(instr_rdata_i[55]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[48]) );
  SDFFR_X1 L0_buffer_reg_1__22_ ( .D(instr_rdata_i[54]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[47]) );
  SDFFR_X1 L0_buffer_reg_1__21_ ( .D(instr_rdata_i[53]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[46]) );
  SDFFR_X1 L0_buffer_reg_1__20_ ( .D(instr_rdata_i[52]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[45]) );
  SDFFR_X1 L0_buffer_reg_1__19_ ( .D(instr_rdata_i[51]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[44]) );
  SDFFR_X1 L0_buffer_reg_1__18_ ( .D(instr_rdata_i[50]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[43]) );
  SDFFR_X1 L0_buffer_reg_1__17_ ( .D(instr_rdata_i[49]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .QN(n345) );
  SDFFR_X1 L0_buffer_reg_1__16_ ( .D(instr_rdata_i[48]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[42]) );
  SDFFR_X1 L0_buffer_reg_1__15_ ( .D(instr_rdata_i[47]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[41]) );
  SDFFR_X1 L0_buffer_reg_1__14_ ( .D(instr_rdata_i[46]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[40]) );
  SDFFR_X1 L0_buffer_reg_1__13_ ( .D(instr_rdata_i[45]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[39]) );
  SDFFR_X1 L0_buffer_reg_1__12_ ( .D(instr_rdata_i[44]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[38]) );
  SDFFR_X1 L0_buffer_reg_1__11_ ( .D(instr_rdata_i[43]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[37]) );
  SDFFR_X1 L0_buffer_reg_1__10_ ( .D(instr_rdata_i[42]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[36]) );
  SDFFR_X1 L0_buffer_reg_1__9_ ( .D(instr_rdata_i[41]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[35]) );
  SDFFR_X1 L0_buffer_reg_1__8_ ( .D(instr_rdata_i[40]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[34]) );
  SDFFR_X1 L0_buffer_reg_1__7_ ( .D(instr_rdata_i[39]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[33]) );
  SDFFR_X1 L0_buffer_reg_1__6_ ( .D(instr_rdata_i[38]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[32]) );
  SDFFR_X1 L0_buffer_reg_1__5_ ( .D(instr_rdata_i[37]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[31]) );
  SDFFR_X1 L0_buffer_reg_1__4_ ( .D(instr_rdata_i[36]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[30]) );
  SDFFR_X1 L0_buffer_reg_1__3_ ( .D(instr_rdata_i[35]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[29]) );
  SDFFR_X1 L0_buffer_reg_1__2_ ( .D(instr_rdata_i[34]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[28]) );
  SDFFR_X1 L0_buffer_reg_1__1_ ( .D(n717), .SI(1'b0), .SE(1'b0), .CK(n720), 
        .RN(rst_n), .QN(n344) );
  SDFFR_X1 L0_buffer_reg_1__0_ ( .D(instr_rdata_i[32]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .QN(n343) );
  SDFFR_X1 L0_buffer_reg_0__31_ ( .D(instr_rdata_i[31]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[27]) );
  SDFFR_X1 L0_buffer_reg_0__30_ ( .D(instr_rdata_i[30]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[26]) );
  SDFFR_X1 L0_buffer_reg_0__29_ ( .D(instr_rdata_i[29]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[25]) );
  SDFFR_X1 L0_buffer_reg_0__28_ ( .D(instr_rdata_i[28]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[24]) );
  SDFFR_X1 L0_buffer_reg_0__27_ ( .D(instr_rdata_i[27]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[23]) );
  SDFFR_X1 L0_buffer_reg_0__26_ ( .D(instr_rdata_i[26]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[22]) );
  SDFFR_X1 L0_buffer_reg_0__25_ ( .D(instr_rdata_i[25]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[21]) );
  SDFFR_X1 L0_buffer_reg_0__24_ ( .D(instr_rdata_i[24]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[20]) );
  SDFFR_X1 L0_buffer_reg_0__23_ ( .D(instr_rdata_i[23]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[19]) );
  SDFFR_X1 L0_buffer_reg_0__22_ ( .D(instr_rdata_i[22]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[18]) );
  SDFFR_X1 L0_buffer_reg_0__21_ ( .D(instr_rdata_i[21]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[17]) );
  SDFFR_X1 L0_buffer_reg_0__20_ ( .D(instr_rdata_i[20]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[16]) );
  SDFFR_X1 L0_buffer_reg_0__19_ ( .D(instr_rdata_i[19]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[15]) );
  SDFFR_X1 L0_buffer_reg_0__18_ ( .D(instr_rdata_i[18]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[14]) );
  SDFFR_X1 L0_buffer_reg_0__17_ ( .D(n718), .SI(1'b0), .SE(1'b0), .CK(n720), 
        .RN(rst_n), .QN(n342) );
  SDFFR_X1 L0_buffer_reg_0__16_ ( .D(n719), .SI(1'b0), .SE(1'b0), .CK(n720), 
        .RN(rst_n), .QN(n341) );
  SDFFR_X1 L0_buffer_reg_0__15_ ( .D(instr_rdata_i[15]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[13]) );
  SDFFR_X1 L0_buffer_reg_0__14_ ( .D(instr_rdata_i[14]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[12]) );
  SDFFR_X1 L0_buffer_reg_0__13_ ( .D(instr_rdata_i[13]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[11]) );
  SDFFR_X1 L0_buffer_reg_0__12_ ( .D(instr_rdata_i[12]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[10]) );
  SDFFR_X1 L0_buffer_reg_0__11_ ( .D(instr_rdata_i[11]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[9]) );
  SDFFR_X1 L0_buffer_reg_0__10_ ( .D(instr_rdata_i[10]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[8]) );
  SDFFR_X1 L0_buffer_reg_0__9_ ( .D(instr_rdata_i[9]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[7]) );
  SDFFR_X1 L0_buffer_reg_0__8_ ( .D(instr_rdata_i[8]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[6]) );
  SDFFR_X1 L0_buffer_reg_0__7_ ( .D(instr_rdata_i[7]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[5]) );
  SDFFR_X1 L0_buffer_reg_0__6_ ( .D(instr_rdata_i[6]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[4]) );
  SDFFR_X1 L0_buffer_reg_0__5_ ( .D(instr_rdata_i[5]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[3]) );
  SDFFR_X1 L0_buffer_reg_0__4_ ( .D(instr_rdata_i[4]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[2]) );
  SDFFR_X1 L0_buffer_reg_0__3_ ( .D(instr_rdata_i[3]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[1]) );
  SDFFR_X1 L0_buffer_reg_0__2_ ( .D(instr_rdata_i[2]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .Q(L0_buffer[0]) );
  SDFFR_X1 L0_buffer_reg_0__1_ ( .D(instr_rdata_i[1]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .QN(n340) );
  SDFFR_X1 L0_buffer_reg_0__0_ ( .D(instr_rdata_i[0]), .SI(1'b0), .SE(1'b0), 
        .CK(n720), .RN(rst_n), .QN(n339) );
  CLKBUF_X3 U26 ( .A(n304), .Z(n166) );
  CLKBUF_X3 U28 ( .A(n106), .Z(n307) );
  SNPS_CLOCK_GATE_HIGH_riscv_L0_buffer_RDATA_IN_WIDTH128_0 clk_gate_L0_buffer_reg_0__0_ ( 
        .CLK(clk), .EN(n34), .ENCLK(n720), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_L0_buffer_RDATA_IN_WIDTH128_1 clk_gate_addr_q_reg_2_ ( 
        .CLK(clk), .EN(n388), .ENCLK(n714), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_L0_buffer_RDATA_IN_WIDTH128_2 clk_gate_addr_q_reg_15_ ( 
        .CLK(clk), .EN(n711), .ENCLK(n709), .TE(1'b0) );
  SDFFR_X1 CS_reg_0_ ( .D(n288), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(rst_n), 
        .Q(CS[0]), .QN(n338) );
  SDFFR_X1 CS_reg_1_ ( .D(n289), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(rst_n), 
        .Q(CS[1]), .QN(n336) );
  AND2_X1 U187 ( .A1(n34), .A2(n196), .ZN(fetch_valid_o) );
  BUF_X1 U10 ( .A(n103), .Z(n159) );
  NAND3_X1 U14 ( .A1(n128), .A2(n126), .A3(n127), .ZN(instr_addr_o[4]) );
  BUF_X2 U4 ( .A(n103), .Z(n153) );
  INV_X4 U5 ( .A(n188), .ZN(n371) );
  CLKBUF_X3 U6 ( .A(n221), .Z(n367) );
  CLKBUF_X1 U7 ( .A(instr_addr_o[12]), .Z(n377) );
  BUF_X2 U8 ( .A(n87), .Z(n314) );
  BUF_X2 U9 ( .A(n304), .Z(n163) );
  OAI21_X1 U11 ( .B1(instr_rvalid_i), .B2(n352), .A(n77), .ZN(rdata_o[112]) );
  CLKBUF_X1 U12 ( .A(instr_addr_o[22]), .Z(n376) );
  CLKBUF_X1 U13 ( .A(instr_addr_o[14]), .Z(n375) );
  INV_X1 U15 ( .A(n34), .ZN(n188) );
  BUF_X8 U16 ( .A(instr_rvalid_i), .Z(n34) );
  NAND3_X1 U17 ( .A1(n69), .A2(n154), .A3(n155), .ZN(instr_addr_o[9]) );
  NAND2_X1 U18 ( .A1(branch_addr_i[9]), .A2(n153), .ZN(n69) );
  NAND3_X1 U19 ( .A1(n372), .A2(n142), .A3(n143), .ZN(instr_addr_o[19]) );
  NAND2_X1 U20 ( .A1(branch_addr_i[19]), .A2(n159), .ZN(n372) );
  NAND3_X1 U21 ( .A1(n373), .A2(n125), .A3(n75), .ZN(instr_addr_o[18]) );
  NAND2_X1 U22 ( .A1(branch_addr_i[18]), .A2(n153), .ZN(n373) );
  NAND3_X1 U23 ( .A1(n374), .A2(n149), .A3(n148), .ZN(instr_addr_o[28]) );
  NAND2_X1 U24 ( .A1(branch_addr_i[28]), .A2(n103), .ZN(n374) );
  NAND3_X1 U25 ( .A1(n378), .A2(n105), .A3(n104), .ZN(instr_addr_o[17]) );
  NAND2_X1 U34 ( .A1(branch_addr_i[17]), .A2(n103), .ZN(n378) );
  NAND3_X1 U35 ( .A1(n383), .A2(n58), .A3(n167), .ZN(instr_addr_o[31]) );
  AOI22_X1 U38 ( .A1(n314), .A2(hwlp_addr_i[9]), .B1(n163), .B2(n24), .ZN(n154) );
  CLKBUF_X3 U44 ( .A(n87), .Z(n308) );
  CLKBUF_X1 U48 ( .A(branch_i), .Z(n298) );
  CLKBUF_X1 U50 ( .A(instr_addr_o[11]), .Z(n379) );
  INV_X2 U51 ( .A(n107), .ZN(n162) );
  CLKBUF_X1 U53 ( .A(instr_addr_o[28]), .Z(n380) );
  CLKBUF_X1 U54 ( .A(instr_addr_o[16]), .Z(n56) );
  CLKBUF_X1 U60 ( .A(instr_addr_o[26]), .Z(n55) );
  NAND3_X1 U74 ( .A1(n385), .A2(n129), .A3(n130), .ZN(instr_addr_o[22]) );
  NAND2_X1 U88 ( .A1(branch_addr_i[31]), .A2(n103), .ZN(n383) );
  NAND3_X1 U91 ( .A1(n384), .A2(n70), .A3(n71), .ZN(instr_addr_o[12]) );
  NAND2_X1 U92 ( .A1(branch_addr_i[12]), .A2(n159), .ZN(n384) );
  NAND2_X1 U98 ( .A1(branch_addr_i[22]), .A2(n159), .ZN(n385) );
  NAND2_X1 U122 ( .A1(n102), .A2(n101), .ZN(instr_addr_o[30]) );
  NAND2_X1 U132 ( .A1(branch_addr_i[30]), .A2(n159), .ZN(n102) );
  NAND4_X1 U179 ( .A1(n386), .A2(n185), .A3(n184), .A4(n186), .ZN(instr_req_o)
         );
  NAND2_X1 U208 ( .A1(prefetch_i), .A2(n181), .ZN(n386) );
  NAND2_X1 U214 ( .A1(n317), .A2(n316), .ZN(n387) );
  NOR2_X1 U227 ( .A1(n221), .A2(n166), .ZN(n388) );
  INV_X1 U228 ( .A(n367), .ZN(n711) );
  INV_X1 U763 ( .A(n306), .ZN(n712) );
  INV_X1 U764 ( .A(n313), .ZN(n713) );
  INV_X1 U766 ( .A(n329), .ZN(n716) );
  INV_X1 U767 ( .A(n326), .ZN(n717) );
  INV_X1 U768 ( .A(n324), .ZN(n718) );
  INV_X1 U769 ( .A(n323), .ZN(n719) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_33 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_32 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_31 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_30 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_29 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_28 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_27 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_26 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_25 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_24 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_23 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_22 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_21 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_20 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_19 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_18 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_17 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_16 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_15 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_14 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_13 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_12 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_11 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_10 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_9 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_8 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_7 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_6 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_5 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_4 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_3 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_2 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_1 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_0 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_load_store_unit_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1768, net1771;
  assign net1768 = EN;
  assign net1771 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1768), .SE(net1771), .GCK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_load_store_unit_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1768, net1771;
  assign net1768 = EN;
  assign net1771 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1768), .SE(net1771), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_ex_stage_FPU0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_DIV0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_0 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net15, net18;
  assign net15 = EN;
  assign net18 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net15), .SE(net18), .GCK(ENCLK) );
endmodule


module riscv_mult_SHARED_DSP_MULT0 ( clk, rst_n, enable_i, operator_i, 
        short_signed_i, op_a_i, op_b_i, op_c_i, imm_i, dot_signed_i, 
        dot_op_a_i, dot_op_b_i, dot_op_c_i, is_clpx_i, clpx_shift_i, 
        clpx_img_i, result_o, multicycle_o, ready_o, ex_ready_i, 
        short_subword_i_BAR );
  input [2:0] operator_i;
  input [1:0] short_signed_i;
  input [31:0] op_a_i;
  input [31:0] op_b_i;
  input [31:0] op_c_i;
  input [4:0] imm_i;
  input [1:0] dot_signed_i;
  input [31:0] dot_op_a_i;
  input [31:0] dot_op_b_i;
  input [31:0] dot_op_c_i;
  input [1:0] clpx_shift_i;
  output [31:0] result_o;
  input clk, rst_n, enable_i, is_clpx_i, clpx_img_i, ex_ready_i,
         short_subword_i_BAR;
  output multicycle_o, ready_o;
  wire   mulh_carry_q, n464, n465, n466, n467, n2, n4, n5, n6, n10, n12, n15,
         n16, n17, n19, n20, n21, n22, n23, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n109, n110, n111, n113, n114,
         n115, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n128, n129, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6097, n6098, n6099, n6100, n6101, n6102, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160;
  wire   [2:0] mulh_CS;

  NOR2_X1 U6 ( .A1(n2058), .A2(n2057), .ZN(n2768) );
  NAND2_X2 U7 ( .A1(n2876), .A2(n5922), .ZN(n3128) );
  AOI21_X2 U18 ( .B1(n1026), .B2(n813), .A(n812), .ZN(n979) );
  OAI21_X1 U20 ( .B1(n6126), .B2(n2874), .A(n2), .ZN(n145) );
  NAND2_X1 U21 ( .A1(n6126), .A2(op_b_i[1]), .ZN(n2) );
  XNOR2_X1 U23 ( .A(n4), .B(n262), .ZN(n259) );
  XNOR2_X1 U24 ( .A(n264), .B(n263), .ZN(n4) );
  XNOR2_X1 U26 ( .A(n1023), .B(n5), .ZN(n4977) );
  AND2_X1 U27 ( .A1(n1025), .A2(n1039), .ZN(n5) );
  MUX2_X1 U33 ( .A(op_b_i[29]), .B(op_b_i[13]), .S(n146), .Z(n897) );
  INV_X1 U36 ( .A(n1608), .ZN(n69) );
  BUF_X1 U37 ( .A(n949), .Z(n70) );
  BUF_X1 U38 ( .A(n1128), .Z(n4587) );
  CLKBUF_X2 U39 ( .A(n1095), .Z(n16) );
  CLKBUF_X2 U40 ( .A(n1117), .Z(n4683) );
  NAND2_X2 U41 ( .A1(n2398), .A2(n6010), .ZN(n2867) );
  BUF_X1 U42 ( .A(n1130), .Z(n58) );
  INV_X1 U44 ( .A(n41), .ZN(n19) );
  INV_X1 U45 ( .A(n43), .ZN(n21) );
  INV_X1 U48 ( .A(n42), .ZN(n20) );
  INV_X2 U49 ( .A(n4137), .ZN(n10) );
  NAND2_X1 U51 ( .A1(n5083), .A2(n23), .ZN(n5114) );
  NAND2_X2 U52 ( .A1(n2402), .A2(n2401), .ZN(n2585) );
  NAND2_X2 U55 ( .A1(n4337), .A2(n5635), .ZN(n3241) );
  INV_X1 U56 ( .A(n3402), .ZN(n26) );
  BUF_X1 U59 ( .A(n1087), .Z(n1123) );
  AOI211_X1 U62 ( .C1(n2831), .C2(n5348), .A(n5023), .B(n5346), .ZN(n5604) );
  AND3_X1 U63 ( .A1(n2283), .A2(n86), .A3(n85), .ZN(n5575) );
  AND3_X1 U64 ( .A1(n1767), .A2(n4916), .A3(n1766), .ZN(n2273) );
  NOR2_X1 U65 ( .A1(n2060), .A2(n2059), .ZN(n2775) );
  NOR2_X1 U66 ( .A1(n635), .A2(n634), .ZN(n2305) );
  NAND2_X1 U68 ( .A1(n1133), .A2(n2112), .ZN(n2113) );
  BUF_X2 U70 ( .A(n1098), .Z(n2147) );
  BUF_X2 U71 ( .A(n114), .Z(n542) );
  BUF_X2 U72 ( .A(n128), .Z(n779) );
  BUF_X2 U73 ( .A(n113), .Z(n653) );
  BUF_X2 U74 ( .A(n125), .Z(n730) );
  BUF_X2 U75 ( .A(n1113), .Z(n17) );
  MUX2_X1 U77 ( .A(op_a_i[16]), .B(op_a_i[0]), .S(n149), .Z(n199) );
  INV_X1 U78 ( .A(n40), .ZN(n52) );
  INV_X1 U79 ( .A(n44), .ZN(n51) );
  INV_X2 U80 ( .A(n6101), .ZN(n5796) );
  NAND2_X1 U81 ( .A1(n2868), .A2(n5936), .ZN(n5934) );
  AND2_X1 U82 ( .A1(n5115), .A2(dot_signed_i[0]), .ZN(n5085) );
  INV_X1 U86 ( .A(n3533), .ZN(n63) );
  INV_X1 U88 ( .A(n67), .ZN(n68) );
  INV_X1 U89 ( .A(n3411), .ZN(n61) );
  INV_X1 U90 ( .A(n71), .ZN(n72) );
  INV_X1 U91 ( .A(n2486), .ZN(n60) );
  INV_X1 U93 ( .A(n1089), .ZN(n23) );
  INV_X2 U98 ( .A(n2840), .ZN(n2525) );
  NAND2_X1 U99 ( .A1(n2553), .A2(n3511), .ZN(n3514) );
  NAND2_X1 U100 ( .A1(n2419), .A2(n3715), .ZN(n3717) );
  NAND2_X1 U102 ( .A1(n2405), .A2(n3711), .ZN(n3713) );
  NAND2_X1 U104 ( .A1(n2849), .A2(n3534), .ZN(n3510) );
  NAND2_X1 U105 ( .A1(n2981), .A2(n6034), .ZN(n6032) );
  INV_X2 U107 ( .A(n2442), .ZN(n25) );
  INV_X2 U108 ( .A(n3386), .ZN(n27) );
  INV_X2 U109 ( .A(n2847), .ZN(n28) );
  INV_X2 U110 ( .A(op_b_i[0]), .ZN(n5635) );
  INV_X2 U112 ( .A(n3016), .ZN(n30) );
  NAND2_X2 U116 ( .A1(n6115), .A2(n122), .ZN(n991) );
  NAND2_X1 U117 ( .A1(n32), .A2(n31), .ZN(n705) );
  NAND2_X1 U118 ( .A1(n657), .A2(n656), .ZN(n31) );
  OAI21_X1 U119 ( .B1(n657), .B2(n656), .A(n655), .ZN(n32) );
  XNOR2_X1 U120 ( .A(n33), .B(n657), .ZN(n670) );
  XNOR2_X1 U121 ( .A(n655), .B(n656), .ZN(n33) );
  XNOR2_X1 U122 ( .A(n848), .B(n123), .ZN(n34) );
  XNOR2_X1 U123 ( .A(n848), .B(n123), .ZN(n35) );
  XNOR2_X1 U124 ( .A(n848), .B(n123), .ZN(n922) );
  XNOR2_X1 U125 ( .A(n1000), .B(n46), .ZN(n4962) );
  OAI21_X1 U126 ( .B1(n89), .B2(n87), .A(n94), .ZN(n93) );
  OR2_X1 U127 ( .A1(n1400), .A2(n88), .ZN(n87) );
  INV_X1 U128 ( .A(n1112), .ZN(n88) );
  OAI21_X1 U129 ( .B1(n991), .B2(n160), .A(n47), .ZN(n76) );
  AOI22_X1 U130 ( .A1(n76), .A2(n74), .B1(n195), .B2(n194), .ZN(n73) );
  OR2_X1 U131 ( .A1(n195), .A2(n194), .ZN(n74) );
  CLKBUF_X1 U132 ( .A(n969), .Z(n2713) );
  XNOR2_X1 U133 ( .A(n1067), .B(n45), .ZN(n4956) );
  AOI21_X1 U134 ( .B1(n2292), .B2(n1064), .A(n1063), .ZN(n1067) );
  NOR2_X1 U135 ( .A1(n2831), .A2(n6095), .ZN(n6098) );
  OAI21_X1 U136 ( .B1(n1887), .B2(n1886), .A(n93), .ZN(n92) );
  OAI21_X1 U137 ( .B1(n207), .B2(n204), .A(n205), .ZN(n141) );
  XNOR2_X1 U138 ( .A(n93), .B(n90), .ZN(n1881) );
  XNOR2_X1 U139 ( .A(n1886), .B(n1887), .ZN(n90) );
  OR2_X1 U141 ( .A1(n680), .A2(n681), .ZN(n82) );
  XNOR2_X1 U142 ( .A(n76), .B(n75), .ZN(n307) );
  XNOR2_X1 U143 ( .A(n195), .B(n194), .ZN(n75) );
  XNOR2_X1 U144 ( .A(n217), .B(n216), .ZN(n239) );
  INV_X1 U145 ( .A(n73), .ZN(n238) );
  XNOR2_X1 U146 ( .A(n679), .B(n83), .ZN(n707) );
  XNOR2_X1 U147 ( .A(n680), .B(n681), .ZN(n83) );
  INV_X1 U148 ( .A(n2135), .ZN(n2131) );
  INV_X1 U149 ( .A(n283), .ZN(n279) );
  NOR2_X1 U150 ( .A1(n633), .A2(n632), .ZN(n2312) );
  NOR2_X1 U152 ( .A1(n637), .A2(n636), .ZN(n2298) );
  OR2_X1 U154 ( .A1(n5794), .A2(n5386), .ZN(n5203) );
  NOR2_X1 U155 ( .A1(n2796), .A2(n2795), .ZN(n4889) );
  INV_X1 U156 ( .A(n5345), .ZN(n5544) );
  OAI21_X1 U157 ( .B1(n2829), .B2(n4965), .A(n4964), .ZN(n5897) );
  OAI21_X1 U158 ( .B1(n5575), .B2(n5894), .A(n2666), .ZN(n2667) );
  AOI21_X1 U159 ( .B1(n5439), .B2(n5158), .A(n2765), .ZN(n2783) );
  INV_X1 U160 ( .A(n5602), .ZN(n5377) );
  INV_X1 U161 ( .A(n5427), .ZN(n5553) );
  INV_X2 U162 ( .A(n3889), .ZN(n5919) );
  XNOR2_X1 U164 ( .A(n12), .B(n3407), .ZN(n5108) );
  XOR2_X1 U165 ( .A(n2879), .B(op_a_i[5]), .Z(n37) );
  XNOR2_X1 U166 ( .A(n1916), .B(n1132), .ZN(n2112) );
  NOR2_X2 U167 ( .A1(n2285), .A2(n1116), .ZN(n38) );
  NAND2_X2 U168 ( .A1(n2872), .A2(n2871), .ZN(n5822) );
  INV_X1 U169 ( .A(is_clpx_i), .ZN(n2658) );
  INV_X2 U170 ( .A(n2658), .ZN(n1661) );
  INV_X2 U171 ( .A(n3900), .ZN(n5922) );
  XOR2_X1 U172 ( .A(n2879), .B(op_a_i[4]), .Z(n39) );
  XOR2_X1 U173 ( .A(n2879), .B(op_a_i[10]), .Z(n40) );
  XOR2_X1 U174 ( .A(n2879), .B(op_a_i[6]), .Z(n41) );
  XOR2_X1 U175 ( .A(n2879), .B(op_a_i[8]), .Z(n42) );
  XOR2_X1 U176 ( .A(n2879), .B(op_a_i[9]), .Z(n43) );
  XOR2_X1 U177 ( .A(n2879), .B(op_a_i[11]), .Z(n44) );
  AND2_X1 U178 ( .A1(n1066), .A2(n1065), .ZN(n45) );
  AND2_X1 U179 ( .A1(n999), .A2(n2684), .ZN(n46) );
  OR2_X1 U180 ( .A1(n159), .A2(n6115), .ZN(n47) );
  XOR2_X1 U181 ( .A(n897), .B(n121), .Z(n48) );
  NOR2_X2 U182 ( .A1(n2272), .A2(clpx_shift_i[1]), .ZN(n5519) );
  INV_X1 U183 ( .A(n2112), .ZN(n49) );
  INV_X1 U184 ( .A(n5108), .ZN(n53) );
  INV_X2 U185 ( .A(n5325), .ZN(n5302) );
  XNOR2_X2 U186 ( .A(n6119), .B(op_a_i[15]), .ZN(n5914) );
  XNOR2_X2 U187 ( .A(n6118), .B(op_a_i[14]), .ZN(n5844) );
  XNOR2_X2 U188 ( .A(dot_op_b_i[26]), .B(dot_op_b_i[25]), .ZN(n3711) );
  XNOR2_X2 U189 ( .A(dot_op_b_i[28]), .B(dot_op_b_i[27]), .ZN(n3715) );
  XNOR2_X2 U190 ( .A(dot_op_b_i[2]), .B(dot_op_b_i[1]), .ZN(n3549) );
  XNOR2_X2 U191 ( .A(dot_op_b_i[10]), .B(dot_op_b_i[9]), .ZN(n3493) );
  XNOR2_X2 U192 ( .A(dot_op_b_i[12]), .B(dot_op_b_i[11]), .ZN(n3511) );
  XNOR2_X2 U193 ( .A(dot_op_b_i[4]), .B(dot_op_b_i[3]), .ZN(n3536) );
  XNOR2_X2 U194 ( .A(dot_op_b_i[14]), .B(dot_op_b_i[13]), .ZN(n3534) );
  XNOR2_X2 U195 ( .A(op_b_i[22]), .B(op_b_i[21]), .ZN(n5983) );
  XOR2_X1 U196 ( .A(n57), .B(n1111), .Z(n5112) );
  XNOR2_X1 U198 ( .A(n6118), .B(op_a_i[13]), .ZN(n65) );
  XNOR2_X1 U199 ( .A(n6118), .B(op_a_i[13]), .ZN(n66) );
  NOR2_X2 U201 ( .A1(clpx_shift_i[0]), .A2(clpx_shift_i[1]), .ZN(n5521) );
  INV_X1 U202 ( .A(n5999), .ZN(n67) );
  XNOR2_X1 U203 ( .A(n12), .B(dot_op_a_i[19]), .ZN(n1916) );
  OAI21_X1 U204 ( .B1(n146), .B2(n6073), .A(n120), .ZN(n949) );
  INV_X2 U205 ( .A(n5327), .ZN(n5304) );
  XNOR2_X2 U206 ( .A(op_b_i[18]), .B(op_b_i[17]), .ZN(n6034) );
  XNOR2_X2 U207 ( .A(n3312), .B(dot_op_a_i[15]), .ZN(n5116) );
  XNOR2_X2 U208 ( .A(n5108), .B(n17), .ZN(n5109) );
  XNOR2_X2 U209 ( .A(n167), .B(n949), .ZN(n2675) );
  AND3_X1 U210 ( .A1(n949), .A2(n166), .A3(short_signed_i[1]), .ZN(n167) );
  XNOR2_X2 U211 ( .A(op_b_i[16]), .B(op_b_i[15]), .ZN(n5917) );
  XNOR2_X2 U212 ( .A(n2879), .B(op_a_i[2]), .ZN(n5848) );
  XNOR2_X2 U213 ( .A(n2879), .B(op_a_i[1]), .ZN(n6002) );
  XNOR2_X2 U214 ( .A(op_b_i[14]), .B(op_b_i[13]), .ZN(n5927) );
  XNOR2_X2 U215 ( .A(dot_op_a_i[11]), .B(dot_op_a_i[12]), .ZN(n4829) );
  XNOR2_X2 U216 ( .A(dot_op_a_i[5]), .B(dot_op_a_i[6]), .ZN(n2246) );
  XNOR2_X2 U217 ( .A(dot_op_a_i[14]), .B(dot_op_a_i[13]), .ZN(n5123) );
  XNOR2_X2 U218 ( .A(dot_op_a_i[2]), .B(dot_op_a_i[1]), .ZN(n1903) );
  XNOR2_X2 U219 ( .A(dot_op_a_i[8]), .B(dot_op_a_i[7]), .ZN(n4629) );
  XNOR2_X2 U220 ( .A(dot_op_a_i[9]), .B(dot_op_a_i[10]), .ZN(n4745) );
  XNOR2_X2 U221 ( .A(dot_op_a_i[3]), .B(dot_op_a_i[4]), .ZN(n2079) );
  XNOR2_X2 U222 ( .A(n1128), .B(n1085), .ZN(n4731) );
  INV_X1 U224 ( .A(n5936), .ZN(n71) );
  AND2_X1 U225 ( .A1(n5573), .A2(n5490), .ZN(n2780) );
  NAND2_X1 U226 ( .A1(n5578), .A2(n5427), .ZN(n2669) );
  NOR2_X1 U227 ( .A1(n1078), .A2(n77), .ZN(n5578) );
  NAND2_X1 U228 ( .A1(n79), .A2(n78), .ZN(n77) );
  NAND2_X1 U229 ( .A1(n5348), .A2(n5794), .ZN(n78) );
  INV_X1 U230 ( .A(n5346), .ZN(n79) );
  NOR2_X1 U231 ( .A1(n802), .A2(n801), .ZN(n1018) );
  NAND2_X1 U232 ( .A1(n81), .A2(n80), .ZN(n724) );
  NAND2_X1 U233 ( .A1(n680), .A2(n681), .ZN(n80) );
  NAND2_X1 U234 ( .A1(n679), .A2(n82), .ZN(n81) );
  INV_X1 U235 ( .A(clpx_img_i), .ZN(n84) );
  AOI21_X1 U236 ( .B1(n5097), .B2(n5096), .A(n5095), .ZN(n5147) );
  XNOR2_X2 U237 ( .A(n1081), .B(n1098), .ZN(n4660) );
  OAI21_X2 U238 ( .B1(n4962), .B2(n5554), .A(n1015), .ZN(n2829) );
  XNOR2_X1 U239 ( .A(n283), .B(n282), .ZN(n218) );
  NAND2_X1 U240 ( .A1(n84), .A2(is_clpx_i), .ZN(n1089) );
  NAND2_X1 U241 ( .A1(n5602), .A2(n5490), .ZN(n85) );
  NAND2_X1 U242 ( .A1(n5588), .A2(n5463), .ZN(n86) );
  INV_X1 U244 ( .A(n6114), .ZN(n89) );
  NAND2_X1 U245 ( .A1(n92), .A2(n91), .ZN(n1911) );
  NAND2_X1 U246 ( .A1(n1886), .A2(n1887), .ZN(n91) );
  OR2_X1 U247 ( .A1(n1817), .A2(n6114), .ZN(n94) );
  MUX2_X2 U251 ( .A(op_b_i[27]), .B(op_b_i[11]), .S(n146), .Z(n848) );
  AND2_X1 U252 ( .A1(n193), .A2(n192), .ZN(n95) );
  XOR2_X1 U253 ( .A(n192), .B(n193), .Z(n96) );
  AND2_X1 U254 ( .A1(n1849), .A2(n1848), .ZN(n97) );
  XOR2_X1 U255 ( .A(n1849), .B(n1848), .Z(n98) );
  AND2_X1 U256 ( .A1(n3581), .A2(n3582), .ZN(n99) );
  XOR2_X1 U257 ( .A(n3582), .B(n3581), .Z(n100) );
  AND2_X1 U258 ( .A1(n1073), .A2(n1072), .ZN(n101) );
  OR2_X1 U259 ( .A1(n806), .A2(n805), .ZN(n102) );
  AND2_X1 U260 ( .A1(n3607), .A2(n3608), .ZN(n103) );
  XOR2_X1 U261 ( .A(n3608), .B(n3607), .Z(n104) );
  OR2_X1 U262 ( .A1(n1441), .A2(n1442), .ZN(n105) );
  OR2_X1 U263 ( .A1(n4889), .A2(n5894), .ZN(n106) );
  OAI21_X1 U264 ( .B1(n217), .B2(n215), .A(n214), .ZN(n135) );
  INV_X1 U265 ( .A(n282), .ZN(n278) );
  INV_X1 U266 ( .A(n2134), .ZN(n2130) );
  XNOR2_X1 U267 ( .A(n1442), .B(n1441), .ZN(n1299) );
  XNOR2_X1 U268 ( .A(n218), .B(n281), .ZN(n286) );
  XNOR2_X1 U269 ( .A(n1440), .B(n1299), .ZN(n1763) );
  XNOR2_X1 U270 ( .A(n2135), .B(n2134), .ZN(n1997) );
  XNOR2_X1 U271 ( .A(n2133), .B(n1997), .ZN(n2062) );
  OR2_X1 U272 ( .A1(n4913), .A2(n4915), .ZN(n1766) );
  XNOR2_X1 U273 ( .A(n1074), .B(n101), .ZN(n4957) );
  NOR2_X1 U274 ( .A1(n109), .A2(mulh_CS[2]), .ZN(n969) );
  AND2_X1 U275 ( .A1(n38), .A2(dot_op_c_i[31]), .ZN(n6097) );
  AND2_X1 U276 ( .A1(n5588), .A2(n5490), .ZN(n2796) );
  OAI222_X1 U277 ( .A1(n5481), .A2(n5386), .B1(n5482), .B2(n5229), .C1(n5700), 
        .C2(n5261), .ZN(n5230) );
  NOR3_X1 U278 ( .A1(n6099), .A2(n6098), .A3(n6097), .ZN(n6100) );
  XNOR2_X1 U280 ( .A(n5147), .B(n5146), .ZN(n5522) );
  AOI21_X1 U281 ( .B1(n2825), .B2(n5158), .A(n2824), .ZN(n2826) );
  OAI211_X1 U283 ( .C1(n5553), .C2(n4893), .A(n106), .B(n2826), .ZN(
        result_o[4]) );
  NOR2_X1 U284 ( .A1(n5208), .A2(mulh_CS[2]), .ZN(multicycle_o) );
  NAND2_X1 U285 ( .A1(n969), .A2(short_subword_i_BAR), .ZN(n110) );
  MUX2_X1 U287 ( .A(op_b_i[18]), .B(op_b_i[2]), .S(n6126), .Z(n107) );
  MUX2_X1 U288 ( .A(op_b_i[19]), .B(op_b_i[3]), .S(n6126), .Z(n114) );
  OR2_X1 U291 ( .A1(n5218), .A2(n6109), .ZN(n5210) );
  NAND2_X1 U292 ( .A1(n5210), .A2(n109), .ZN(n144) );
  NAND2_X1 U293 ( .A1(n144), .A2(n110), .ZN(n149) );
  MUX2_X1 U294 ( .A(op_a_i[30]), .B(op_a_i[14]), .S(n149), .Z(n954) );
  XNOR2_X1 U295 ( .A(n542), .B(n954), .ZN(n131) );
  XNOR2_X1 U297 ( .A(n542), .B(n985), .ZN(n181) );
  OAI22_X1 U298 ( .A1(n6135), .A2(n131), .B1(n6132), .B2(n181), .ZN(n174) );
  MUX2_X1 U299 ( .A(op_b_i[22]), .B(op_b_i[6]), .S(n6126), .Z(n111) );
  MUX2_X1 U300 ( .A(op_b_i[23]), .B(op_b_i[7]), .S(n6126), .Z(n125) );
  MUX2_X1 U302 ( .A(op_b_i[21]), .B(op_b_i[5]), .S(n6126), .Z(n113) );
  MUX2_X1 U304 ( .A(op_a_i[26]), .B(op_a_i[10]), .S(n149), .Z(n846) );
  XNOR2_X1 U305 ( .A(n730), .B(n846), .ZN(n139) );
  MUX2_X1 U306 ( .A(op_a_i[27]), .B(op_a_i[11]), .S(n149), .Z(n874) );
  XNOR2_X1 U307 ( .A(n730), .B(n874), .ZN(n164) );
  OAI22_X1 U308 ( .A1(n737), .A2(n139), .B1(n6136), .B2(n164), .ZN(n173) );
  MUX2_X1 U309 ( .A(op_b_i[20]), .B(op_b_i[4]), .S(n6126), .Z(n115) );
  MUX2_X1 U312 ( .A(op_a_i[28]), .B(op_a_i[12]), .S(n149), .Z(n902) );
  XNOR2_X1 U313 ( .A(n653), .B(n902), .ZN(n133) );
  MUX2_X1 U314 ( .A(op_a_i[29]), .B(op_a_i[13]), .S(n149), .Z(n918) );
  XNOR2_X1 U315 ( .A(n653), .B(n918), .ZN(n165) );
  OAI22_X1 U316 ( .A1(n6155), .A2(n133), .B1(n6152), .B2(n165), .ZN(n172) );
  INV_X1 U317 ( .A(operator_i[0]), .ZN(n117) );
  INV_X1 U318 ( .A(operator_i[1]), .ZN(n5212) );
  NOR3_X1 U319 ( .A1(n117), .A2(n5212), .A3(operator_i[2]), .ZN(n150) );
  INV_X1 U320 ( .A(imm_i[1]), .ZN(n118) );
  NAND3_X1 U321 ( .A1(n150), .A2(imm_i[0]), .A3(n118), .ZN(n895) );
  INV_X1 U322 ( .A(imm_i[3]), .ZN(n522) );
  INV_X1 U323 ( .A(imm_i[2]), .ZN(n727) );
  NAND3_X1 U324 ( .A1(n522), .A2(n727), .A3(imm_i[4]), .ZN(n183) );
  NOR2_X1 U325 ( .A1(n895), .A2(n183), .ZN(n138) );
  INV_X1 U326 ( .A(imm_i[0]), .ZN(n119) );
  NAND3_X1 U327 ( .A1(n150), .A2(n118), .A3(n119), .ZN(n880) );
  NOR2_X1 U328 ( .A1(n880), .A2(n183), .ZN(n158) );
  NAND3_X1 U329 ( .A1(n150), .A2(imm_i[1]), .A3(n119), .ZN(n916) );
  NOR2_X1 U330 ( .A1(n916), .A2(n183), .ZN(n184) );
  XNOR2_X1 U331 ( .A(n184), .B(op_c_i[17]), .ZN(n170) );
  MUX2_X1 U332 ( .A(op_b_i[30]), .B(op_b_i[14]), .S(n146), .Z(n121) );
  INV_X1 U333 ( .A(op_b_i[31]), .ZN(n6073) );
  NAND2_X1 U334 ( .A1(n146), .A2(op_b_i[15]), .ZN(n120) );
  XOR2_X1 U335 ( .A(n121), .B(n949), .Z(n122) );
  MUX2_X1 U336 ( .A(op_a_i[18]), .B(op_a_i[2]), .S(n149), .Z(n532) );
  XNOR2_X1 U337 ( .A(n70), .B(n532), .ZN(n136) );
  MUX2_X1 U338 ( .A(op_a_i[19]), .B(op_a_i[3]), .S(n149), .Z(n517) );
  XNOR2_X1 U339 ( .A(n70), .B(n517), .ZN(n182) );
  OAI22_X1 U340 ( .A1(n991), .A2(n136), .B1(n6115), .B2(n182), .ZN(n169) );
  MUX2_X1 U341 ( .A(op_b_i[28]), .B(op_b_i[12]), .S(n6126), .Z(n123) );
  XOR2_X1 U342 ( .A(n123), .B(n897), .Z(n124) );
  MUX2_X1 U343 ( .A(op_a_i[20]), .B(op_a_i[4]), .S(n149), .Z(n645) );
  XNOR2_X1 U344 ( .A(n6), .B(n645), .ZN(n142) );
  MUX2_X1 U345 ( .A(op_a_i[21]), .B(op_a_i[5]), .S(n149), .Z(n690) );
  XNOR2_X1 U346 ( .A(n6), .B(n690), .ZN(n179) );
  OAI22_X1 U347 ( .A1(n921), .A2(n142), .B1(n35), .B2(n179), .ZN(n177) );
  MUX2_X1 U348 ( .A(op_b_i[24]), .B(op_b_i[8]), .S(n6126), .Z(n126) );
  MUX2_X1 U349 ( .A(op_b_i[25]), .B(op_b_i[9]), .S(n6126), .Z(n128) );
  MUX2_X1 U351 ( .A(op_a_i[24]), .B(op_a_i[8]), .S(n149), .Z(n782) );
  XNOR2_X1 U352 ( .A(n779), .B(n782), .ZN(n143) );
  MUX2_X1 U353 ( .A(op_a_i[25]), .B(op_a_i[9]), .S(n149), .Z(n822) );
  XNOR2_X1 U354 ( .A(n779), .B(n822), .ZN(n185) );
  OAI22_X1 U355 ( .A1(n831), .A2(n143), .B1(n832), .B2(n185), .ZN(n176) );
  MUX2_X1 U356 ( .A(op_b_i[26]), .B(op_b_i[10]), .S(n6126), .Z(n129) );
  MUX2_X1 U359 ( .A(op_a_i[22]), .B(op_a_i[6]), .S(n149), .Z(n714) );
  XNOR2_X1 U360 ( .A(n848), .B(n714), .ZN(n132) );
  MUX2_X1 U361 ( .A(op_a_i[23]), .B(op_a_i[7]), .S(n149), .Z(n734) );
  XNOR2_X1 U362 ( .A(n848), .B(n734), .ZN(n180) );
  OAI22_X1 U363 ( .A1(n870), .A2(n132), .B1(n6156), .B2(n180), .ZN(n175) );
  XNOR2_X1 U364 ( .A(n542), .B(n918), .ZN(n148) );
  OAI22_X1 U365 ( .A1(n6134), .A2(n148), .B1(n6132), .B2(n131), .ZN(n217) );
  XNOR2_X1 U366 ( .A(n848), .B(n690), .ZN(n202) );
  OAI22_X1 U367 ( .A1(n6158), .A2(n202), .B1(n6156), .B2(n132), .ZN(n215) );
  XNOR2_X1 U368 ( .A(n653), .B(n874), .ZN(n147) );
  OAI22_X1 U369 ( .A1(n6154), .A2(n147), .B1(n6152), .B2(n133), .ZN(n214) );
  NAND2_X1 U370 ( .A1(n217), .A2(n215), .ZN(n134) );
  NAND2_X1 U371 ( .A1(n135), .A2(n134), .ZN(n163) );
  MUX2_X1 U372 ( .A(op_a_i[17]), .B(op_a_i[1]), .S(n149), .Z(n541) );
  XNOR2_X1 U373 ( .A(n70), .B(n541), .ZN(n200) );
  OAI22_X1 U374 ( .A1(n991), .A2(n200), .B1(n6115), .B2(n136), .ZN(n207) );
  FA_X1 U375 ( .A(n138), .B(op_c_i[16]), .CI(n137), .CO(n171), .S(n204) );
  XNOR2_X1 U376 ( .A(n730), .B(n822), .ZN(n212) );
  OAI22_X1 U377 ( .A1(n737), .A2(n212), .B1(n6136), .B2(n139), .ZN(n205) );
  NAND2_X1 U378 ( .A1(n207), .A2(n204), .ZN(n140) );
  NAND2_X1 U379 ( .A1(n141), .A2(n140), .ZN(n162) );
  XNOR2_X1 U380 ( .A(n6), .B(n517), .ZN(n197) );
  OAI22_X1 U381 ( .A1(n921), .A2(n197), .B1(n35), .B2(n142), .ZN(n153) );
  XNOR2_X1 U382 ( .A(n779), .B(n734), .ZN(n208) );
  OAI22_X1 U383 ( .A1(n6151), .A2(n208), .B1(n6148), .B2(n143), .ZN(n152) );
  XNOR2_X1 U386 ( .A(n2673), .B(n533), .ZN(n187) );
  MUX2_X1 U387 ( .A(op_b_i[16]), .B(op_b_i[0]), .S(n6126), .Z(n526) );
  XNOR2_X1 U390 ( .A(n533), .B(n985), .ZN(n210) );
  OAI22_X1 U391 ( .A1(n187), .A2(n549), .B1(n552), .B2(n210), .ZN(n151) );
  XNOR2_X1 U392 ( .A(n653), .B(n846), .ZN(n154) );
  OAI22_X1 U393 ( .A1(n6155), .A2(n154), .B1(n6152), .B2(n147), .ZN(n306) );
  XNOR2_X1 U394 ( .A(n542), .B(n902), .ZN(n155) );
  OAI22_X1 U395 ( .A1(n6135), .A2(n155), .B1(n6132), .B2(n148), .ZN(n305) );
  AND2_X1 U396 ( .A1(n199), .A2(n48), .ZN(n300) );
  NAND3_X1 U397 ( .A1(n150), .A2(imm_i[1]), .A3(imm_i[0]), .ZN(n952) );
  NOR2_X1 U398 ( .A1(n727), .A2(imm_i[4]), .ZN(n462) );
  NAND2_X1 U399 ( .A1(n462), .A2(imm_i[3]), .ZN(n230) );
  NOR2_X1 U400 ( .A1(n952), .A2(n230), .ZN(n157) );
  NOR2_X1 U401 ( .A1(n916), .A2(n230), .ZN(n231) );
  XNOR2_X1 U402 ( .A(n533), .B(n918), .ZN(n232) );
  XNOR2_X1 U403 ( .A(n533), .B(n954), .ZN(n211) );
  OAI22_X1 U404 ( .A1(n552), .A2(n232), .B1(n211), .B2(n549), .ZN(n298) );
  FA_X1 U405 ( .A(n153), .B(n152), .CI(n151), .CO(n161), .S(n293) );
  XNOR2_X1 U406 ( .A(n779), .B(n690), .ZN(n235) );
  XNOR2_X1 U407 ( .A(n779), .B(n714), .ZN(n209) );
  OAI22_X1 U408 ( .A1(n831), .A2(n235), .B1(n6148), .B2(n209), .ZN(n297) );
  XNOR2_X1 U409 ( .A(n653), .B(n822), .ZN(n234) );
  OAI22_X1 U410 ( .A1(n686), .A2(n234), .B1(n6152), .B2(n154), .ZN(n296) );
  XNOR2_X1 U411 ( .A(n730), .B(n734), .ZN(n323) );
  XNOR2_X1 U412 ( .A(n730), .B(n782), .ZN(n213) );
  OAI22_X1 U413 ( .A1(n737), .A2(n323), .B1(n6136), .B2(n213), .ZN(n295) );
  XNOR2_X1 U414 ( .A(n6), .B(n541), .ZN(n228) );
  XNOR2_X1 U415 ( .A(n6), .B(n532), .ZN(n198) );
  OAI22_X1 U416 ( .A1(n921), .A2(n228), .B1(n922), .B2(n198), .ZN(n303) );
  XNOR2_X1 U417 ( .A(n542), .B(n874), .ZN(n227) );
  OAI22_X1 U418 ( .A1(n6134), .A2(n227), .B1(n6132), .B2(n155), .ZN(n302) );
  XNOR2_X1 U419 ( .A(n848), .B(n517), .ZN(n233) );
  XNOR2_X1 U420 ( .A(n848), .B(n645), .ZN(n203) );
  OAI22_X1 U421 ( .A1(n6159), .A2(n233), .B1(n6156), .B2(n203), .ZN(n301) );
  FA_X1 U422 ( .A(n157), .B(op_c_i[14]), .CI(n156), .CO(n195), .S(n299) );
  HA_X1 U423 ( .A(n158), .B(op_c_i[15]), .CO(n137), .S(n194) );
  INV_X1 U424 ( .A(n949), .ZN(n160) );
  OR2_X1 U425 ( .A1(n199), .A2(n160), .ZN(n159) );
  FA_X1 U426 ( .A(n163), .B(n162), .CI(n161), .CO(n261), .S(n245) );
  XNOR2_X1 U427 ( .A(n730), .B(n902), .ZN(n256) );
  OAI22_X1 U428 ( .A1(n6139), .A2(n164), .B1(n6136), .B2(n256), .ZN(n249) );
  XNOR2_X1 U429 ( .A(n653), .B(n954), .ZN(n268) );
  OAI22_X1 U430 ( .A1(n6155), .A2(n165), .B1(n6152), .B2(n268), .ZN(n248) );
  INV_X1 U431 ( .A(n532), .ZN(n168) );
  NOR2_X1 U432 ( .A1(n168), .A2(n2675), .ZN(n247) );
  FA_X1 U433 ( .A(n171), .B(n170), .CI(n169), .CO(n263), .S(n190) );
  FA_X1 U434 ( .A(n174), .B(n173), .CI(n172), .CO(n262), .S(n191) );
  FA_X1 U435 ( .A(n177), .B(n176), .CI(n175), .CO(n264), .S(n189) );
  XNOR2_X1 U436 ( .A(n6), .B(n714), .ZN(n254) );
  OAI22_X1 U437 ( .A1(n921), .A2(n179), .B1(n922), .B2(n254), .ZN(n277) );
  XNOR2_X1 U438 ( .A(n848), .B(n782), .ZN(n267) );
  OAI22_X1 U439 ( .A1(n870), .A2(n180), .B1(n6156), .B2(n267), .ZN(n276) );
  XNOR2_X1 U440 ( .A(n2673), .B(n542), .ZN(n269) );
  OAI22_X1 U441 ( .A1(n6134), .A2(n181), .B1(n269), .B2(n6132), .ZN(n275) );
  XNOR2_X1 U442 ( .A(n70), .B(n645), .ZN(n253) );
  OAI22_X1 U443 ( .A1(n991), .A2(n182), .B1(n6115), .B2(n253), .ZN(n273) );
  NOR2_X1 U444 ( .A1(n952), .A2(n183), .ZN(n252) );
  INV_X1 U445 ( .A(op_c_i[18]), .ZN(n251) );
  OR2_X1 U446 ( .A1(n184), .A2(op_c_i[17]), .ZN(n250) );
  XNOR2_X1 U447 ( .A(n779), .B(n846), .ZN(n255) );
  OAI22_X1 U448 ( .A1(n6150), .A2(n185), .B1(n6148), .B2(n255), .ZN(n271) );
  INV_X1 U449 ( .A(n541), .ZN(n186) );
  NOR2_X1 U450 ( .A1(n186), .A2(n2675), .ZN(n193) );
  AOI21_X1 U451 ( .B1(n552), .B2(n549), .A(n187), .ZN(n188) );
  INV_X1 U452 ( .A(n188), .ZN(n192) );
  FA_X1 U453 ( .A(n191), .B(n190), .CI(n189), .CO(n282), .S(n246) );
  INV_X1 U454 ( .A(n2675), .ZN(n196) );
  AND2_X1 U455 ( .A1(n199), .A2(n196), .ZN(n237) );
  OAI22_X1 U456 ( .A1(n921), .A2(n198), .B1(n35), .B2(n197), .ZN(n224) );
  XNOR2_X1 U457 ( .A(n70), .B(n199), .ZN(n201) );
  OAI22_X1 U458 ( .A1(n991), .A2(n201), .B1(n6115), .B2(n200), .ZN(n223) );
  OAI22_X1 U459 ( .A1(n6158), .A2(n203), .B1(n6156), .B2(n202), .ZN(n222) );
  XNOR2_X1 U460 ( .A(n205), .B(n204), .ZN(n206) );
  XNOR2_X1 U461 ( .A(n207), .B(n206), .ZN(n241) );
  OAI22_X1 U462 ( .A1(n6150), .A2(n209), .B1(n6148), .B2(n208), .ZN(n221) );
  OAI22_X1 U463 ( .A1(n552), .A2(n211), .B1(n210), .B2(n549), .ZN(n220) );
  OAI22_X1 U464 ( .A1(n6138), .A2(n213), .B1(n6136), .B2(n212), .ZN(n219) );
  XNOR2_X1 U465 ( .A(n215), .B(n214), .ZN(n216) );
  FA_X1 U466 ( .A(n221), .B(n220), .CI(n219), .CO(n240), .S(n338) );
  FA_X1 U467 ( .A(n224), .B(n223), .CI(n222), .CO(n236), .S(n337) );
  INV_X1 U468 ( .A(n6), .ZN(n226) );
  OR2_X1 U469 ( .A1(n199), .A2(n226), .ZN(n225) );
  OAI22_X1 U470 ( .A1(n921), .A2(n226), .B1(n225), .B2(n35), .ZN(n335) );
  XNOR2_X1 U471 ( .A(n542), .B(n846), .ZN(n325) );
  OAI22_X1 U472 ( .A1(n562), .A2(n325), .B1(n560), .B2(n227), .ZN(n334) );
  XNOR2_X1 U473 ( .A(n6), .B(n199), .ZN(n229) );
  OAI22_X1 U474 ( .A1(n921), .A2(n229), .B1(n35), .B2(n228), .ZN(n333) );
  NOR2_X1 U475 ( .A1(n895), .A2(n230), .ZN(n321) );
  NOR2_X1 U476 ( .A1(n880), .A2(n230), .ZN(n355) );
  HA_X1 U477 ( .A(n231), .B(op_c_i[13]), .CO(n156), .S(n331) );
  XNOR2_X1 U478 ( .A(n533), .B(n902), .ZN(n322) );
  OAI22_X1 U479 ( .A1(n552), .A2(n322), .B1(n232), .B2(n549), .ZN(n330) );
  XNOR2_X1 U480 ( .A(n848), .B(n532), .ZN(n324) );
  OAI22_X1 U481 ( .A1(n870), .A2(n324), .B1(n871), .B2(n233), .ZN(n329) );
  XNOR2_X1 U482 ( .A(n653), .B(n782), .ZN(n353) );
  OAI22_X1 U483 ( .A1(n686), .A2(n353), .B1(n687), .B2(n234), .ZN(n328) );
  XNOR2_X1 U484 ( .A(n779), .B(n645), .ZN(n326) );
  OAI22_X1 U485 ( .A1(n6150), .A2(n326), .B1(n6148), .B2(n235), .ZN(n327) );
  FA_X1 U486 ( .A(n238), .B(n237), .CI(n236), .CO(n243), .S(n311) );
  FA_X1 U487 ( .A(n241), .B(n240), .CI(n239), .CO(n242), .S(n310) );
  FA_X1 U488 ( .A(n96), .B(n243), .CI(n242), .CO(n281), .S(n290) );
  FA_X1 U489 ( .A(n246), .B(n245), .CI(n244), .CO(n288), .S(n289) );
  FA_X1 U490 ( .A(n249), .B(n248), .CI(n247), .CO(n669), .S(n260) );
  FA_X1 U491 ( .A(n252), .B(n251), .CI(n250), .CO(n650), .S(n272) );
  NAND3_X1 U492 ( .A1(n522), .A2(imm_i[2]), .A3(imm_i[4]), .ZN(n725) );
  NOR2_X1 U493 ( .A1(n880), .A2(n725), .ZN(n665) );
  XNOR2_X1 U494 ( .A(n690), .B(n70), .ZN(n664) );
  OAI22_X1 U495 ( .A1(n991), .A2(n253), .B1(n6115), .B2(n664), .ZN(n648) );
  XNOR2_X1 U496 ( .A(n6), .B(n734), .ZN(n652) );
  OAI22_X1 U497 ( .A1(n921), .A2(n254), .B1(n922), .B2(n652), .ZN(n663) );
  XNOR2_X1 U498 ( .A(n779), .B(n874), .ZN(n647) );
  OAI22_X1 U499 ( .A1(n6151), .A2(n255), .B1(n6148), .B2(n647), .ZN(n662) );
  XNOR2_X1 U500 ( .A(n730), .B(n918), .ZN(n651) );
  OAI22_X1 U501 ( .A1(n6139), .A2(n256), .B1(n6136), .B2(n651), .ZN(n661) );
  FA_X1 U502 ( .A(n258), .B(n257), .CI(n95), .CO(n643), .S(n283) );
  FA_X1 U503 ( .A(n261), .B(n260), .CI(n259), .CO(n642), .S(n287) );
  OAI21_X1 U504 ( .B1(n264), .B2(n263), .A(n262), .ZN(n266) );
  NAND2_X1 U505 ( .A1(n264), .A2(n263), .ZN(n265) );
  NAND2_X1 U506 ( .A1(n266), .A2(n265), .ZN(n672) );
  XNOR2_X1 U507 ( .A(n848), .B(n822), .ZN(n666) );
  OAI22_X1 U508 ( .A1(n6159), .A2(n267), .B1(n6156), .B2(n666), .ZN(n660) );
  XNOR2_X1 U509 ( .A(n653), .B(n985), .ZN(n654) );
  OAI22_X1 U510 ( .A1(n6154), .A2(n268), .B1(n6152), .B2(n654), .ZN(n659) );
  AOI21_X1 U511 ( .B1(n6132), .B2(n6134), .A(n269), .ZN(n270) );
  INV_X1 U512 ( .A(n270), .ZN(n658) );
  FA_X1 U513 ( .A(n273), .B(n272), .CI(n271), .CO(n657), .S(n257) );
  INV_X1 U514 ( .A(n517), .ZN(n274) );
  NOR2_X1 U515 ( .A1(n274), .A2(n2675), .ZN(n656) );
  FA_X1 U516 ( .A(n277), .B(n276), .CI(n275), .CO(n655), .S(n258) );
  NAND2_X1 U517 ( .A1(n279), .A2(n278), .ZN(n280) );
  NAND2_X1 U518 ( .A1(n281), .A2(n280), .ZN(n285) );
  NAND2_X1 U519 ( .A1(n283), .A2(n282), .ZN(n284) );
  NAND2_X1 U520 ( .A1(n285), .A2(n284), .ZN(n673) );
  FA_X1 U521 ( .A(n288), .B(n287), .CI(n286), .CO(n636), .S(n635) );
  NOR2_X1 U522 ( .A1(n2305), .A2(n2298), .ZN(n639) );
  FA_X1 U523 ( .A(n291), .B(n290), .CI(n289), .CO(n634), .S(n633) );
  FA_X1 U524 ( .A(n294), .B(n293), .CI(n292), .CO(n244), .S(n315) );
  FA_X1 U525 ( .A(n297), .B(n296), .CI(n295), .CO(n309), .S(n362) );
  FA_X1 U526 ( .A(n300), .B(n299), .CI(n298), .CO(n304), .S(n361) );
  FA_X1 U527 ( .A(n303), .B(n302), .CI(n301), .CO(n308), .S(n360) );
  FA_X1 U528 ( .A(n306), .B(n305), .CI(n304), .CO(n294), .S(n340) );
  FA_X1 U529 ( .A(n309), .B(n308), .CI(n307), .CO(n292), .S(n339) );
  FA_X1 U530 ( .A(n312), .B(n311), .CI(n310), .CO(n291), .S(n313) );
  FA_X1 U531 ( .A(n315), .B(n314), .CI(n313), .CO(n632), .S(n631) );
  FA_X1 U532 ( .A(n318), .B(n317), .CI(n316), .CO(n336), .S(n365) );
  INV_X1 U533 ( .A(n922), .ZN(n319) );
  AND2_X1 U534 ( .A1(n199), .A2(n319), .ZN(n350) );
  FA_X1 U535 ( .A(n321), .B(op_c_i[12]), .CI(n320), .CO(n332), .S(n349) );
  XNOR2_X1 U536 ( .A(n533), .B(n874), .ZN(n356) );
  OAI22_X1 U537 ( .A1(n552), .A2(n356), .B1(n322), .B2(n549), .ZN(n348) );
  XNOR2_X1 U538 ( .A(n730), .B(n714), .ZN(n351) );
  OAI22_X1 U539 ( .A1(n6138), .A2(n351), .B1(n6136), .B2(n323), .ZN(n358) );
  XNOR2_X1 U540 ( .A(n848), .B(n541), .ZN(n346) );
  OAI22_X1 U541 ( .A1(n6159), .A2(n346), .B1(n6156), .B2(n324), .ZN(n378) );
  XNOR2_X1 U542 ( .A(n542), .B(n822), .ZN(n345) );
  OAI22_X1 U543 ( .A1(n6135), .A2(n345), .B1(n6132), .B2(n325), .ZN(n377) );
  XNOR2_X1 U544 ( .A(n779), .B(n517), .ZN(n342) );
  OAI22_X1 U545 ( .A1(n6150), .A2(n342), .B1(n6148), .B2(n326), .ZN(n376) );
  FA_X1 U546 ( .A(n329), .B(n328), .CI(n327), .CO(n316), .S(n384) );
  FA_X1 U547 ( .A(n332), .B(n331), .CI(n330), .CO(n317), .S(n383) );
  FA_X1 U548 ( .A(n335), .B(n334), .CI(n333), .CO(n318), .S(n382) );
  FA_X1 U549 ( .A(n338), .B(n337), .CI(n336), .CO(n312), .S(n413) );
  FA_X1 U550 ( .A(n341), .B(n340), .CI(n339), .CO(n314), .S(n412) );
  NOR2_X1 U551 ( .A1(n631), .A2(n630), .ZN(n2310) );
  NOR2_X1 U552 ( .A1(n2312), .A2(n2310), .ZN(n2304) );
  NAND2_X1 U553 ( .A1(n639), .A2(n2304), .ZN(n641) );
  XNOR2_X1 U554 ( .A(n779), .B(n532), .ZN(n366) );
  OAI22_X1 U555 ( .A1(n6151), .A2(n366), .B1(n6148), .B2(n342), .ZN(n396) );
  XNOR2_X1 U556 ( .A(n653), .B(n714), .ZN(n400) );
  XNOR2_X1 U557 ( .A(n653), .B(n734), .ZN(n354) );
  OAI22_X1 U558 ( .A1(n6154), .A2(n400), .B1(n6152), .B2(n354), .ZN(n395) );
  XNOR2_X1 U559 ( .A(n730), .B(n645), .ZN(n368) );
  XNOR2_X1 U560 ( .A(n730), .B(n690), .ZN(n352) );
  OAI22_X1 U561 ( .A1(n6139), .A2(n368), .B1(n6136), .B2(n352), .ZN(n394) );
  INV_X1 U562 ( .A(n848), .ZN(n344) );
  OR2_X1 U563 ( .A1(n199), .A2(n344), .ZN(n343) );
  OAI22_X1 U564 ( .A1(n6159), .A2(n344), .B1(n343), .B2(n6156), .ZN(n393) );
  XNOR2_X1 U565 ( .A(n542), .B(n782), .ZN(n367) );
  OAI22_X1 U566 ( .A1(n6135), .A2(n367), .B1(n6132), .B2(n345), .ZN(n392) );
  XNOR2_X1 U567 ( .A(n848), .B(n199), .ZN(n347) );
  OAI22_X1 U568 ( .A1(n6158), .A2(n347), .B1(n6156), .B2(n346), .ZN(n391) );
  FA_X1 U569 ( .A(n350), .B(n349), .CI(n348), .CO(n359), .S(n406) );
  OAI22_X1 U570 ( .A1(n6138), .A2(n352), .B1(n6136), .B2(n351), .ZN(n381) );
  OAI22_X1 U571 ( .A1(n6154), .A2(n354), .B1(n6152), .B2(n353), .ZN(n380) );
  NOR2_X1 U572 ( .A1(imm_i[4]), .A2(imm_i[2]), .ZN(n523) );
  NAND2_X1 U573 ( .A1(n523), .A2(imm_i[3]), .ZN(n397) );
  NOR2_X1 U574 ( .A1(n952), .A2(n397), .ZN(n371) );
  NOR2_X1 U575 ( .A1(n916), .A2(n397), .ZN(n398) );
  HA_X1 U576 ( .A(n355), .B(op_c_i[11]), .CO(n320), .S(n374) );
  XNOR2_X1 U577 ( .A(n533), .B(n846), .ZN(n372) );
  OAI22_X1 U578 ( .A1(n552), .A2(n372), .B1(n356), .B2(n549), .ZN(n373) );
  FA_X1 U579 ( .A(n359), .B(n358), .CI(n357), .CO(n364), .S(n385) );
  FA_X1 U580 ( .A(n362), .B(n361), .CI(n360), .CO(n341), .S(n416) );
  FA_X1 U581 ( .A(n365), .B(n364), .CI(n363), .CO(n414), .S(n415) );
  XNOR2_X1 U582 ( .A(n779), .B(n541), .ZN(n404) );
  OAI22_X1 U583 ( .A1(n6150), .A2(n404), .B1(n6148), .B2(n366), .ZN(n423) );
  XNOR2_X1 U584 ( .A(n542), .B(n734), .ZN(n403) );
  OAI22_X1 U585 ( .A1(n6135), .A2(n403), .B1(n6132), .B2(n367), .ZN(n422) );
  XNOR2_X1 U586 ( .A(n730), .B(n517), .ZN(n427) );
  OAI22_X1 U587 ( .A1(n6138), .A2(n427), .B1(n6136), .B2(n368), .ZN(n421) );
  INV_X1 U588 ( .A(n871), .ZN(n369) );
  AND2_X1 U589 ( .A1(n199), .A2(n369), .ZN(n426) );
  FA_X1 U590 ( .A(n371), .B(op_c_i[10]), .CI(n370), .CO(n375), .S(n425) );
  XNOR2_X1 U591 ( .A(n533), .B(n822), .ZN(n399) );
  OAI22_X1 U592 ( .A1(n552), .A2(n399), .B1(n372), .B2(n549), .ZN(n424) );
  FA_X1 U593 ( .A(n375), .B(n374), .CI(n373), .CO(n379), .S(n418) );
  FA_X1 U594 ( .A(n378), .B(n377), .CI(n376), .CO(n357), .S(n410) );
  FA_X1 U595 ( .A(n381), .B(n380), .CI(n379), .CO(n386), .S(n409) );
  FA_X1 U596 ( .A(n384), .B(n383), .CI(n382), .CO(n363), .S(n389) );
  FA_X1 U597 ( .A(n387), .B(n386), .CI(n385), .CO(n417), .S(n388) );
  OR2_X1 U598 ( .A1(n623), .A2(n622), .ZN(n2335) );
  FA_X1 U599 ( .A(n390), .B(n389), .CI(n388), .CO(n622), .S(n621) );
  FA_X1 U600 ( .A(n393), .B(n392), .CI(n391), .CO(n407), .S(n435) );
  FA_X1 U601 ( .A(n396), .B(n395), .CI(n394), .CO(n408), .S(n434) );
  NOR2_X1 U602 ( .A1(n895), .A2(n397), .ZN(n431) );
  NOR2_X1 U603 ( .A1(n880), .A2(n397), .ZN(n463) );
  HA_X1 U604 ( .A(n398), .B(op_c_i[9]), .CO(n370), .S(n440) );
  XNOR2_X1 U605 ( .A(n533), .B(n782), .ZN(n432) );
  OAI22_X1 U606 ( .A1(n552), .A2(n432), .B1(n399), .B2(n549), .ZN(n439) );
  XNOR2_X1 U607 ( .A(n653), .B(n690), .ZN(n428) );
  OAI22_X1 U608 ( .A1(n6154), .A2(n428), .B1(n6152), .B2(n400), .ZN(n437) );
  INV_X1 U609 ( .A(n779), .ZN(n402) );
  OR2_X1 U610 ( .A1(n199), .A2(n402), .ZN(n401) );
  OAI22_X1 U611 ( .A1(n6151), .A2(n402), .B1(n401), .B2(n6148), .ZN(n447) );
  XNOR2_X1 U612 ( .A(n542), .B(n714), .ZN(n443) );
  OAI22_X1 U613 ( .A1(n6134), .A2(n443), .B1(n6132), .B2(n403), .ZN(n446) );
  XNOR2_X1 U614 ( .A(n779), .B(n199), .ZN(n405) );
  OAI22_X1 U615 ( .A1(n6151), .A2(n405), .B1(n6148), .B2(n404), .ZN(n445) );
  FA_X1 U616 ( .A(n408), .B(n407), .CI(n406), .CO(n387), .S(n476) );
  FA_X1 U617 ( .A(n411), .B(n410), .CI(n409), .CO(n390), .S(n475) );
  NOR2_X1 U618 ( .A1(n621), .A2(n620), .ZN(n2333) );
  INV_X1 U619 ( .A(n2333), .ZN(n2339) );
  NAND2_X1 U620 ( .A1(n2335), .A2(n2339), .ZN(n2327) );
  FA_X1 U621 ( .A(n414), .B(n413), .CI(n412), .CO(n630), .S(n627) );
  FA_X1 U622 ( .A(n417), .B(n416), .CI(n415), .CO(n626), .S(n623) );
  NOR2_X1 U623 ( .A1(n627), .A2(n626), .ZN(n2328) );
  NOR2_X1 U624 ( .A1(n2327), .A2(n2328), .ZN(n629) );
  FA_X1 U625 ( .A(n420), .B(n419), .CI(n418), .CO(n411), .S(n480) );
  FA_X1 U626 ( .A(n423), .B(n422), .CI(n421), .CO(n420), .S(n450) );
  FA_X1 U627 ( .A(n426), .B(n425), .CI(n424), .CO(n419), .S(n449) );
  XNOR2_X1 U628 ( .A(n730), .B(n532), .ZN(n442) );
  OAI22_X1 U629 ( .A1(n6139), .A2(n442), .B1(n6136), .B2(n427), .ZN(n456) );
  XNOR2_X1 U630 ( .A(n653), .B(n645), .ZN(n444) );
  OAI22_X1 U631 ( .A1(n6155), .A2(n444), .B1(n6152), .B2(n428), .ZN(n455) );
  INV_X1 U632 ( .A(n832), .ZN(n429) );
  AND2_X1 U633 ( .A1(n199), .A2(n429), .ZN(n471) );
  FA_X1 U634 ( .A(n431), .B(op_c_i[8]), .CI(n430), .CO(n441), .S(n470) );
  XNOR2_X1 U635 ( .A(n533), .B(n734), .ZN(n468) );
  OAI22_X1 U636 ( .A1(n552), .A2(n468), .B1(n432), .B2(n549), .ZN(n469) );
  FA_X1 U637 ( .A(n435), .B(n434), .CI(n433), .CO(n477), .S(n478) );
  FA_X1 U638 ( .A(n438), .B(n437), .CI(n436), .CO(n433), .S(n453) );
  FA_X1 U639 ( .A(n441), .B(n440), .CI(n439), .CO(n438), .S(n474) );
  XNOR2_X1 U640 ( .A(n730), .B(n541), .ZN(n460) );
  OAI22_X1 U641 ( .A1(n6139), .A2(n460), .B1(n6136), .B2(n442), .ZN(n595) );
  XNOR2_X1 U642 ( .A(n542), .B(n690), .ZN(n459) );
  OAI22_X1 U643 ( .A1(n6134), .A2(n459), .B1(n6132), .B2(n443), .ZN(n594) );
  XNOR2_X1 U644 ( .A(n653), .B(n517), .ZN(n492) );
  OAI22_X1 U645 ( .A1(n6154), .A2(n492), .B1(n6152), .B2(n444), .ZN(n593) );
  FA_X1 U646 ( .A(n447), .B(n446), .CI(n445), .CO(n436), .S(n472) );
  FA_X1 U647 ( .A(n450), .B(n449), .CI(n448), .CO(n479), .S(n451) );
  NOR2_X1 U648 ( .A1(n614), .A2(n613), .ZN(n2352) );
  FA_X1 U649 ( .A(n453), .B(n452), .CI(n451), .CO(n613), .S(n612) );
  FA_X1 U650 ( .A(n456), .B(n455), .CI(n454), .CO(n448), .S(n589) );
  INV_X1 U651 ( .A(n730), .ZN(n458) );
  OR2_X1 U652 ( .A1(n199), .A2(n458), .ZN(n457) );
  OAI22_X1 U653 ( .A1(n6138), .A2(n458), .B1(n457), .B2(n6136), .ZN(n486) );
  XNOR2_X1 U654 ( .A(n542), .B(n645), .ZN(n481) );
  OAI22_X1 U655 ( .A1(n6135), .A2(n481), .B1(n6132), .B2(n459), .ZN(n485) );
  XNOR2_X1 U656 ( .A(n730), .B(n199), .ZN(n461) );
  OAI22_X1 U657 ( .A1(n6139), .A2(n461), .B1(n6136), .B2(n460), .ZN(n484) );
  NAND2_X1 U658 ( .A1(n462), .A2(n522), .ZN(n482) );
  NOR2_X1 U659 ( .A1(n952), .A2(n482), .ZN(n489) );
  NOR2_X1 U660 ( .A1(n916), .A2(n482), .ZN(n483) );
  HA_X1 U661 ( .A(n463), .B(op_c_i[7]), .CO(n430), .S(n495) );
  XNOR2_X1 U662 ( .A(n533), .B(n714), .ZN(n490) );
  OAI22_X1 U663 ( .A1(n552), .A2(n490), .B1(n468), .B2(n549), .ZN(n494) );
  FA_X1 U664 ( .A(n471), .B(n470), .CI(n469), .CO(n454), .S(n596) );
  FA_X1 U665 ( .A(n474), .B(n473), .CI(n472), .CO(n452), .S(n587) );
  NOR2_X1 U666 ( .A1(n612), .A2(n611), .ZN(n2350) );
  NOR2_X1 U667 ( .A1(n2352), .A2(n2350), .ZN(n2367) );
  FA_X1 U668 ( .A(n477), .B(n476), .CI(n475), .CO(n620), .S(n616) );
  FA_X1 U669 ( .A(n480), .B(n479), .CI(n478), .CO(n615), .S(n614) );
  OR2_X1 U670 ( .A1(n616), .A2(n615), .ZN(n2370) );
  NAND2_X1 U671 ( .A1(n2367), .A2(n2370), .ZN(n619) );
  XNOR2_X1 U672 ( .A(n653), .B(n541), .ZN(n503) );
  XNOR2_X1 U673 ( .A(n653), .B(n532), .ZN(n493) );
  OAI22_X1 U674 ( .A1(n6155), .A2(n503), .B1(n6152), .B2(n493), .ZN(n507) );
  XNOR2_X1 U675 ( .A(n542), .B(n517), .ZN(n502) );
  OAI22_X1 U676 ( .A1(n6135), .A2(n502), .B1(n6132), .B2(n481), .ZN(n506) );
  NOR2_X1 U677 ( .A1(n895), .A2(n482), .ZN(n516) );
  NOR2_X1 U678 ( .A1(n880), .A2(n482), .ZN(n547) );
  HA_X1 U679 ( .A(n483), .B(op_c_i[5]), .CO(n488), .S(n512) );
  XNOR2_X1 U680 ( .A(n533), .B(n645), .ZN(n518) );
  XNOR2_X1 U681 ( .A(n533), .B(n690), .ZN(n491) );
  OAI22_X1 U682 ( .A1(n552), .A2(n518), .B1(n491), .B2(n549), .ZN(n511) );
  FA_X1 U683 ( .A(n486), .B(n485), .CI(n484), .CO(n598), .S(n603) );
  INV_X1 U684 ( .A(n738), .ZN(n487) );
  AND2_X1 U685 ( .A1(n199), .A2(n487), .ZN(n499) );
  FA_X1 U686 ( .A(n489), .B(op_c_i[6]), .CI(n488), .CO(n496), .S(n498) );
  OAI22_X1 U687 ( .A1(n552), .A2(n491), .B1(n490), .B2(n549), .ZN(n497) );
  OAI22_X1 U688 ( .A1(n6154), .A2(n493), .B1(n6152), .B2(n492), .ZN(n591) );
  FA_X1 U689 ( .A(n496), .B(n495), .CI(n494), .CO(n597), .S(n590) );
  FA_X1 U690 ( .A(n499), .B(n498), .CI(n497), .CO(n592), .S(n510) );
  INV_X1 U691 ( .A(n653), .ZN(n501) );
  OR2_X1 U692 ( .A1(n199), .A2(n501), .ZN(n500) );
  OAI22_X1 U693 ( .A1(n6154), .A2(n501), .B1(n500), .B2(n6152), .ZN(n521) );
  XNOR2_X1 U694 ( .A(n542), .B(n532), .ZN(n559) );
  OAI22_X1 U695 ( .A1(n6134), .A2(n559), .B1(n6132), .B2(n502), .ZN(n520) );
  XNOR2_X1 U696 ( .A(n653), .B(n199), .ZN(n504) );
  OAI22_X1 U697 ( .A1(n6155), .A2(n504), .B1(n6152), .B2(n503), .ZN(n519) );
  FA_X1 U698 ( .A(n507), .B(n506), .CI(n505), .CO(n604), .S(n508) );
  OR2_X1 U699 ( .A1(n583), .A2(n582), .ZN(n2382) );
  FA_X1 U700 ( .A(n510), .B(n509), .CI(n508), .CO(n582), .S(n581) );
  FA_X1 U701 ( .A(n513), .B(n512), .CI(n511), .CO(n505), .S(n573) );
  INV_X1 U702 ( .A(n687), .ZN(n514) );
  AND2_X1 U703 ( .A1(n199), .A2(n514), .ZN(n565) );
  FA_X1 U704 ( .A(n516), .B(op_c_i[4]), .CI(n515), .CO(n513), .S(n564) );
  XNOR2_X1 U705 ( .A(n533), .B(n517), .ZN(n550) );
  OAI22_X1 U706 ( .A1(n552), .A2(n550), .B1(n518), .B2(n549), .ZN(n563) );
  FA_X1 U707 ( .A(n521), .B(n520), .CI(n519), .CO(n509), .S(n571) );
  OR2_X1 U708 ( .A1(n581), .A2(n580), .ZN(n2388) );
  NAND2_X1 U709 ( .A1(n2382), .A2(n2388), .ZN(n586) );
  NAND2_X1 U710 ( .A1(n523), .A2(n522), .ZN(n531) );
  NOR2_X1 U711 ( .A1(n916), .A2(n531), .ZN(n536) );
  XNOR2_X1 U712 ( .A(n533), .B(n541), .ZN(n534) );
  OAI22_X1 U713 ( .A1(n552), .A2(n199), .B1(n534), .B2(n549), .ZN(n535) );
  INV_X1 U714 ( .A(n533), .ZN(n524) );
  OR2_X1 U715 ( .A1(n199), .A2(n524), .ZN(n525) );
  NAND2_X1 U716 ( .A1(n525), .A2(n552), .ZN(n527) );
  OR2_X1 U717 ( .A1(n528), .A2(n527), .ZN(n5249) );
  NOR2_X1 U718 ( .A1(n895), .A2(n531), .ZN(n5253) );
  AND2_X1 U719 ( .A1(n199), .A2(n526), .ZN(n5252) );
  NAND2_X1 U720 ( .A1(n528), .A2(n527), .ZN(n5248) );
  INV_X1 U721 ( .A(n5248), .ZN(n529) );
  AOI21_X1 U722 ( .B1(n5249), .B2(n5250), .A(n529), .ZN(n5247) );
  INV_X1 U723 ( .A(n560), .ZN(n530) );
  AND2_X1 U724 ( .A1(n199), .A2(n530), .ZN(n546) );
  NOR2_X1 U725 ( .A1(n952), .A2(n531), .ZN(n548) );
  XNOR2_X1 U726 ( .A(n533), .B(n532), .ZN(n551) );
  OAI22_X1 U727 ( .A1(n552), .A2(n534), .B1(n551), .B2(n549), .ZN(n544) );
  FA_X1 U728 ( .A(n536), .B(op_c_i[1]), .CI(n535), .CO(n537), .S(n528) );
  NOR2_X1 U729 ( .A1(n538), .A2(n537), .ZN(n5243) );
  NAND2_X1 U730 ( .A1(n538), .A2(n537), .ZN(n5244) );
  OAI21_X1 U731 ( .B1(n5247), .B2(n5243), .A(n5244), .ZN(n2743) );
  INV_X1 U732 ( .A(n542), .ZN(n540) );
  OR2_X1 U733 ( .A1(n199), .A2(n540), .ZN(n539) );
  OAI22_X1 U734 ( .A1(n6135), .A2(n540), .B1(n539), .B2(n6132), .ZN(n568) );
  XNOR2_X1 U735 ( .A(n542), .B(n199), .ZN(n543) );
  XNOR2_X1 U736 ( .A(n542), .B(n541), .ZN(n561) );
  OAI22_X1 U737 ( .A1(n6134), .A2(n543), .B1(n6132), .B2(n561), .ZN(n567) );
  FA_X1 U738 ( .A(n546), .B(n545), .CI(n544), .CO(n566), .S(n538) );
  HA_X1 U739 ( .A(n547), .B(op_c_i[3]), .CO(n515), .S(n558) );
  HA_X1 U740 ( .A(n548), .B(op_c_i[2]), .CO(n557), .S(n545) );
  OAI22_X1 U741 ( .A1(n552), .A2(n551), .B1(n550), .B2(n549), .ZN(n556) );
  OR2_X1 U742 ( .A1(n554), .A2(n553), .ZN(n2742) );
  NAND2_X1 U743 ( .A1(n554), .A2(n553), .ZN(n2741) );
  INV_X1 U744 ( .A(n2741), .ZN(n555) );
  AOI21_X1 U745 ( .B1(n2743), .B2(n2742), .A(n555), .ZN(n2739) );
  FA_X1 U746 ( .A(n558), .B(n557), .CI(n556), .CO(n576), .S(n553) );
  OAI22_X1 U747 ( .A1(n6134), .A2(n561), .B1(n6132), .B2(n559), .ZN(n575) );
  FA_X1 U748 ( .A(n565), .B(n564), .CI(n563), .CO(n572), .S(n574) );
  FA_X1 U749 ( .A(n568), .B(n567), .CI(n566), .CO(n569), .S(n554) );
  NOR2_X1 U750 ( .A1(n570), .A2(n569), .ZN(n2736) );
  NAND2_X1 U751 ( .A1(n570), .A2(n569), .ZN(n2737) );
  OAI21_X1 U752 ( .B1(n2739), .B2(n2736), .A(n2737), .ZN(n2394) );
  FA_X1 U753 ( .A(n573), .B(n572), .CI(n571), .CO(n580), .S(n578) );
  FA_X1 U754 ( .A(n576), .B(n575), .CI(n574), .CO(n577), .S(n570) );
  OR2_X1 U755 ( .A1(n578), .A2(n577), .ZN(n2392) );
  NAND2_X1 U756 ( .A1(n578), .A2(n577), .ZN(n2391) );
  INV_X1 U757 ( .A(n2391), .ZN(n579) );
  AOI21_X1 U758 ( .B1(n2394), .B2(n2392), .A(n579), .ZN(n2383) );
  NAND2_X1 U759 ( .A1(n581), .A2(n580), .ZN(n2387) );
  INV_X1 U760 ( .A(n2387), .ZN(n2384) );
  NAND2_X1 U761 ( .A1(n583), .A2(n582), .ZN(n2381) );
  INV_X1 U762 ( .A(n2381), .ZN(n584) );
  AOI21_X1 U763 ( .B1(n2382), .B2(n2384), .A(n584), .ZN(n585) );
  OAI21_X1 U764 ( .B1(n586), .B2(n2383), .A(n585), .ZN(n2360) );
  FA_X1 U765 ( .A(n589), .B(n588), .CI(n587), .CO(n611), .S(n608) );
  FA_X1 U766 ( .A(n592), .B(n591), .CI(n590), .CO(n601), .S(n602) );
  FA_X1 U767 ( .A(n595), .B(n594), .CI(n593), .CO(n473), .S(n600) );
  FA_X1 U768 ( .A(n598), .B(n597), .CI(n596), .CO(n588), .S(n599) );
  NOR2_X1 U769 ( .A1(n608), .A2(n607), .ZN(n2361) );
  FA_X1 U770 ( .A(n601), .B(n600), .CI(n599), .CO(n607), .S(n606) );
  FA_X1 U771 ( .A(n604), .B(n603), .CI(n602), .CO(n605), .S(n583) );
  NOR2_X1 U772 ( .A1(n606), .A2(n605), .ZN(n2376) );
  NOR2_X1 U773 ( .A1(n2361), .A2(n2376), .ZN(n610) );
  NAND2_X1 U774 ( .A1(n606), .A2(n605), .ZN(n2377) );
  NAND2_X1 U775 ( .A1(n608), .A2(n607), .ZN(n2362) );
  OAI21_X1 U776 ( .B1(n2361), .B2(n2377), .A(n2362), .ZN(n609) );
  AOI21_X1 U777 ( .B1(n2360), .B2(n610), .A(n609), .ZN(n2349) );
  NAND2_X1 U778 ( .A1(n612), .A2(n611), .ZN(n2357) );
  NAND2_X1 U779 ( .A1(n614), .A2(n613), .ZN(n2353) );
  OAI21_X1 U780 ( .B1(n2352), .B2(n2357), .A(n2353), .ZN(n2366) );
  NAND2_X1 U781 ( .A1(n616), .A2(n615), .ZN(n2369) );
  INV_X1 U782 ( .A(n2369), .ZN(n617) );
  AOI21_X1 U783 ( .B1(n2366), .B2(n2370), .A(n617), .ZN(n618) );
  OAI21_X1 U784 ( .B1(n619), .B2(n2349), .A(n618), .ZN(n2325) );
  NAND2_X1 U785 ( .A1(n621), .A2(n620), .ZN(n2338) );
  INV_X1 U786 ( .A(n2338), .ZN(n625) );
  NAND2_X1 U787 ( .A1(n623), .A2(n622), .ZN(n2334) );
  INV_X1 U788 ( .A(n2334), .ZN(n624) );
  AOI21_X1 U789 ( .B1(n2335), .B2(n625), .A(n624), .ZN(n2326) );
  NAND2_X1 U790 ( .A1(n627), .A2(n626), .ZN(n2329) );
  OAI21_X1 U791 ( .B1(n2326), .B2(n2328), .A(n2329), .ZN(n628) );
  AOI21_X1 U792 ( .B1(n629), .B2(n2325), .A(n628), .ZN(n2294) );
  NAND2_X1 U793 ( .A1(n631), .A2(n630), .ZN(n2321) );
  NAND2_X1 U794 ( .A1(n633), .A2(n632), .ZN(n2313) );
  OAI21_X1 U795 ( .B1(n2312), .B2(n2321), .A(n2313), .ZN(n2303) );
  NAND2_X1 U796 ( .A1(n635), .A2(n634), .ZN(n2306) );
  NAND2_X1 U797 ( .A1(n637), .A2(n636), .ZN(n2299) );
  OAI21_X1 U798 ( .B1(n2298), .B2(n2306), .A(n2299), .ZN(n638) );
  AOI21_X1 U799 ( .B1(n639), .B2(n2303), .A(n638), .ZN(n640) );
  OAI21_X1 U800 ( .B1(n641), .B2(n2294), .A(n640), .ZN(n1002) );
  FA_X1 U801 ( .A(n644), .B(n643), .CI(n642), .CO(n710), .S(n675) );
  INV_X1 U802 ( .A(n645), .ZN(n646) );
  NOR2_X1 U803 ( .A1(n646), .A2(n2675), .ZN(n681) );
  XNOR2_X1 U804 ( .A(n779), .B(n902), .ZN(n684) );
  OAI22_X1 U805 ( .A1(n6150), .A2(n647), .B1(n6148), .B2(n684), .ZN(n680) );
  FA_X1 U806 ( .A(n650), .B(n649), .CI(n648), .CO(n679), .S(n668) );
  XNOR2_X1 U807 ( .A(n730), .B(n954), .ZN(n689) );
  OAI22_X1 U808 ( .A1(n6138), .A2(n651), .B1(n6136), .B2(n689), .ZN(n694) );
  XNOR2_X1 U809 ( .A(n6), .B(n782), .ZN(n682) );
  OAI22_X1 U810 ( .A1(n921), .A2(n652), .B1(n35), .B2(n682), .ZN(n693) );
  XNOR2_X1 U811 ( .A(n2673), .B(n653), .ZN(n685) );
  OAI22_X1 U812 ( .A1(n6155), .A2(n654), .B1(n685), .B2(n6152), .ZN(n692) );
  FA_X1 U813 ( .A(n660), .B(n659), .CI(n658), .CO(n704), .S(n671) );
  FA_X1 U814 ( .A(n663), .B(n662), .CI(n661), .CO(n703), .S(n667) );
  XNOR2_X1 U815 ( .A(n70), .B(n714), .ZN(n701) );
  OAI22_X1 U816 ( .A1(n991), .A2(n664), .B1(n6115), .B2(n701), .ZN(n697) );
  NOR2_X1 U817 ( .A1(n895), .A2(n725), .ZN(n700) );
  INV_X1 U818 ( .A(op_c_i[20]), .ZN(n699) );
  FA_X1 U819 ( .A(op_c_i[19]), .B(op_c_i[18]), .CI(n665), .CO(n698), .S(n649)
         );
  XNOR2_X1 U820 ( .A(n848), .B(n846), .ZN(n683) );
  OAI22_X1 U821 ( .A1(n6159), .A2(n666), .B1(n6156), .B2(n683), .ZN(n695) );
  FA_X1 U822 ( .A(n669), .B(n668), .CI(n667), .CO(n677), .S(n644) );
  FA_X1 U823 ( .A(n672), .B(n671), .CI(n670), .CO(n676), .S(n674) );
  FA_X1 U824 ( .A(n673), .B(n674), .CI(n675), .CO(n799), .S(n637) );
  NOR2_X1 U825 ( .A1(n800), .A2(n799), .ZN(n1016) );
  FA_X1 U826 ( .A(n678), .B(n677), .CI(n676), .CO(n798), .S(n708) );
  XNOR2_X1 U827 ( .A(n6), .B(n822), .ZN(n729) );
  OAI22_X1 U828 ( .A1(n921), .A2(n682), .B1(n922), .B2(n729), .ZN(n718) );
  XNOR2_X1 U829 ( .A(n848), .B(n874), .ZN(n745) );
  OAI22_X1 U830 ( .A1(n6159), .A2(n683), .B1(n6156), .B2(n745), .ZN(n717) );
  XNOR2_X1 U831 ( .A(n779), .B(n918), .ZN(n728) );
  OAI22_X1 U832 ( .A1(n6151), .A2(n684), .B1(n6148), .B2(n728), .ZN(n716) );
  AOI21_X1 U833 ( .B1(n6152), .B2(n686), .A(n685), .ZN(n688) );
  INV_X1 U834 ( .A(n688), .ZN(n754) );
  XNOR2_X1 U835 ( .A(n730), .B(n985), .ZN(n731) );
  OAI22_X1 U836 ( .A1(n6139), .A2(n689), .B1(n6136), .B2(n731), .ZN(n753) );
  INV_X1 U837 ( .A(n690), .ZN(n691) );
  NOR2_X1 U838 ( .A1(n691), .A2(n2675), .ZN(n752) );
  FA_X1 U839 ( .A(n694), .B(n693), .CI(n692), .CO(n721), .S(n706) );
  FA_X1 U840 ( .A(n697), .B(n696), .CI(n695), .CO(n720), .S(n702) );
  FA_X1 U841 ( .A(n700), .B(n699), .CI(n698), .CO(n713), .S(n696) );
  NOR2_X1 U842 ( .A1(n916), .A2(n725), .ZN(n726) );
  XNOR2_X1 U843 ( .A(n70), .B(n734), .ZN(n741) );
  OAI22_X1 U844 ( .A1(n991), .A2(n701), .B1(n6115), .B2(n741), .ZN(n711) );
  FA_X1 U845 ( .A(n704), .B(n703), .CI(n702), .CO(n759), .S(n678) );
  FA_X1 U846 ( .A(n707), .B(n706), .CI(n705), .CO(n758), .S(n709) );
  FA_X1 U847 ( .A(n710), .B(n709), .CI(n708), .CO(n801), .S(n800) );
  NOR2_X1 U848 ( .A1(n1016), .A2(n1018), .ZN(n1024) );
  FA_X1 U849 ( .A(n713), .B(n712), .CI(n711), .CO(n748), .S(n719) );
  INV_X1 U850 ( .A(n714), .ZN(n715) );
  NOR2_X1 U851 ( .A1(n715), .A2(n2675), .ZN(n747) );
  FA_X1 U852 ( .A(n718), .B(n717), .CI(n716), .CO(n746), .S(n723) );
  FA_X1 U853 ( .A(n721), .B(n720), .CI(n719), .CO(n765), .S(n760) );
  FA_X1 U854 ( .A(n724), .B(n723), .CI(n722), .CO(n764), .S(n797) );
  NOR2_X1 U855 ( .A1(n952), .A2(n725), .ZN(n743) );
  FA_X1 U856 ( .A(op_c_i[20]), .B(op_c_i[21]), .CI(n726), .CO(n742), .S(n712)
         );
  AND2_X1 U857 ( .A1(imm_i[4]), .A2(imm_i[3]), .ZN(n879) );
  NAND2_X1 U858 ( .A1(n879), .A2(n727), .ZN(n854) );
  NOR2_X1 U859 ( .A1(n880), .A2(n854), .ZN(n777) );
  XNOR2_X1 U860 ( .A(n782), .B(n70), .ZN(n740) );
  XNOR2_X1 U861 ( .A(n70), .B(n822), .ZN(n776) );
  OAI22_X1 U862 ( .A1(n991), .A2(n740), .B1(n6115), .B2(n776), .ZN(n773) );
  XNOR2_X1 U863 ( .A(n779), .B(n954), .ZN(n732) );
  OAI22_X1 U864 ( .A1(n6151), .A2(n728), .B1(n6148), .B2(n732), .ZN(n757) );
  XNOR2_X1 U865 ( .A(n6), .B(n846), .ZN(n733) );
  OAI22_X1 U866 ( .A1(n921), .A2(n729), .B1(n922), .B2(n733), .ZN(n756) );
  XNOR2_X1 U867 ( .A(n2673), .B(n730), .ZN(n736) );
  OAI22_X1 U868 ( .A1(n737), .A2(n731), .B1(n736), .B2(n738), .ZN(n755) );
  XNOR2_X1 U869 ( .A(n779), .B(n985), .ZN(n780) );
  OAI22_X1 U870 ( .A1(n6150), .A2(n732), .B1(n6148), .B2(n780), .ZN(n772) );
  XNOR2_X1 U871 ( .A(n848), .B(n902), .ZN(n744) );
  XNOR2_X1 U872 ( .A(n848), .B(n918), .ZN(n781) );
  OAI22_X1 U873 ( .A1(n6158), .A2(n744), .B1(n6156), .B2(n781), .ZN(n771) );
  XNOR2_X1 U874 ( .A(n6), .B(n874), .ZN(n778) );
  OAI22_X1 U875 ( .A1(n921), .A2(n733), .B1(n922), .B2(n778), .ZN(n770) );
  INV_X1 U876 ( .A(n734), .ZN(n735) );
  NOR2_X1 U877 ( .A1(n735), .A2(n2675), .ZN(n786) );
  AOI21_X1 U878 ( .B1(n6136), .B2(n6138), .A(n736), .ZN(n739) );
  INV_X1 U879 ( .A(n739), .ZN(n785) );
  OAI22_X1 U880 ( .A1(n991), .A2(n741), .B1(n6115), .B2(n740), .ZN(n751) );
  FA_X1 U881 ( .A(n743), .B(n4082), .CI(n742), .CO(n775), .S(n750) );
  OAI22_X1 U882 ( .A1(n6158), .A2(n745), .B1(n6156), .B2(n744), .ZN(n749) );
  FA_X1 U883 ( .A(n748), .B(n747), .CI(n746), .CO(n768), .S(n766) );
  FA_X1 U884 ( .A(n751), .B(n750), .CI(n749), .CO(n784), .S(n763) );
  FA_X1 U885 ( .A(n754), .B(n753), .CI(n752), .CO(n762), .S(n722) );
  FA_X1 U886 ( .A(n757), .B(n756), .CI(n755), .CO(n788), .S(n761) );
  FA_X1 U887 ( .A(n760), .B(n759), .CI(n758), .CO(n795), .S(n796) );
  FA_X1 U888 ( .A(n761), .B(n762), .CI(n763), .CO(n767), .S(n794) );
  FA_X1 U889 ( .A(n766), .B(n765), .CI(n764), .CO(n792), .S(n793) );
  FA_X1 U890 ( .A(n769), .B(n768), .CI(n767), .CO(n842), .S(n790) );
  FA_X1 U891 ( .A(n772), .B(n771), .CI(n770), .CO(n839), .S(n787) );
  FA_X1 U892 ( .A(n775), .B(n774), .CI(n773), .CO(n838), .S(n789) );
  XNOR2_X1 U893 ( .A(n70), .B(n846), .ZN(n827) );
  OAI22_X1 U894 ( .A1(n991), .A2(n776), .B1(n6115), .B2(n827), .ZN(n821) );
  NOR2_X1 U895 ( .A1(n895), .A2(n854), .ZN(n826) );
  INV_X1 U896 ( .A(op_c_i[24]), .ZN(n825) );
  FA_X1 U897 ( .A(op_c_i[22]), .B(op_c_i[23]), .CI(n777), .CO(n824), .S(n774)
         );
  XNOR2_X1 U898 ( .A(n6), .B(n902), .ZN(n829) );
  OAI22_X1 U899 ( .A1(n921), .A2(n778), .B1(n922), .B2(n829), .ZN(n819) );
  XNOR2_X1 U900 ( .A(n2673), .B(n779), .ZN(n830) );
  OAI22_X1 U901 ( .A1(n6151), .A2(n780), .B1(n830), .B2(n6148), .ZN(n836) );
  XNOR2_X1 U902 ( .A(n848), .B(n954), .ZN(n828) );
  OAI22_X1 U903 ( .A1(n6158), .A2(n781), .B1(n6156), .B2(n828), .ZN(n835) );
  INV_X1 U904 ( .A(n782), .ZN(n783) );
  NOR2_X1 U905 ( .A1(n783), .A2(n2675), .ZN(n834) );
  FA_X1 U906 ( .A(n786), .B(n785), .CI(n784), .CO(n817), .S(n769) );
  FA_X1 U907 ( .A(n789), .B(n788), .CI(n787), .CO(n816), .S(n791) );
  FA_X1 U908 ( .A(n792), .B(n791), .CI(n790), .CO(n807), .S(n806) );
  OR2_X1 U909 ( .A1(n808), .A2(n807), .ZN(n1034) );
  NAND2_X1 U910 ( .A1(n102), .A2(n1034), .ZN(n811) );
  FA_X1 U911 ( .A(n795), .B(n794), .CI(n793), .CO(n805), .S(n804) );
  FA_X1 U912 ( .A(n796), .B(n797), .CI(n798), .CO(n803), .S(n802) );
  NOR2_X1 U913 ( .A1(n804), .A2(n803), .ZN(n1040) );
  NOR2_X1 U914 ( .A1(n811), .A2(n1040), .ZN(n813) );
  NAND2_X1 U915 ( .A1(n1024), .A2(n813), .ZN(n2683) );
  INV_X1 U916 ( .A(n2683), .ZN(n815) );
  NAND2_X1 U917 ( .A1(n800), .A2(n799), .ZN(n2289) );
  NAND2_X1 U918 ( .A1(n802), .A2(n801), .ZN(n1019) );
  OAI21_X1 U919 ( .B1(n1018), .B2(n2289), .A(n1019), .ZN(n1026) );
  NAND2_X1 U920 ( .A1(n804), .A2(n803), .ZN(n1039) );
  NAND2_X1 U921 ( .A1(n806), .A2(n805), .ZN(n1044) );
  INV_X1 U922 ( .A(n1044), .ZN(n1027) );
  NAND2_X1 U923 ( .A1(n808), .A2(n807), .ZN(n1033) );
  INV_X1 U924 ( .A(n1033), .ZN(n809) );
  AOI21_X1 U925 ( .B1(n1034), .B2(n1027), .A(n809), .ZN(n810) );
  OAI21_X1 U926 ( .B1(n811), .B2(n1039), .A(n810), .ZN(n812) );
  INV_X1 U927 ( .A(n979), .ZN(n814) );
  AOI21_X1 U928 ( .B1(n1002), .B2(n815), .A(n814), .ZN(n1049) );
  FA_X1 U929 ( .A(n818), .B(n817), .CI(n816), .CO(n865), .S(n840) );
  FA_X1 U930 ( .A(n821), .B(n820), .CI(n819), .CO(n862), .S(n837) );
  INV_X1 U931 ( .A(n822), .ZN(n823) );
  NOR2_X1 U932 ( .A1(n823), .A2(n2675), .ZN(n861) );
  FA_X1 U933 ( .A(n826), .B(n825), .CI(n824), .CO(n852), .S(n820) );
  NOR2_X1 U934 ( .A1(n916), .A2(n854), .ZN(n855) );
  XNOR2_X1 U935 ( .A(n874), .B(n70), .ZN(n853) );
  OAI22_X1 U936 ( .A1(n991), .A2(n827), .B1(n6115), .B2(n853), .ZN(n850) );
  XNOR2_X1 U937 ( .A(n848), .B(n985), .ZN(n849) );
  OAI22_X1 U938 ( .A1(n6159), .A2(n828), .B1(n6156), .B2(n849), .ZN(n859) );
  XNOR2_X1 U939 ( .A(n6), .B(n918), .ZN(n856) );
  OAI22_X1 U940 ( .A1(n921), .A2(n829), .B1(n922), .B2(n856), .ZN(n858) );
  AOI21_X1 U941 ( .B1(n6148), .B2(n6150), .A(n830), .ZN(n833) );
  INV_X1 U942 ( .A(n833), .ZN(n857) );
  FA_X1 U943 ( .A(n836), .B(n835), .CI(n834), .CO(n844), .S(n818) );
  FA_X1 U944 ( .A(n839), .B(n838), .CI(n837), .CO(n843), .S(n841) );
  FA_X1 U945 ( .A(n842), .B(n841), .CI(n840), .CO(n930), .S(n808) );
  NOR2_X1 U946 ( .A1(n931), .A2(n930), .ZN(n1069) );
  INV_X1 U947 ( .A(n1069), .ZN(n1050) );
  FA_X1 U948 ( .A(n845), .B(n844), .CI(n843), .CO(n890), .S(n863) );
  INV_X1 U949 ( .A(n846), .ZN(n847) );
  NOR2_X1 U950 ( .A1(n847), .A2(n2675), .ZN(n887) );
  XNOR2_X1 U951 ( .A(n2673), .B(n848), .ZN(n869) );
  OAI22_X1 U952 ( .A1(n6158), .A2(n849), .B1(n869), .B2(n6156), .ZN(n886) );
  FA_X1 U953 ( .A(n852), .B(n851), .CI(n850), .CO(n885), .S(n860) );
  XNOR2_X1 U954 ( .A(n70), .B(n902), .ZN(n881) );
  OAI22_X1 U955 ( .A1(n991), .A2(n853), .B1(n6115), .B2(n881), .ZN(n884) );
  NOR2_X1 U956 ( .A1(n952), .A2(n854), .ZN(n878) );
  INV_X1 U957 ( .A(op_c_i[26]), .ZN(n877) );
  FA_X1 U958 ( .A(op_c_i[25]), .B(op_c_i[24]), .CI(n855), .CO(n876), .S(n851)
         );
  XNOR2_X1 U959 ( .A(n6), .B(n954), .ZN(n873) );
  OAI22_X1 U960 ( .A1(n921), .A2(n856), .B1(n35), .B2(n873), .ZN(n882) );
  FA_X1 U961 ( .A(n859), .B(n858), .CI(n857), .CO(n867), .S(n845) );
  FA_X1 U962 ( .A(n862), .B(n861), .CI(n860), .CO(n866), .S(n864) );
  FA_X1 U963 ( .A(n865), .B(n864), .CI(n863), .CO(n932), .S(n931) );
  OR2_X1 U964 ( .A1(n933), .A2(n932), .ZN(n1073) );
  NAND2_X1 U965 ( .A1(n1050), .A2(n1073), .ZN(n2672) );
  FA_X1 U966 ( .A(n868), .B(n867), .CI(n866), .CO(n909), .S(n888) );
  AOI21_X1 U967 ( .B1(n6156), .B2(n6159), .A(n869), .ZN(n872) );
  INV_X1 U968 ( .A(n872), .ZN(n906) );
  XNOR2_X1 U969 ( .A(n6), .B(n985), .ZN(n898) );
  OAI22_X1 U970 ( .A1(n921), .A2(n873), .B1(n922), .B2(n898), .ZN(n905) );
  INV_X1 U971 ( .A(n874), .ZN(n875) );
  NOR2_X1 U972 ( .A1(n875), .A2(n2675), .ZN(n904) );
  FA_X1 U973 ( .A(n878), .B(n877), .CI(n876), .CO(n901), .S(n883) );
  NAND2_X1 U974 ( .A1(n879), .A2(imm_i[2]), .ZN(n951) );
  NOR2_X1 U975 ( .A1(n880), .A2(n951), .ZN(n896) );
  XNOR2_X1 U976 ( .A(n70), .B(n918), .ZN(n894) );
  OAI22_X1 U977 ( .A1(n991), .A2(n881), .B1(n6115), .B2(n894), .ZN(n899) );
  FA_X1 U978 ( .A(n884), .B(n883), .CI(n882), .CO(n892), .S(n868) );
  FA_X1 U979 ( .A(n887), .B(n886), .CI(n885), .CO(n891), .S(n889) );
  FA_X1 U980 ( .A(n890), .B(n889), .CI(n888), .CO(n936), .S(n933) );
  NOR2_X1 U981 ( .A1(n937), .A2(n936), .ZN(n1054) );
  FA_X1 U982 ( .A(n893), .B(n892), .CI(n891), .CO(n929), .S(n907) );
  XNOR2_X1 U983 ( .A(n954), .B(n70), .ZN(n917) );
  OAI22_X1 U984 ( .A1(n991), .A2(n894), .B1(n6115), .B2(n917), .ZN(n926) );
  NOR2_X1 U985 ( .A1(n895), .A2(n951), .ZN(n915) );
  INV_X1 U986 ( .A(op_c_i[28]), .ZN(n914) );
  FA_X1 U987 ( .A(op_c_i[26]), .B(op_c_i[27]), .CI(n896), .CO(n913), .S(n900)
         );
  XNOR2_X1 U988 ( .A(n2673), .B(n6), .ZN(n920) );
  OAI22_X1 U989 ( .A1(n921), .A2(n898), .B1(n920), .B2(n922), .ZN(n924) );
  FA_X1 U990 ( .A(n901), .B(n900), .CI(n899), .CO(n912), .S(n893) );
  INV_X1 U991 ( .A(n902), .ZN(n903) );
  NOR2_X1 U992 ( .A1(n903), .A2(n2675), .ZN(n911) );
  FA_X1 U993 ( .A(n906), .B(n905), .CI(n904), .CO(n910), .S(n908) );
  FA_X1 U994 ( .A(n909), .B(n908), .CI(n907), .CO(n938), .S(n937) );
  OR2_X1 U995 ( .A1(n939), .A2(n938), .ZN(n1066) );
  FA_X1 U996 ( .A(n912), .B(n911), .CI(n910), .CO(n964), .S(n927) );
  FA_X1 U997 ( .A(n915), .B(n914), .CI(n913), .CO(n958), .S(n925) );
  NOR2_X1 U998 ( .A1(n916), .A2(n951), .ZN(n953) );
  XNOR2_X1 U999 ( .A(n70), .B(n985), .ZN(n950) );
  OAI22_X1 U1000 ( .A1(n991), .A2(n917), .B1(n6115), .B2(n950), .ZN(n956) );
  INV_X1 U1001 ( .A(n918), .ZN(n919) );
  NOR2_X1 U1002 ( .A1(n919), .A2(n2675), .ZN(n961) );
  AOI21_X1 U1003 ( .B1(n35), .B2(n921), .A(n920), .ZN(n923) );
  INV_X1 U1004 ( .A(n923), .ZN(n960) );
  FA_X1 U1005 ( .A(n926), .B(n925), .CI(n924), .CO(n959), .S(n928) );
  FA_X1 U1006 ( .A(n929), .B(n928), .CI(n927), .CO(n940), .S(n939) );
  OR2_X1 U1007 ( .A1(n941), .A2(n940), .ZN(n1009) );
  NAND2_X1 U1008 ( .A1(n1066), .A2(n1009), .ZN(n944) );
  NOR2_X1 U1009 ( .A1(n1054), .A2(n944), .ZN(n2671) );
  INV_X1 U1010 ( .A(n2671), .ZN(n946) );
  NOR2_X1 U1011 ( .A1(n2672), .A2(n946), .ZN(n973) );
  INV_X1 U1012 ( .A(n973), .ZN(n948) );
  NAND2_X1 U1013 ( .A1(n931), .A2(n930), .ZN(n1068) );
  INV_X1 U1014 ( .A(n1068), .ZN(n935) );
  NAND2_X1 U1015 ( .A1(n933), .A2(n932), .ZN(n1072) );
  INV_X1 U1016 ( .A(n1072), .ZN(n934) );
  AOI21_X1 U1017 ( .B1(n1073), .B2(n935), .A(n934), .ZN(n2692) );
  NAND2_X1 U1018 ( .A1(n937), .A2(n936), .ZN(n1055) );
  NAND2_X1 U1019 ( .A1(n939), .A2(n938), .ZN(n1065) );
  INV_X1 U1020 ( .A(n1065), .ZN(n1003) );
  NAND2_X1 U1021 ( .A1(n941), .A2(n940), .ZN(n1008) );
  INV_X1 U1022 ( .A(n1008), .ZN(n942) );
  AOI21_X1 U1023 ( .B1(n1003), .B2(n1009), .A(n942), .ZN(n943) );
  OAI21_X1 U1024 ( .B1(n944), .B2(n1055), .A(n943), .ZN(n2689) );
  INV_X1 U1025 ( .A(n2689), .ZN(n945) );
  OAI21_X1 U1026 ( .B1(n2692), .B2(n946), .A(n945), .ZN(n976) );
  INV_X1 U1027 ( .A(n976), .ZN(n947) );
  OAI21_X1 U1028 ( .B1(n1049), .B2(n948), .A(n947), .ZN(n968) );
  XNOR2_X1 U1029 ( .A(n2673), .B(n70), .ZN(n990) );
  OAI22_X1 U1030 ( .A1(n990), .A2(n6115), .B1(n991), .B2(n950), .ZN(n984) );
  NOR2_X1 U1031 ( .A1(n952), .A2(n951), .ZN(n989) );
  INV_X1 U1032 ( .A(op_c_i[30]), .ZN(n988) );
  FA_X1 U1033 ( .A(op_c_i[28]), .B(op_c_i[29]), .CI(n953), .CO(n987), .S(n957)
         );
  INV_X1 U1034 ( .A(n954), .ZN(n955) );
  NOR2_X1 U1035 ( .A1(n955), .A2(n2675), .ZN(n982) );
  FA_X1 U1036 ( .A(n958), .B(n957), .CI(n956), .CO(n995), .S(n963) );
  FA_X1 U1037 ( .A(n961), .B(n960), .CI(n959), .CO(n994), .S(n962) );
  FA_X1 U1038 ( .A(n964), .B(n963), .CI(n962), .CO(n965), .S(n941) );
  NOR2_X1 U1039 ( .A1(n966), .A2(n965), .ZN(n2670) );
  INV_X1 U1040 ( .A(n2670), .ZN(n975) );
  NAND2_X1 U1041 ( .A1(n966), .A2(n965), .ZN(n2685) );
  NAND2_X1 U1042 ( .A1(n975), .A2(n2685), .ZN(n967) );
  XNOR2_X1 U1043 ( .A(n968), .B(n967), .ZN(n4963) );
  NAND2_X1 U1044 ( .A1(n2713), .A2(imm_i[0]), .ZN(n1037) );
  INV_X1 U1045 ( .A(n1037), .ZN(n970) );
  NAND2_X1 U1046 ( .A1(n2713), .A2(imm_i[1]), .ZN(n4965) );
  NAND2_X1 U1047 ( .A1(n970), .A2(n4965), .ZN(n5327) );
  NAND2_X1 U1048 ( .A1(n4963), .A2(n5304), .ZN(n1014) );
  INV_X1 U1049 ( .A(n4965), .ZN(n972) );
  AND2_X1 U1050 ( .A1(n972), .A2(n1037), .ZN(n5331) );
  NAND2_X1 U1051 ( .A1(n2713), .A2(short_signed_i[0]), .ZN(n971) );
  NAND2_X1 U1052 ( .A1(n971), .A2(n5218), .ZN(n1015) );
  AND2_X1 U1053 ( .A1(n972), .A2(n1015), .ZN(n1001) );
  NAND2_X1 U1054 ( .A1(n973), .A2(n975), .ZN(n978) );
  NOR2_X1 U1055 ( .A1(n2683), .A2(n978), .ZN(n981) );
  INV_X1 U1056 ( .A(n2685), .ZN(n974) );
  AOI21_X1 U1057 ( .B1(n976), .B2(n975), .A(n974), .ZN(n977) );
  OAI21_X1 U1058 ( .B1(n979), .B2(n978), .A(n977), .ZN(n980) );
  AOI21_X1 U1059 ( .B1(n1002), .B2(n981), .A(n980), .ZN(n1000) );
  FA_X1 U1060 ( .A(n984), .B(n983), .CI(n982), .CO(n2682), .S(n996) );
  INV_X1 U1061 ( .A(n985), .ZN(n986) );
  NOR2_X1 U1062 ( .A1(n986), .A2(n2675), .ZN(n2681) );
  FA_X1 U1063 ( .A(n989), .B(n988), .CI(n987), .CO(n2679), .S(n983) );
  AOI21_X1 U1064 ( .B1(n6115), .B2(n991), .A(n990), .ZN(n993) );
  INV_X1 U1065 ( .A(n993), .ZN(n2677) );
  FA_X1 U1066 ( .A(n996), .B(n995), .CI(n994), .CO(n997), .S(n966) );
  NOR2_X1 U1067 ( .A1(n998), .A2(n997), .ZN(n2686) );
  INV_X1 U1068 ( .A(n2686), .ZN(n999) );
  NAND2_X1 U1069 ( .A1(n998), .A2(n997), .ZN(n2684) );
  OAI21_X1 U1070 ( .B1(n5331), .B2(n1001), .A(n4962), .ZN(n1013) );
  NOR2_X1 U1072 ( .A1(n2672), .A2(n1054), .ZN(n1059) );
  NAND2_X1 U1073 ( .A1(n1059), .A2(n1066), .ZN(n1005) );
  NOR2_X1 U1074 ( .A1(n2683), .A2(n1005), .ZN(n1007) );
  OAI21_X1 U1075 ( .B1(n2692), .B2(n1054), .A(n1055), .ZN(n1060) );
  AOI21_X1 U1076 ( .B1(n1060), .B2(n1066), .A(n1003), .ZN(n1004) );
  OAI21_X1 U1077 ( .B1(n979), .B2(n1005), .A(n1004), .ZN(n1006) );
  AOI21_X1 U1078 ( .B1(n2292), .B2(n1007), .A(n1006), .ZN(n1011) );
  NAND2_X1 U1079 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1080 ( .A(n1011), .B(n1010), .Z(n4958) );
  NAND2_X1 U1081 ( .A1(n4965), .A2(n1037), .ZN(n5325) );
  NAND2_X1 U1082 ( .A1(n4958), .A2(n5302), .ZN(n1012) );
  AND3_X1 U1083 ( .A1(n1014), .A2(n1013), .A3(n1012), .ZN(n5794) );
  INV_X1 U1084 ( .A(n2713), .ZN(n5554) );
  NAND2_X1 U1085 ( .A1(n2713), .A2(imm_i[3]), .ZN(n2830) );
  INV_X1 U1086 ( .A(n2830), .ZN(n2288) );
  NAND2_X1 U1087 ( .A1(n2713), .A2(imm_i[2]), .ZN(n2716) );
  AND2_X1 U1088 ( .A1(n2288), .A2(n2716), .ZN(n5264) );
  AOI21_X1 U1089 ( .B1(n2829), .B2(n2288), .A(n5264), .ZN(n2792) );
  INV_X1 U1090 ( .A(n2792), .ZN(n5348) );
  INV_X1 U1091 ( .A(n1016), .ZN(n2290) );
  INV_X1 U1092 ( .A(n2289), .ZN(n1017) );
  AOI21_X1 U1093 ( .B1(n2292), .B2(n2290), .A(n1017), .ZN(n1022) );
  INV_X1 U1094 ( .A(n1018), .ZN(n1020) );
  NAND2_X1 U1095 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1096 ( .A(n1022), .B(n1021), .Z(n5009) );
  INV_X1 U1097 ( .A(n5009), .ZN(n2723) );
  AOI21_X1 U1098 ( .B1(n2292), .B2(n1024), .A(n1026), .ZN(n1023) );
  INV_X1 U1099 ( .A(n1040), .ZN(n1025) );
  INV_X1 U1100 ( .A(n1024), .ZN(n1038) );
  NAND2_X1 U1101 ( .A1(n1025), .A2(n102), .ZN(n1030) );
  NOR2_X1 U1102 ( .A1(n1038), .A2(n1030), .ZN(n1032) );
  INV_X1 U1103 ( .A(n1026), .ZN(n1041) );
  INV_X1 U1104 ( .A(n1039), .ZN(n1028) );
  AOI21_X1 U1105 ( .B1(n1028), .B2(n102), .A(n1027), .ZN(n1029) );
  OAI21_X1 U1106 ( .B1(n1041), .B2(n1030), .A(n1029), .ZN(n1031) );
  AOI21_X1 U1107 ( .B1(n2292), .B2(n1032), .A(n1031), .ZN(n1036) );
  NAND2_X1 U1108 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1109 ( .A(n1036), .B(n1035), .Z(n4976) );
  NOR2_X1 U1110 ( .A1(n4965), .A2(n1037), .ZN(n5311) );
  INV_X1 U1111 ( .A(n5311), .ZN(n5334) );
  INV_X1 U1112 ( .A(n5334), .ZN(n5008) );
  AOI22_X1 U1113 ( .A1(n5304), .A2(n4977), .B1(n4976), .B2(n5008), .ZN(n1048)
         );
  NOR2_X1 U1114 ( .A1(n1038), .A2(n1040), .ZN(n1043) );
  OAI21_X1 U1115 ( .B1(n1041), .B2(n1040), .A(n1039), .ZN(n1042) );
  AOI21_X1 U1116 ( .B1(n2292), .B2(n1043), .A(n1042), .ZN(n1046) );
  NAND2_X1 U1117 ( .A1(n102), .A2(n1044), .ZN(n1045) );
  XOR2_X1 U1118 ( .A(n1046), .B(n1045), .Z(n4975) );
  NAND2_X1 U1119 ( .A1(n4975), .A2(n5331), .ZN(n1047) );
  OAI211_X1 U1120 ( .C1(n5325), .C2(n2723), .A(n1048), .B(n1047), .ZN(n5512)
         );
  AND2_X1 U1121 ( .A1(n2716), .A2(n2830), .ZN(n5384) );
  INV_X1 U1122 ( .A(n5384), .ZN(n5344) );
  INV_X1 U1123 ( .A(n1049), .ZN(n5221) );
  NAND2_X1 U1124 ( .A1(n1050), .A2(n1068), .ZN(n1051) );
  XNOR2_X1 U1125 ( .A(n5221), .B(n1051), .ZN(n4974) );
  NOR2_X1 U1126 ( .A1(n2683), .A2(n2672), .ZN(n1053) );
  OAI21_X1 U1127 ( .B1(n979), .B2(n2672), .A(n2692), .ZN(n1052) );
  AOI21_X1 U1128 ( .B1(n2292), .B2(n1053), .A(n1052), .ZN(n1058) );
  INV_X1 U1129 ( .A(n1054), .ZN(n1056) );
  NAND2_X1 U1130 ( .A1(n1056), .A2(n1055), .ZN(n1057) );
  XOR2_X1 U1131 ( .A(n1058), .B(n1057), .Z(n4959) );
  AOI22_X1 U1132 ( .A1(n4974), .A2(n5302), .B1(n4959), .B2(n5331), .ZN(n1076)
         );
  INV_X1 U1133 ( .A(n1059), .ZN(n1062) );
  NOR2_X1 U1134 ( .A1(n2683), .A2(n1062), .ZN(n1064) );
  INV_X1 U1135 ( .A(n1060), .ZN(n1061) );
  OAI21_X1 U1136 ( .B1(n979), .B2(n1062), .A(n1061), .ZN(n1063) );
  NOR2_X1 U1137 ( .A1(n2683), .A2(n1069), .ZN(n1071) );
  OAI21_X1 U1138 ( .B1(n979), .B2(n1069), .A(n1068), .ZN(n1070) );
  AOI21_X1 U1139 ( .B1(n2292), .B2(n1071), .A(n1070), .ZN(n1074) );
  AOI22_X1 U1140 ( .A1(n4956), .A2(n5008), .B1(n4957), .B2(n5304), .ZN(n1075)
         );
  AND2_X1 U1141 ( .A1(n1076), .A2(n1075), .ZN(n4894) );
  OR2_X1 U1142 ( .A1(n2288), .A2(n2716), .ZN(n5386) );
  INV_X1 U1143 ( .A(n5386), .ZN(n5257) );
  NAND2_X1 U1144 ( .A1(n4894), .A2(n5257), .ZN(n1077) );
  OAI21_X1 U1145 ( .B1(n5512), .B2(n5344), .A(n1077), .ZN(n1078) );
  NOR2_X1 U1146 ( .A1(n2792), .A2(n2716), .ZN(n5346) );
  AND2_X1 U1147 ( .A1(n6108), .A2(mulh_CS[0]), .ZN(n5215) );
  AOI21_X1 U1148 ( .B1(n2713), .B2(imm_i[4]), .A(n5215), .ZN(n2287) );
  INV_X1 U1149 ( .A(n2287), .ZN(n1079) );
  NAND2_X1 U1150 ( .A1(operator_i[2]), .A2(operator_i[0]), .ZN(n2284) );
  AND2_X1 U1151 ( .A1(n2284), .A2(operator_i[1]), .ZN(n2286) );
  AND2_X1 U1152 ( .A1(n1079), .A2(n2286), .ZN(n5427) );
  INV_X1 U1153 ( .A(clpx_shift_i[1]), .ZN(n1080) );
  NOR2_X1 U1154 ( .A1(n1080), .A2(clpx_shift_i[0]), .ZN(n5463) );
  INV_X1 U1155 ( .A(n23), .ZN(n1116) );
  XNOR2_X1 U1156 ( .A(n1116), .B(dot_op_a_i[24]), .ZN(n1081) );
  XNOR2_X1 U1157 ( .A(n1116), .B(dot_op_a_i[25]), .ZN(n1128) );
  XOR2_X1 U1158 ( .A(n1081), .B(n1128), .Z(n1082) );
  XNOR2_X1 U1159 ( .A(n1116), .B(dot_op_a_i[23]), .ZN(n1098) );
  NAND2_X1 U1160 ( .A1(n1082), .A2(n4660), .ZN(n4661) );
  MUX2_X1 U1161 ( .A(dot_op_b_i[21]), .B(dot_op_b_i[5]), .S(n1087), .Z(n2109)
         );
  XNOR2_X1 U1162 ( .A(n2109), .B(n4587), .ZN(n1129) );
  MUX2_X1 U1163 ( .A(dot_op_b_i[22]), .B(dot_op_b_i[6]), .S(n1123), .Z(n2153)
         );
  XNOR2_X1 U1164 ( .A(n2153), .B(n4587), .ZN(n1289) );
  OAI22_X1 U1165 ( .A1(n4661), .A2(n1129), .B1(n4660), .B2(n1289), .ZN(n1107)
         );
  XNOR2_X1 U1166 ( .A(n1131), .B(dot_op_a_i[18]), .ZN(n1083) );
  XOR2_X1 U1167 ( .A(n1083), .B(n1916), .Z(n1084) );
  XNOR2_X1 U1168 ( .A(n12), .B(dot_op_a_i[17]), .ZN(n1095) );
  MUX2_X1 U1170 ( .A(dot_op_b_i[27]), .B(dot_op_b_i[11]), .S(n1087), .Z(n4740)
         );
  XNOR2_X1 U1171 ( .A(n4740), .B(n69), .ZN(n1160) );
  MUX2_X1 U1172 ( .A(dot_op_b_i[28]), .B(dot_op_b_i[12]), .S(n1123), .Z(n4780)
         );
  XNOR2_X1 U1173 ( .A(n4780), .B(n69), .ZN(n1287) );
  OAI22_X1 U1174 ( .A1(n1931), .A2(n1160), .B1(n6122), .B2(n1287), .ZN(n1106)
         );
  XNOR2_X1 U1175 ( .A(n1116), .B(dot_op_a_i[27]), .ZN(n1117) );
  XNOR2_X1 U1176 ( .A(n1116), .B(dot_op_a_i[26]), .ZN(n1085) );
  XOR2_X1 U1177 ( .A(n4683), .B(n1085), .Z(n1086) );
  MUX2_X1 U1179 ( .A(dot_op_b_i[19]), .B(dot_op_b_i[3]), .S(n1123), .Z(n1819)
         );
  XNOR2_X1 U1180 ( .A(n4683), .B(n1819), .ZN(n1134) );
  MUX2_X1 U1181 ( .A(dot_op_b_i[20]), .B(dot_op_b_i[4]), .S(n1087), .Z(n1784)
         );
  XNOR2_X1 U1182 ( .A(n4683), .B(n1784), .ZN(n1138) );
  OAI22_X1 U1183 ( .A1(n4732), .A2(n1134), .B1(n1138), .B2(n4731), .ZN(n1105)
         );
  INV_X1 U1185 ( .A(n5123), .ZN(n1088) );
  AND2_X1 U1186 ( .A1(n1093), .A2(n1088), .ZN(n1104) );
  INV_X1 U1187 ( .A(dot_op_b_i[30]), .ZN(n1090) );
  INV_X1 U1188 ( .A(dot_op_c_i[14]), .ZN(n3195) );
  OAI22_X1 U1189 ( .A1(n1131), .A2(n1090), .B1(n1661), .B2(n3195), .ZN(n1103)
         );
  INV_X1 U1190 ( .A(dot_op_b_i[31]), .ZN(n2925) );
  INV_X1 U1191 ( .A(dot_op_c_i[15]), .ZN(n3076) );
  OAI22_X1 U1192 ( .A1(n1131), .A2(n2925), .B1(n1661), .B2(n3076), .ZN(n1423)
         );
  OR2_X1 U1193 ( .A1(n1093), .A2(n2848), .ZN(n1092) );
  XOR2_X1 U1194 ( .A(dot_op_a_i[14]), .B(dot_op_a_i[15]), .Z(n1091) );
  NAND2_X1 U1195 ( .A1(n1091), .A2(n5123), .ZN(n5124) );
  OAI22_X1 U1196 ( .A1(n1092), .A2(n5123), .B1(n5124), .B2(n2848), .ZN(n1422)
         );
  MUX2_X1 U1197 ( .A(dot_op_b_i[1]), .B(dot_op_b_i[17]), .S(n1087), .Z(n1812)
         );
  XNOR2_X1 U1198 ( .A(n1812), .B(n1803), .ZN(n1402) );
  XNOR2_X1 U1199 ( .A(n1093), .B(n1803), .ZN(n1094) );
  OAI22_X1 U1200 ( .A1(n1402), .A2(n5123), .B1(n1094), .B2(n5124), .ZN(n1421)
         );
  MUX2_X1 U1201 ( .A(dot_op_b_i[14]), .B(dot_op_b_i[30]), .S(n1123), .Z(n5076)
         );
  INV_X1 U1202 ( .A(dot_op_a_i[1]), .ZN(n1628) );
  XNOR2_X1 U1203 ( .A(n5076), .B(n1612), .ZN(n1127) );
  MUX2_X1 U1204 ( .A(dot_op_b_i[15]), .B(dot_op_b_i[31]), .S(n1123), .Z(n5115)
         );
  XNOR2_X1 U1205 ( .A(n5115), .B(n1612), .ZN(n1408) );
  OAI22_X1 U1206 ( .A1(n1127), .A2(n1778), .B1(n1408), .B2(n1777), .ZN(n1420)
         );
  XNOR2_X1 U1207 ( .A(n1131), .B(dot_op_a_i[16]), .ZN(n1663) );
  INV_X1 U1208 ( .A(n1663), .ZN(n1889) );
  NAND2_X1 U1209 ( .A1(n16), .A2(n1889), .ZN(n1890) );
  MUX2_X1 U1210 ( .A(dot_op_b_i[30]), .B(dot_op_b_i[14]), .S(n1087), .Z(n5078)
         );
  XNOR2_X1 U1211 ( .A(n5078), .B(n16), .ZN(n1101) );
  MUX2_X1 U1212 ( .A(dot_op_b_i[31]), .B(dot_op_b_i[15]), .S(n1087), .Z(n5107)
         );
  XNOR2_X1 U1213 ( .A(n5107), .B(n16), .ZN(n1414) );
  OAI22_X1 U1214 ( .A1(n1890), .A2(n1101), .B1(n1414), .B2(n1889), .ZN(n1419)
         );
  MUX2_X1 U1215 ( .A(dot_op_b_i[5]), .B(dot_op_b_i[21]), .S(n1123), .Z(n2103)
         );
  INV_X1 U1216 ( .A(dot_op_a_i[9]), .ZN(n1313) );
  XNOR2_X1 U1217 ( .A(n2103), .B(n1307), .ZN(n1207) );
  XOR2_X1 U1218 ( .A(dot_op_a_i[8]), .B(dot_op_a_i[9]), .Z(n1096) );
  NAND2_X1 U1219 ( .A1(n1096), .A2(n4629), .ZN(n4630) );
  MUX2_X1 U1220 ( .A(dot_op_b_i[6]), .B(dot_op_b_i[22]), .S(n1087), .Z(n2169)
         );
  XNOR2_X1 U1221 ( .A(n2169), .B(n1307), .ZN(n1110) );
  OAI22_X1 U1222 ( .A1(n1207), .A2(n4630), .B1(n1110), .B2(n4629), .ZN(n1151)
         );
  MUX2_X1 U1223 ( .A(dot_op_b_i[11]), .B(dot_op_b_i[27]), .S(n1123), .Z(n4742)
         );
  XNOR2_X1 U1224 ( .A(n4742), .B(n1808), .ZN(n1158) );
  XOR2_X1 U1225 ( .A(dot_op_a_i[2]), .B(dot_op_a_i[3]), .Z(n1097) );
  NAND2_X1 U1226 ( .A1(n1097), .A2(n1903), .ZN(n1901) );
  MUX2_X1 U1227 ( .A(dot_op_b_i[12]), .B(dot_op_b_i[28]), .S(n1087), .Z(n4795)
         );
  XNOR2_X1 U1228 ( .A(n4795), .B(n1808), .ZN(n1108) );
  OAI22_X1 U1229 ( .A1(n1158), .A2(n1901), .B1(n1108), .B2(n1903), .ZN(n1150)
         );
  XNOR2_X1 U1230 ( .A(n1131), .B(dot_op_a_i[21]), .ZN(n1130) );
  XNOR2_X1 U1231 ( .A(n12), .B(dot_op_a_i[22]), .ZN(n1099) );
  MUX2_X1 U1235 ( .A(dot_op_b_i[23]), .B(dot_op_b_i[7]), .S(n1087), .Z(n2226)
         );
  XNOR2_X1 U1236 ( .A(n2226), .B(n2147), .ZN(n1203) );
  MUX2_X1 U1237 ( .A(dot_op_b_i[24]), .B(dot_op_b_i[8]), .S(n1087), .Z(n4590)
         );
  XNOR2_X1 U1238 ( .A(n4590), .B(n2147), .ZN(n1124) );
  OAI22_X1 U1239 ( .A1(n6130), .A2(n1203), .B1(n6128), .B2(n1124), .ZN(n1149)
         );
  MUX2_X1 U1240 ( .A(dot_op_b_i[29]), .B(dot_op_b_i[13]), .S(n1087), .Z(n4841)
         );
  XNOR2_X1 U1241 ( .A(n4841), .B(n16), .ZN(n1241) );
  OAI22_X1 U1242 ( .A1(n1890), .A2(n1241), .B1(n1101), .B2(n1889), .ZN(n1145)
         );
  MUX2_X1 U1243 ( .A(dot_op_b_i[9]), .B(dot_op_b_i[25]), .S(n1087), .Z(n4655)
         );
  XNOR2_X1 U1244 ( .A(n4655), .B(n1785), .ZN(n1159) );
  XOR2_X1 U1245 ( .A(dot_op_a_i[5]), .B(dot_op_a_i[4]), .Z(n1102) );
  NAND2_X1 U1246 ( .A1(n1102), .A2(n2079), .ZN(n2080) );
  MUX2_X1 U1247 ( .A(dot_op_b_i[10]), .B(dot_op_b_i[26]), .S(n1087), .Z(n4673)
         );
  XNOR2_X1 U1248 ( .A(n4673), .B(n1785), .ZN(n1288) );
  OAI22_X1 U1249 ( .A1(n1159), .A2(n2080), .B1(n1288), .B2(n2079), .ZN(n1144)
         );
  HA_X1 U1250 ( .A(n1104), .B(n1103), .CO(n1424), .S(n1143) );
  FA_X1 U1251 ( .A(n1107), .B(n1106), .CI(n1105), .CO(n1388), .S(n1152) );
  MUX2_X1 U1252 ( .A(dot_op_b_i[13]), .B(dot_op_b_i[29]), .S(n1123), .Z(n4839)
         );
  XNOR2_X1 U1253 ( .A(n4839), .B(n1808), .ZN(n1396) );
  OAI22_X1 U1254 ( .A1(n1108), .A2(n1901), .B1(n1396), .B2(n1903), .ZN(n1430)
         );
  MUX2_X1 U1255 ( .A(dot_op_b_i[4]), .B(dot_op_b_i[20]), .S(n1087), .Z(n1804)
         );
  XNOR2_X1 U1256 ( .A(n1804), .B(n4679), .ZN(n1135) );
  XOR2_X1 U1257 ( .A(dot_op_a_i[11]), .B(dot_op_a_i[10]), .Z(n1109) );
  NAND2_X1 U1258 ( .A1(n1109), .A2(n4745), .ZN(n4746) );
  XNOR2_X1 U1259 ( .A(n2103), .B(n4679), .ZN(n1401) );
  OAI22_X1 U1260 ( .A1(n1135), .A2(n4746), .B1(n1401), .B2(n4745), .ZN(n1429)
         );
  MUX2_X1 U1261 ( .A(dot_op_b_i[7]), .B(dot_op_b_i[23]), .S(n1087), .Z(n2214)
         );
  XNOR2_X1 U1262 ( .A(n2214), .B(n1307), .ZN(n1395) );
  OAI22_X1 U1263 ( .A1(n1110), .A2(n4630), .B1(n1395), .B2(n4629), .ZN(n1428)
         );
  XNOR2_X1 U1264 ( .A(n12), .B(dot_op_a_i[30]), .ZN(n1111) );
  XNOR2_X1 U1265 ( .A(n12), .B(dot_op_a_i[31]), .ZN(n1113) );
  XOR2_X1 U1266 ( .A(n1111), .B(n17), .Z(n1112) );
  XNOR2_X1 U1267 ( .A(n1126), .B(n17), .ZN(n1114) );
  MUX2_X1 U1268 ( .A(dot_op_b_i[17]), .B(dot_op_b_i[1]), .S(n1087), .Z(n1781)
         );
  XNOR2_X1 U1269 ( .A(n1781), .B(n17), .ZN(n1400) );
  OAI22_X1 U1270 ( .A1(n5113), .A2(n1114), .B1(n1400), .B2(n6114), .ZN(n1427)
         );
  MUX2_X1 U1271 ( .A(dot_op_b_i[8]), .B(dot_op_b_i[24]), .S(n1123), .Z(n4592)
         );
  XNOR2_X1 U1272 ( .A(n4592), .B(n28), .ZN(n1136) );
  XOR2_X1 U1273 ( .A(n28), .B(dot_op_a_i[6]), .Z(n1115) );
  NAND2_X1 U1274 ( .A1(n2246), .A2(n1115), .ZN(n2247) );
  XNOR2_X1 U1275 ( .A(n4655), .B(n28), .ZN(n1411) );
  OAI22_X1 U1276 ( .A1(n1136), .A2(n2247), .B1(n1411), .B2(n2246), .ZN(n1426)
         );
  XNOR2_X1 U1277 ( .A(n1116), .B(dot_op_a_i[28]), .ZN(n1118) );
  MUX2_X1 U1279 ( .A(dot_op_b_i[18]), .B(dot_op_b_i[2]), .S(n1087), .Z(n1905)
         );
  XNOR2_X1 U1280 ( .A(n1905), .B(n6111), .ZN(n1137) );
  XNOR2_X1 U1281 ( .A(n1819), .B(n6111), .ZN(n1403) );
  OAI22_X1 U1282 ( .A1(n6125), .A2(n1137), .B1(n6123), .B2(n1403), .ZN(n1425)
         );
  INV_X1 U1283 ( .A(n17), .ZN(n1121) );
  OR2_X1 U1284 ( .A1(n1126), .A2(n1121), .ZN(n1120) );
  OAI22_X1 U1285 ( .A1(n5113), .A2(n1121), .B1(n1120), .B2(n6114), .ZN(n1433)
         );
  MUX2_X1 U1286 ( .A(dot_op_b_i[2]), .B(dot_op_b_i[18]), .S(n1123), .Z(n1770)
         );
  XNOR2_X1 U1287 ( .A(n1770), .B(n30), .ZN(n1125) );
  XOR2_X1 U1288 ( .A(n30), .B(dot_op_a_i[12]), .Z(n1122) );
  NAND2_X1 U1289 ( .A1(n4829), .A2(n1122), .ZN(n4830) );
  MUX2_X1 U1290 ( .A(dot_op_b_i[3]), .B(dot_op_b_i[19]), .S(n1087), .Z(n1825)
         );
  XNOR2_X1 U1291 ( .A(n1825), .B(n30), .ZN(n1398) );
  OAI22_X1 U1292 ( .A1(n1125), .A2(n4830), .B1(n1398), .B2(n4829), .ZN(n1432)
         );
  MUX2_X1 U1293 ( .A(dot_op_b_i[25]), .B(dot_op_b_i[9]), .S(n1123), .Z(n4657)
         );
  XNOR2_X1 U1294 ( .A(n4657), .B(n2147), .ZN(n1397) );
  OAI22_X1 U1295 ( .A1(n6131), .A2(n1124), .B1(n6128), .B2(n1397), .ZN(n1431)
         );
  XNOR2_X1 U1296 ( .A(n1812), .B(n30), .ZN(n1244) );
  OAI22_X1 U1297 ( .A1(n1125), .A2(n4829), .B1(n1244), .B2(n4830), .ZN(n1142)
         );
  AND2_X1 U1298 ( .A1(n1126), .A2(n89), .ZN(n1141) );
  XNOR2_X1 U1299 ( .A(n4839), .B(n1612), .ZN(n1201) );
  OAI22_X1 U1300 ( .A1(n1201), .A2(n1778), .B1(n1127), .B2(n1777), .ZN(n1140)
         );
  XNOR2_X1 U1301 ( .A(n1784), .B(n4587), .ZN(n1222) );
  OAI22_X1 U1302 ( .A1(n4661), .A2(n1222), .B1(n4660), .B2(n1129), .ZN(n1157)
         );
  XNOR2_X1 U1303 ( .A(n1131), .B(dot_op_a_i[20]), .ZN(n1132) );
  XOR2_X1 U1304 ( .A(n1130), .B(n1132), .Z(n1133) );
  XNOR2_X1 U1305 ( .A(n58), .B(n4590), .ZN(n1186) );
  XNOR2_X1 U1306 ( .A(n58), .B(n4657), .ZN(n1253) );
  OAI22_X1 U1307 ( .A1(n2113), .A2(n1186), .B1(n1253), .B2(n50), .ZN(n1156) );
  XNOR2_X1 U1308 ( .A(n4683), .B(n1905), .ZN(n1220) );
  OAI22_X1 U1309 ( .A1(n4732), .A2(n1220), .B1(n1134), .B2(n4731), .ZN(n1155)
         );
  XNOR2_X1 U1310 ( .A(n1825), .B(n4679), .ZN(n1199) );
  OAI22_X1 U1311 ( .A1(n1199), .A2(n4746), .B1(n1135), .B2(n4745), .ZN(n1148)
         );
  XNOR2_X1 U1312 ( .A(n2214), .B(n28), .ZN(n1205) );
  OAI22_X1 U1313 ( .A1(n1205), .A2(n2247), .B1(n1136), .B2(n2246), .ZN(n1147)
         );
  XNOR2_X1 U1314 ( .A(n1781), .B(n6111), .ZN(n1209) );
  OAI22_X1 U1315 ( .A1(n4845), .A2(n1209), .B1(n6123), .B2(n1137), .ZN(n1146)
         );
  XNOR2_X1 U1316 ( .A(n4683), .B(n2109), .ZN(n1409) );
  OAI22_X1 U1317 ( .A1(n4732), .A2(n1138), .B1(n1409), .B2(n4731), .ZN(n1385)
         );
  MUX2_X1 U1318 ( .A(dot_op_b_i[26]), .B(dot_op_b_i[10]), .S(n1087), .Z(n4681)
         );
  XNOR2_X1 U1319 ( .A(n58), .B(n4681), .ZN(n1252) );
  XNOR2_X1 U1320 ( .A(n58), .B(n4740), .ZN(n1415) );
  OAI22_X1 U1321 ( .A1(n2113), .A2(n1252), .B1(n1415), .B2(n50), .ZN(n1384) );
  FA_X1 U1322 ( .A(n1142), .B(n1141), .CI(n1140), .CO(n1383), .S(n1230) );
  FA_X1 U1323 ( .A(n1145), .B(n1144), .CI(n1143), .CO(n1382), .S(n1153) );
  FA_X1 U1324 ( .A(n1148), .B(n1147), .CI(n1146), .CO(n1381), .S(n1228) );
  FA_X1 U1325 ( .A(n1151), .B(n1150), .CI(n1149), .CO(n1380), .S(n1154) );
  FA_X1 U1326 ( .A(n1154), .B(n1153), .CI(n1152), .CO(n1393), .S(n1338) );
  FA_X1 U1327 ( .A(n1157), .B(n1156), .CI(n1155), .CO(n1229), .S(n1332) );
  XNOR2_X1 U1328 ( .A(n4673), .B(n1808), .ZN(n1184) );
  OAI22_X1 U1329 ( .A1(n1184), .A2(n1901), .B1(n1158), .B2(n1903), .ZN(n1213)
         );
  XNOR2_X1 U1330 ( .A(n4592), .B(n1785), .ZN(n1169) );
  OAI22_X1 U1331 ( .A1(n1169), .A2(n2080), .B1(n1159), .B2(n2079), .ZN(n1212)
         );
  XNOR2_X1 U1332 ( .A(n4681), .B(n69), .ZN(n1182) );
  OAI22_X1 U1333 ( .A1(n1931), .A2(n1182), .B1(n6122), .B2(n1160), .ZN(n1211)
         );
  XNOR2_X1 U1334 ( .A(n1804), .B(n28), .ZN(n1266) );
  XNOR2_X1 U1335 ( .A(n2103), .B(n28), .ZN(n1162) );
  OAI22_X1 U1336 ( .A1(n1266), .A2(n2247), .B1(n1162), .B2(n2246), .ZN(n1277)
         );
  XNOR2_X1 U1337 ( .A(n4673), .B(n1612), .ZN(n1194) );
  XNOR2_X1 U1338 ( .A(n4742), .B(n1612), .ZN(n1163) );
  OAI22_X1 U1339 ( .A1(n1194), .A2(n1778), .B1(n1163), .B2(n1777), .ZN(n1276)
         );
  XNOR2_X1 U1340 ( .A(n1770), .B(n1307), .ZN(n1192) );
  XNOR2_X1 U1341 ( .A(n1825), .B(n1307), .ZN(n1171) );
  OAI22_X1 U1342 ( .A1(n1192), .A2(n4630), .B1(n1171), .B2(n4629), .ZN(n1275)
         );
  XNOR2_X1 U1343 ( .A(n4681), .B(n16), .ZN(n1195) );
  XNOR2_X1 U1344 ( .A(n4740), .B(n16), .ZN(n1165) );
  OAI22_X1 U1345 ( .A1(n1890), .A2(n1195), .B1(n1165), .B2(n1889), .ZN(n1280)
         );
  XNOR2_X1 U1346 ( .A(n1812), .B(n4679), .ZN(n1166) );
  XNOR2_X1 U1347 ( .A(n1093), .B(n4679), .ZN(n1161) );
  OAI22_X1 U1348 ( .A1(n1166), .A2(n4745), .B1(n1161), .B2(n4746), .ZN(n1279)
         );
  XNOR2_X1 U1349 ( .A(n1784), .B(n2147), .ZN(n1268) );
  XNOR2_X1 U1350 ( .A(n2109), .B(n2147), .ZN(n1172) );
  OAI22_X1 U1351 ( .A1(n6131), .A2(n1268), .B1(n6128), .B2(n1172), .ZN(n1278)
         );
  XNOR2_X1 U1352 ( .A(n2169), .B(n1785), .ZN(n1267) );
  XNOR2_X1 U1353 ( .A(n2214), .B(n1785), .ZN(n1170) );
  OAI22_X1 U1354 ( .A1(n1267), .A2(n2080), .B1(n1170), .B2(n2079), .ZN(n1283)
         );
  XNOR2_X1 U1355 ( .A(n4592), .B(n1808), .ZN(n1196) );
  XNOR2_X1 U1356 ( .A(n4655), .B(n1808), .ZN(n1185) );
  OAI22_X1 U1357 ( .A1(n1196), .A2(n1901), .B1(n1185), .B2(n1903), .ZN(n1282)
         );
  XNOR2_X1 U1358 ( .A(n4590), .B(n69), .ZN(n1270) );
  XNOR2_X1 U1359 ( .A(n4657), .B(n69), .ZN(n1183) );
  OAI22_X1 U1360 ( .A1(n1931), .A2(n1270), .B1(n6122), .B2(n1183), .ZN(n1281)
         );
  XNOR2_X1 U1361 ( .A(n2169), .B(n28), .ZN(n1206) );
  OAI22_X1 U1362 ( .A1(n1162), .A2(n2247), .B1(n1206), .B2(n2246), .ZN(n1191)
         );
  XNOR2_X1 U1363 ( .A(n4795), .B(dot_op_a_i[1]), .ZN(n1202) );
  OAI22_X1 U1364 ( .A1(n1163), .A2(n1778), .B1(n1202), .B2(n1777), .ZN(n1190)
         );
  INV_X1 U1365 ( .A(n4844), .ZN(n1164) );
  AND2_X1 U1366 ( .A1(n1126), .A2(n1164), .ZN(n1189) );
  XNOR2_X1 U1367 ( .A(n4780), .B(n16), .ZN(n1242) );
  OAI22_X1 U1368 ( .A1(n1890), .A2(n1165), .B1(n1242), .B2(n1889), .ZN(n1175)
         );
  XNOR2_X1 U1369 ( .A(n1770), .B(n4679), .ZN(n1200) );
  OAI22_X1 U1370 ( .A1(n1200), .A2(n4745), .B1(n1166), .B2(n4746), .ZN(n1174)
         );
  INV_X1 U1371 ( .A(n4829), .ZN(n1167) );
  AND2_X1 U1372 ( .A1(n1093), .A2(n1167), .ZN(n1238) );
  INV_X1 U1373 ( .A(dot_op_b_i[28]), .ZN(n1168) );
  INV_X1 U1374 ( .A(dot_op_c_i[12]), .ZN(n3662) );
  OAI22_X1 U1375 ( .A1(n1131), .A2(n1168), .B1(n1661), .B2(n3662), .ZN(n1237)
         );
  OAI22_X1 U1376 ( .A1(n1170), .A2(n2080), .B1(n1169), .B2(n2079), .ZN(n1181)
         );
  XNOR2_X1 U1377 ( .A(n1804), .B(n1307), .ZN(n1208) );
  OAI22_X1 U1378 ( .A1(n1171), .A2(n4630), .B1(n1208), .B2(n4629), .ZN(n1180)
         );
  XNOR2_X1 U1379 ( .A(n2153), .B(n2147), .ZN(n1204) );
  OAI22_X1 U1380 ( .A1(n6130), .A2(n1172), .B1(n6128), .B2(n1204), .ZN(n1179)
         );
  FA_X1 U1381 ( .A(n1175), .B(n1174), .CI(n1173), .CO(n1247), .S(n1302) );
  INV_X1 U1382 ( .A(n4683), .ZN(n1177) );
  OR2_X1 U1383 ( .A1(n1126), .A2(n1177), .ZN(n1176) );
  OAI22_X1 U1384 ( .A1(n4732), .A2(n1177), .B1(n1176), .B2(n4731), .ZN(n1320)
         );
  XNOR2_X1 U1385 ( .A(n58), .B(n2153), .ZN(n1271) );
  XNOR2_X1 U1386 ( .A(n58), .B(n2226), .ZN(n1187) );
  OAI22_X1 U1387 ( .A1(n2113), .A2(n1271), .B1(n1187), .B2(n50), .ZN(n1319) );
  XNOR2_X1 U1388 ( .A(n4683), .B(n1126), .ZN(n1178) );
  XNOR2_X1 U1389 ( .A(n4683), .B(n1781), .ZN(n1221) );
  OAI22_X1 U1390 ( .A1(n4732), .A2(n1178), .B1(n1221), .B2(n4731), .ZN(n1318)
         );
  FA_X1 U1391 ( .A(n1181), .B(n1180), .CI(n1179), .CO(n1246), .S(n1300) );
  OAI22_X1 U1392 ( .A1(n1931), .A2(n1183), .B1(n6122), .B2(n1182), .ZN(n1234)
         );
  OAI22_X1 U1393 ( .A1(n1185), .A2(n1901), .B1(n1184), .B2(n1903), .ZN(n1233)
         );
  XNOR2_X1 U1394 ( .A(n1234), .B(n1233), .ZN(n1188) );
  OAI22_X1 U1395 ( .A1(n2113), .A2(n1187), .B1(n1186), .B2(n50), .ZN(n1232) );
  XNOR2_X1 U1396 ( .A(n1188), .B(n1232), .ZN(n1370) );
  FA_X1 U1397 ( .A(n1191), .B(n1190), .CI(n1189), .CO(n1248), .S(n1369) );
  XNOR2_X1 U1398 ( .A(n1812), .B(n1307), .ZN(n1309) );
  OAI22_X1 U1399 ( .A1(n1192), .A2(n4629), .B1(n1309), .B2(n4630), .ZN(n1323)
         );
  INV_X1 U1400 ( .A(n4731), .ZN(n1193) );
  AND2_X1 U1401 ( .A1(n1126), .A2(n1193), .ZN(n1322) );
  XNOR2_X1 U1402 ( .A(n4655), .B(n1612), .ZN(n1316) );
  OAI22_X1 U1403 ( .A1(n1316), .A2(n1778), .B1(n1194), .B2(n1777), .ZN(n1321)
         );
  XNOR2_X1 U1404 ( .A(n1905), .B(n4587), .ZN(n1269) );
  XNOR2_X1 U1405 ( .A(n1819), .B(n4587), .ZN(n1223) );
  OAI22_X1 U1406 ( .A1(n4661), .A2(n1269), .B1(n4660), .B2(n1223), .ZN(n1352)
         );
  XNOR2_X1 U1407 ( .A(n4657), .B(n16), .ZN(n1306) );
  OAI22_X1 U1408 ( .A1(n1890), .A2(n1306), .B1(n1195), .B2(n1889), .ZN(n1359)
         );
  XNOR2_X1 U1409 ( .A(n2214), .B(n1808), .ZN(n1325) );
  OAI22_X1 U1410 ( .A1(n1325), .A2(n1901), .B1(n1196), .B2(n1903), .ZN(n1358)
         );
  INV_X1 U1411 ( .A(n4745), .ZN(n1197) );
  AND2_X1 U1412 ( .A1(n1093), .A2(n1197), .ZN(n1225) );
  INV_X1 U1413 ( .A(dot_op_b_i[26]), .ZN(n1198) );
  INV_X1 U1414 ( .A(dot_op_c_i[10]), .ZN(n3568) );
  OAI22_X1 U1415 ( .A1(n1131), .A2(n1198), .B1(n1661), .B2(n3568), .ZN(n1224)
         );
  OAI22_X1 U1416 ( .A1(n1200), .A2(n4746), .B1(n1199), .B2(n4745), .ZN(n1216)
         );
  OAI22_X1 U1417 ( .A1(n1202), .A2(n1778), .B1(n1201), .B2(n1777), .ZN(n1215)
         );
  OAI22_X1 U1418 ( .A1(n2234), .A2(n1204), .B1(n6128), .B2(n1203), .ZN(n1214)
         );
  OAI22_X1 U1419 ( .A1(n1206), .A2(n2247), .B1(n1205), .B2(n2246), .ZN(n1219)
         );
  OAI22_X1 U1420 ( .A1(n1208), .A2(n4630), .B1(n1207), .B2(n4629), .ZN(n1218)
         );
  XNOR2_X1 U1421 ( .A(n1126), .B(n6111), .ZN(n1210) );
  OAI22_X1 U1422 ( .A1(n4845), .A2(n1210), .B1(n6123), .B2(n1209), .ZN(n1217)
         );
  FA_X1 U1423 ( .A(n1213), .B(n1212), .CI(n1211), .CO(n1290), .S(n1331) );
  FA_X1 U1424 ( .A(n1216), .B(n1215), .CI(n1214), .CO(n1292), .S(n1259) );
  FA_X1 U1425 ( .A(n1219), .B(n1218), .CI(n1217), .CO(n1291), .S(n1258) );
  OAI22_X1 U1426 ( .A1(n4732), .A2(n1221), .B1(n1220), .B2(n4731), .ZN(n1274)
         );
  OAI22_X1 U1427 ( .A1(n4661), .A2(n1223), .B1(n4660), .B2(n1222), .ZN(n1273)
         );
  HA_X1 U1428 ( .A(n1225), .B(n1224), .CO(n1265), .S(n1357) );
  INV_X1 U1429 ( .A(dot_op_b_i[27]), .ZN(n1226) );
  INV_X1 U1430 ( .A(dot_op_c_i[11]), .ZN(n3640) );
  OAI22_X1 U1431 ( .A1(n1131), .A2(n1226), .B1(n1661), .B2(n3640), .ZN(n1264)
         );
  OR2_X1 U1432 ( .A1(n1093), .A2(n3084), .ZN(n1227) );
  OAI22_X1 U1433 ( .A1(n1227), .A2(n4745), .B1(n4746), .B2(n3084), .ZN(n1263)
         );
  FA_X1 U1434 ( .A(n1230), .B(n1229), .CI(n1228), .CO(n1391), .S(n1296) );
  OR2_X1 U1435 ( .A1(n1234), .A2(n1233), .ZN(n1231) );
  NAND2_X1 U1436 ( .A1(n1232), .A2(n1231), .ZN(n1236) );
  NAND2_X1 U1437 ( .A1(n1234), .A2(n1233), .ZN(n1235) );
  NAND2_X1 U1438 ( .A1(n1236), .A2(n1235), .ZN(n1262) );
  HA_X1 U1439 ( .A(n1238), .B(n1237), .CO(n1251), .S(n1173) );
  INV_X1 U1440 ( .A(dot_op_b_i[29]), .ZN(n1239) );
  INV_X1 U1441 ( .A(dot_op_c_i[13]), .ZN(n3300) );
  OAI22_X1 U1442 ( .A1(n1131), .A2(n1239), .B1(n1661), .B2(n3300), .ZN(n1250)
         );
  OR2_X1 U1443 ( .A1(n1093), .A2(n3016), .ZN(n1240) );
  OAI22_X1 U1444 ( .A1(n1240), .A2(n4829), .B1(n4830), .B2(n3016), .ZN(n1249)
         );
  OAI22_X1 U1445 ( .A1(n1890), .A2(n1242), .B1(n1241), .B2(n1889), .ZN(n1256)
         );
  XNOR2_X1 U1446 ( .A(n1093), .B(n30), .ZN(n1243) );
  OAI22_X1 U1447 ( .A1(n1244), .A2(n4829), .B1(n1243), .B2(n4830), .ZN(n1255)
         );
  OR2_X1 U1448 ( .A1(n1126), .A2(n36), .ZN(n1245) );
  OAI22_X1 U1449 ( .A1(n4845), .A2(n36), .B1(n6123), .B2(n1245), .ZN(n1254) );
  FA_X1 U1450 ( .A(n1248), .B(n1247), .CI(n1246), .CO(n1294), .S(n1335) );
  FA_X1 U1451 ( .A(n1251), .B(n1250), .CI(n1249), .CO(n1286), .S(n1261) );
  OAI22_X1 U1452 ( .A1(n2113), .A2(n1253), .B1(n1252), .B2(n50), .ZN(n1285) );
  FA_X1 U1453 ( .A(n1256), .B(n1255), .CI(n1254), .CO(n1284), .S(n1260) );
  FA_X1 U1454 ( .A(n1259), .B(n1258), .CI(n1257), .CO(n1297), .S(n1347) );
  FA_X1 U1455 ( .A(n1262), .B(n1261), .CI(n1260), .CO(n1295), .S(n1346) );
  FA_X1 U1456 ( .A(n1265), .B(n1264), .CI(n1263), .CO(n1272), .S(n1350) );
  XNOR2_X1 U1457 ( .A(n1825), .B(n28), .ZN(n1317) );
  OAI22_X1 U1458 ( .A1(n1317), .A2(n2247), .B1(n1266), .B2(n2246), .ZN(n1329)
         );
  XNOR2_X1 U1459 ( .A(n2103), .B(n1785), .ZN(n1315) );
  OAI22_X1 U1460 ( .A1(n1315), .A2(n2080), .B1(n1267), .B2(n2079), .ZN(n1328)
         );
  XNOR2_X1 U1461 ( .A(n1819), .B(n2147), .ZN(n1310) );
  OAI22_X1 U1462 ( .A1(n2234), .A2(n1310), .B1(n6128), .B2(n1268), .ZN(n1327)
         );
  XNOR2_X1 U1463 ( .A(n1781), .B(n4587), .ZN(n1362) );
  OAI22_X1 U1464 ( .A1(n4661), .A2(n1362), .B1(n4660), .B2(n1269), .ZN(n1356)
         );
  XNOR2_X1 U1465 ( .A(n2226), .B(n69), .ZN(n1324) );
  OAI22_X1 U1466 ( .A1(n1931), .A2(n1324), .B1(n6122), .B2(n1270), .ZN(n1355)
         );
  XNOR2_X1 U1467 ( .A(n58), .B(n2109), .ZN(n1326) );
  OAI22_X1 U1468 ( .A1(n2113), .A2(n1326), .B1(n1271), .B2(n50), .ZN(n1354) );
  FA_X1 U1469 ( .A(n1274), .B(n1273), .CI(n1272), .CO(n1257), .S(n1372) );
  FA_X1 U1470 ( .A(n1277), .B(n1276), .CI(n1275), .CO(n1305), .S(n1499) );
  FA_X1 U1471 ( .A(n1280), .B(n1279), .CI(n1278), .CO(n1304), .S(n1498) );
  FA_X1 U1472 ( .A(n1283), .B(n1282), .CI(n1281), .CO(n1303), .S(n1497) );
  FA_X1 U1473 ( .A(n1286), .B(n1285), .CI(n1284), .CO(n1406), .S(n1293) );
  XNOR2_X1 U1474 ( .A(n4841), .B(n69), .ZN(n1407) );
  OAI22_X1 U1475 ( .A1(n1931), .A2(n1287), .B1(n6122), .B2(n1407), .ZN(n1436)
         );
  XNOR2_X1 U1476 ( .A(n4742), .B(n1785), .ZN(n1410) );
  OAI22_X1 U1477 ( .A1(n1288), .A2(n2080), .B1(n1410), .B2(n2079), .ZN(n1435)
         );
  XNOR2_X1 U1478 ( .A(n2226), .B(n4587), .ZN(n1413) );
  OAI22_X1 U1479 ( .A1(n4661), .A2(n1289), .B1(n4660), .B2(n1413), .ZN(n1434)
         );
  FA_X1 U1480 ( .A(n1292), .B(n1291), .CI(n1290), .CO(n1404), .S(n1298) );
  FA_X1 U1481 ( .A(n1295), .B(n1294), .CI(n1293), .CO(n1438), .S(n1340) );
  FA_X1 U1482 ( .A(n1298), .B(n1297), .CI(n1296), .CO(n1437), .S(n1341) );
  FA_X1 U1483 ( .A(n1302), .B(n1301), .CI(n1300), .CO(n1334), .S(n1737) );
  FA_X1 U1484 ( .A(n1305), .B(n1304), .CI(n1303), .CO(n1330), .S(n1736) );
  XNOR2_X1 U1485 ( .A(n4590), .B(n16), .ZN(n1364) );
  OAI22_X1 U1486 ( .A1(n1890), .A2(n1364), .B1(n1306), .B2(n1889), .ZN(n1493)
         );
  XNOR2_X1 U1487 ( .A(n1093), .B(n1307), .ZN(n1308) );
  OAI22_X1 U1488 ( .A1(n1309), .A2(n4629), .B1(n1308), .B2(n4630), .ZN(n1492)
         );
  XNOR2_X1 U1489 ( .A(n1905), .B(n2147), .ZN(n1483) );
  OAI22_X1 U1490 ( .A1(n6130), .A2(n1483), .B1(n6128), .B2(n1310), .ZN(n1491)
         );
  INV_X1 U1491 ( .A(n4629), .ZN(n1311) );
  AND2_X1 U1492 ( .A1(n1093), .A2(n1311), .ZN(n1367) );
  INV_X1 U1493 ( .A(dot_op_b_i[24]), .ZN(n1312) );
  INV_X1 U1494 ( .A(dot_op_c_i[8]), .ZN(n3821) );
  OAI22_X1 U1495 ( .A1(n1131), .A2(n1312), .B1(n1661), .B2(n3821), .ZN(n1366)
         );
  INV_X1 U1496 ( .A(dot_op_c_i[9]), .ZN(n3692) );
  OAI22_X1 U1497 ( .A1(n1131), .A2(n2623), .B1(n1661), .B2(n3692), .ZN(n1486)
         );
  OR2_X1 U1498 ( .A1(n1093), .A2(n1313), .ZN(n1314) );
  OAI22_X1 U1499 ( .A1(n1314), .A2(n4629), .B1(n4630), .B2(n1313), .ZN(n1485)
         );
  XNOR2_X1 U1500 ( .A(n1804), .B(n1785), .ZN(n1481) );
  OAI22_X1 U1501 ( .A1(n1481), .A2(n2080), .B1(n1315), .B2(n2079), .ZN(n1490)
         );
  XNOR2_X1 U1502 ( .A(n4592), .B(dot_op_a_i[1]), .ZN(n1475) );
  OAI22_X1 U1503 ( .A1(n1475), .A2(n1778), .B1(n1316), .B2(n1777), .ZN(n1489)
         );
  XNOR2_X1 U1504 ( .A(n1770), .B(n28), .ZN(n1365) );
  OAI22_X1 U1505 ( .A1(n1365), .A2(n2247), .B1(n1317), .B2(n2246), .ZN(n1488)
         );
  FA_X1 U1506 ( .A(n1320), .B(n1319), .CI(n1318), .CO(n1301), .S(n1501) );
  FA_X1 U1507 ( .A(n1323), .B(n1322), .CI(n1321), .CO(n1353), .S(n1450) );
  XNOR2_X1 U1508 ( .A(n2153), .B(n69), .ZN(n1477) );
  OAI22_X1 U1509 ( .A1(n1931), .A2(n1477), .B1(n6122), .B2(n1324), .ZN(n1496)
         );
  XNOR2_X1 U1510 ( .A(n2169), .B(n1808), .ZN(n1479) );
  OAI22_X1 U1511 ( .A1(n1479), .A2(n1901), .B1(n1325), .B2(n1903), .ZN(n1495)
         );
  XNOR2_X1 U1512 ( .A(n58), .B(n1784), .ZN(n1459) );
  OAI22_X1 U1513 ( .A1(n2113), .A2(n1459), .B1(n1326), .B2(n50), .ZN(n1494) );
  FA_X1 U1514 ( .A(n1329), .B(n1328), .CI(n1327), .CO(n1349), .S(n1448) );
  FA_X1 U1515 ( .A(n1332), .B(n1331), .CI(n1330), .CO(n1337), .S(n1375) );
  FA_X1 U1516 ( .A(n1335), .B(n1334), .CI(n1333), .CO(n1336), .S(n1374) );
  FA_X1 U1517 ( .A(n1338), .B(n1337), .CI(n1336), .CO(n1377), .S(n1343) );
  FA_X1 U1518 ( .A(n1341), .B(n1340), .CI(n1339), .CO(n1442), .S(n1342) );
  OR2_X1 U1519 ( .A1(n1763), .A2(n1762), .ZN(n5161) );
  FA_X1 U1520 ( .A(n1344), .B(n1343), .CI(n1342), .CO(n1762), .S(n1761) );
  FA_X1 U1521 ( .A(n1347), .B(n1346), .CI(n1345), .CO(n1339), .S(n1734) );
  FA_X1 U1522 ( .A(n1350), .B(n1349), .CI(n1348), .CO(n1373), .S(n1470) );
  FA_X1 U1523 ( .A(n1353), .B(n1352), .CI(n1351), .CO(n1368), .S(n1469) );
  FA_X1 U1524 ( .A(n1356), .B(n1355), .CI(n1354), .CO(n1348), .S(n1447) );
  FA_X1 U1525 ( .A(n1359), .B(n1358), .CI(n1357), .CO(n1351), .S(n1446) );
  INV_X1 U1526 ( .A(n4587), .ZN(n1361) );
  OR2_X1 U1527 ( .A1(n1126), .A2(n1361), .ZN(n1360) );
  OAI22_X1 U1528 ( .A1(n4661), .A2(n1361), .B1(n4660), .B2(n1360), .ZN(n1467)
         );
  XNOR2_X1 U1529 ( .A(n1126), .B(n4587), .ZN(n1363) );
  OAI22_X1 U1530 ( .A1(n4661), .A2(n1363), .B1(n4660), .B2(n1362), .ZN(n1466)
         );
  XNOR2_X1 U1531 ( .A(n2226), .B(n16), .ZN(n1461) );
  OAI22_X1 U1532 ( .A1(n1890), .A2(n1461), .B1(n1364), .B2(n1889), .ZN(n1455)
         );
  XNOR2_X1 U1533 ( .A(n1812), .B(n28), .ZN(n1463) );
  OAI22_X1 U1534 ( .A1(n1365), .A2(n2246), .B1(n1463), .B2(n2247), .ZN(n1454)
         );
  HA_X1 U1535 ( .A(n1367), .B(n1366), .CO(n1487), .S(n1453) );
  FA_X1 U1536 ( .A(n1370), .B(n1369), .CI(n1368), .CO(n1333), .S(n1742) );
  FA_X1 U1537 ( .A(n1373), .B(n1372), .CI(n1371), .CO(n1345), .S(n1741) );
  FA_X1 U1538 ( .A(n1376), .B(n1375), .CI(n1374), .CO(n1344), .S(n1732) );
  NOR2_X1 U1539 ( .A1(n1761), .A2(n1760), .ZN(n5159) );
  INV_X1 U1540 ( .A(n5159), .ZN(n5532) );
  NAND2_X1 U1541 ( .A1(n5161), .A2(n5532), .ZN(n4914) );
  FA_X1 U1542 ( .A(n1379), .B(n1378), .CI(n1377), .CO(n2054), .S(n1440) );
  FA_X1 U1543 ( .A(n1382), .B(n1381), .CI(n1380), .CO(n1960), .S(n1389) );
  FA_X1 U1544 ( .A(n1385), .B(n1384), .CI(n1383), .CO(n1959), .S(n1390) );
  FA_X1 U1545 ( .A(n1388), .B(n1387), .CI(n1386), .CO(n1958), .S(n1394) );
  FA_X1 U1546 ( .A(n1391), .B(n1390), .CI(n1389), .CO(n2029), .S(n1378) );
  FA_X1 U1547 ( .A(n1394), .B(n1393), .CI(n1392), .CO(n2028), .S(n1379) );
  XNOR2_X1 U1548 ( .A(n4592), .B(n1307), .ZN(n1793) );
  OAI22_X1 U1549 ( .A1(n1395), .A2(n4630), .B1(n1793), .B2(n4629), .ZN(n1923)
         );
  XNOR2_X1 U1550 ( .A(n5076), .B(n1808), .ZN(n1809) );
  OAI22_X1 U1551 ( .A1(n1396), .A2(n1901), .B1(n1809), .B2(n1903), .ZN(n1922)
         );
  XNOR2_X1 U1552 ( .A(n4681), .B(n2147), .ZN(n1788) );
  OAI22_X1 U1553 ( .A1(n2234), .A2(n1397), .B1(n6128), .B2(n1788), .ZN(n1921)
         );
  XNOR2_X1 U1554 ( .A(n1804), .B(n30), .ZN(n1790) );
  OAI22_X1 U1555 ( .A1(n1398), .A2(n4830), .B1(n1790), .B2(n4829), .ZN(n1887)
         );
  AND2_X1 U1556 ( .A1(dot_op_a_i[31]), .A2(dot_signed_i[1]), .ZN(n3407) );
  INV_X1 U1557 ( .A(n5109), .ZN(n1399) );
  AND2_X1 U1558 ( .A1(n1126), .A2(n1399), .ZN(n1886) );
  XNOR2_X1 U1559 ( .A(n1905), .B(n17), .ZN(n1817) );
  XNOR2_X1 U1560 ( .A(n2169), .B(n4679), .ZN(n1789) );
  OAI22_X1 U1561 ( .A1(n1401), .A2(n4746), .B1(n1789), .B2(n4745), .ZN(n1894)
         );
  XNOR2_X1 U1562 ( .A(n1770), .B(n1803), .ZN(n1786) );
  OAI22_X1 U1563 ( .A1(n1786), .A2(n5123), .B1(n1402), .B2(n5124), .ZN(n1893)
         );
  XNOR2_X1 U1564 ( .A(n1784), .B(n6111), .ZN(n1792) );
  OAI22_X1 U1565 ( .A1(n4845), .A2(n1403), .B1(n4844), .B2(n1792), .ZN(n1892)
         );
  FA_X1 U1566 ( .A(n1406), .B(n1405), .CI(n1404), .CO(n2011), .S(n1439) );
  XNOR2_X1 U1567 ( .A(n5078), .B(n69), .ZN(n1780) );
  OAI22_X1 U1568 ( .A1(n1931), .A2(n1407), .B1(n6122), .B2(n1780), .ZN(n1926)
         );
  XNOR2_X1 U1569 ( .A(n5085), .B(n1612), .ZN(n1776) );
  OAI22_X1 U1570 ( .A1(n1776), .A2(n1777), .B1(n1408), .B2(n1778), .ZN(n1925)
         );
  XNOR2_X1 U1571 ( .A(n4683), .B(n2153), .ZN(n1783) );
  OAI22_X1 U1572 ( .A1(n4732), .A2(n1409), .B1(n1783), .B2(n4731), .ZN(n1924)
         );
  XNOR2_X1 U1573 ( .A(n4795), .B(n1785), .ZN(n1795) );
  OAI22_X1 U1574 ( .A1(n1410), .A2(n2080), .B1(n1795), .B2(n2079), .ZN(n1920)
         );
  XNOR2_X1 U1575 ( .A(n4673), .B(n28), .ZN(n1787) );
  OAI22_X1 U1576 ( .A1(n1411), .A2(n2247), .B1(n1787), .B2(n2246), .ZN(n1919)
         );
  INV_X1 U1577 ( .A(dot_op_c_i[16]), .ZN(n3029) );
  AND2_X1 U1578 ( .A1(n5107), .A2(dot_signed_i[0]), .ZN(n5083) );
  OAI21_X1 U1579 ( .B1(n1661), .B2(n3029), .A(n5114), .ZN(n1815) );
  AND2_X1 U1580 ( .A1(dot_op_a_i[15]), .A2(dot_signed_i[1]), .ZN(n3312) );
  INV_X1 U1581 ( .A(n5116), .ZN(n1412) );
  AND2_X1 U1582 ( .A1(n1093), .A2(n1412), .ZN(n1814) );
  XNOR2_X1 U1583 ( .A(n4590), .B(n4587), .ZN(n1775) );
  OAI22_X1 U1584 ( .A1(n4661), .A2(n1413), .B1(n4660), .B2(n1775), .ZN(n1847)
         );
  XNOR2_X1 U1585 ( .A(n5083), .B(n16), .ZN(n1888) );
  OAI22_X1 U1586 ( .A1(n1888), .A2(n1889), .B1(n1890), .B2(n1414), .ZN(n1846)
         );
  XNOR2_X1 U1587 ( .A(n58), .B(n4780), .ZN(n1774) );
  OAI22_X1 U1588 ( .A1(n2113), .A2(n1415), .B1(n1774), .B2(n50), .ZN(n1845) );
  FA_X1 U1589 ( .A(n1418), .B(n1417), .CI(n1416), .CO(n2009), .S(n1392) );
  FA_X1 U1590 ( .A(n1421), .B(n1420), .CI(n1419), .CO(n1873), .S(n1386) );
  FA_X1 U1591 ( .A(n1424), .B(n1423), .CI(n1422), .CO(n1872), .S(n1387) );
  FA_X1 U1592 ( .A(n1427), .B(n1426), .CI(n1425), .CO(n1871), .S(n1417) );
  FA_X1 U1593 ( .A(n1430), .B(n1429), .CI(n1428), .CO(n1885), .S(n1418) );
  FA_X1 U1594 ( .A(n1433), .B(n1432), .CI(n1431), .CO(n1884), .S(n1416) );
  FA_X1 U1595 ( .A(n1436), .B(n1435), .CI(n1434), .CO(n1883), .S(n1405) );
  FA_X1 U1596 ( .A(n1439), .B(n1438), .CI(n1437), .CO(n2040), .S(n1441) );
  NAND2_X1 U1597 ( .A1(n1440), .A2(n105), .ZN(n1444) );
  NAND2_X1 U1598 ( .A1(n1442), .A2(n1441), .ZN(n1443) );
  NAND2_X1 U1599 ( .A1(n1444), .A2(n1443), .ZN(n1758) );
  NOR2_X1 U1600 ( .A1(n1759), .A2(n1758), .ZN(n4915) );
  NOR2_X1 U1601 ( .A1(n4914), .A2(n4915), .ZN(n1757) );
  FA_X1 U1602 ( .A(n1447), .B(n1446), .CI(n1445), .CO(n1468), .S(n1530) );
  FA_X1 U1603 ( .A(n1450), .B(n1449), .CI(n1448), .CO(n1500), .S(n1529) );
  XNOR2_X1 U1604 ( .A(n1784), .B(n69), .ZN(n1544) );
  XNOR2_X1 U1605 ( .A(n2109), .B(n69), .ZN(n1478) );
  OAI22_X1 U1606 ( .A1(n1931), .A2(n1544), .B1(n6122), .B2(n1478), .ZN(n1577)
         );
  XNOR2_X1 U1607 ( .A(n1770), .B(n1785), .ZN(n1516) );
  XNOR2_X1 U1608 ( .A(n1825), .B(n1785), .ZN(n1482) );
  OAI22_X1 U1609 ( .A1(n1516), .A2(n2080), .B1(n1482), .B2(n2079), .ZN(n1576)
         );
  XNOR2_X1 U1610 ( .A(n58), .B(n1905), .ZN(n1543) );
  XNOR2_X1 U1611 ( .A(n58), .B(n1819), .ZN(n1460) );
  OAI22_X1 U1612 ( .A1(n2113), .A2(n1543), .B1(n1460), .B2(n50), .ZN(n1575) );
  XNOR2_X1 U1613 ( .A(n1804), .B(n1808), .ZN(n1513) );
  XNOR2_X1 U1614 ( .A(n2103), .B(n1808), .ZN(n1480) );
  OAI22_X1 U1615 ( .A1(n1513), .A2(n1901), .B1(n1480), .B2(n1903), .ZN(n1539)
         );
  XNOR2_X1 U1616 ( .A(n2169), .B(n1612), .ZN(n1512) );
  XNOR2_X1 U1617 ( .A(n2214), .B(dot_op_a_i[1]), .ZN(n1476) );
  OAI22_X1 U1618 ( .A1(n1512), .A2(n1778), .B1(n1476), .B2(n1777), .ZN(n1538)
         );
  INV_X1 U1619 ( .A(n2147), .ZN(n1452) );
  OR2_X1 U1620 ( .A1(n1126), .A2(n1452), .ZN(n1451) );
  OAI22_X1 U1621 ( .A1(n6130), .A2(n1452), .B1(n2233), .B2(n1451), .ZN(n1537)
         );
  FA_X1 U1622 ( .A(n1455), .B(n1454), .CI(n1453), .CO(n1465), .S(n1552) );
  INV_X1 U1623 ( .A(n2246), .ZN(n1456) );
  AND2_X1 U1624 ( .A1(n1093), .A2(n1456), .ZN(n1518) );
  INV_X1 U1625 ( .A(dot_op_b_i[22]), .ZN(n1457) );
  INV_X1 U1626 ( .A(dot_op_c_i[6]), .ZN(n3981) );
  OAI22_X1 U1627 ( .A1(n1131), .A2(n1457), .B1(n1661), .B2(n3981), .ZN(n1517)
         );
  INV_X1 U1628 ( .A(dot_op_b_i[23]), .ZN(n2929) );
  INV_X1 U1629 ( .A(dot_op_c_i[7]), .ZN(n3893) );
  OAI22_X1 U1630 ( .A1(n1131), .A2(n2929), .B1(n1661), .B2(n3893), .ZN(n1520)
         );
  OR2_X1 U1631 ( .A1(n1093), .A2(n2847), .ZN(n1458) );
  OAI22_X1 U1632 ( .A1(n1458), .A2(n2246), .B1(n2247), .B2(n2847), .ZN(n1519)
         );
  OAI22_X1 U1633 ( .A1(n2113), .A2(n1460), .B1(n1459), .B2(n2112), .ZN(n1550)
         );
  XNOR2_X1 U1634 ( .A(n2153), .B(n16), .ZN(n1515) );
  OAI22_X1 U1635 ( .A1(n1890), .A2(n1515), .B1(n1461), .B2(n1889), .ZN(n1542)
         );
  XNOR2_X1 U1636 ( .A(n1093), .B(n28), .ZN(n1462) );
  OAI22_X1 U1637 ( .A1(n1463), .A2(n2246), .B1(n1462), .B2(n2247), .ZN(n1541)
         );
  XNOR2_X1 U1638 ( .A(n1126), .B(n2147), .ZN(n1464) );
  XNOR2_X1 U1639 ( .A(n1781), .B(n2147), .ZN(n1484) );
  OAI22_X1 U1640 ( .A1(n6131), .A2(n1464), .B1(n6128), .B2(n1484), .ZN(n1540)
         );
  FA_X1 U1641 ( .A(n1467), .B(n1466), .CI(n1465), .CO(n1445), .S(n1534) );
  FA_X1 U1642 ( .A(n1470), .B(n1469), .CI(n1468), .CO(n1743), .S(n1748) );
  FA_X1 U1643 ( .A(n1473), .B(n1472), .CI(n1471), .CO(n1502), .S(n1505) );
  INV_X1 U1644 ( .A(n4660), .ZN(n1474) );
  AND2_X1 U1645 ( .A1(n1126), .A2(n1474), .ZN(n1508) );
  OAI22_X1 U1646 ( .A1(n1476), .A2(n1778), .B1(n1475), .B2(n1777), .ZN(n1507)
         );
  OAI22_X1 U1647 ( .A1(n1931), .A2(n1478), .B1(n6122), .B2(n1477), .ZN(n1506)
         );
  OAI22_X1 U1648 ( .A1(n1480), .A2(n1901), .B1(n1479), .B2(n1903), .ZN(n1511)
         );
  OAI22_X1 U1649 ( .A1(n1482), .A2(n2080), .B1(n1481), .B2(n2079), .ZN(n1510)
         );
  OAI22_X1 U1650 ( .A1(n6130), .A2(n1484), .B1(n6128), .B2(n1483), .ZN(n1509)
         );
  FA_X1 U1651 ( .A(n1487), .B(n1486), .CI(n1485), .CO(n1472), .S(n1522) );
  FA_X1 U1652 ( .A(n1490), .B(n1489), .CI(n1488), .CO(n1471), .S(n1527) );
  FA_X1 U1653 ( .A(n1493), .B(n1492), .CI(n1491), .CO(n1473), .S(n1526) );
  FA_X1 U1654 ( .A(n1496), .B(n1495), .CI(n1494), .CO(n1449), .S(n1525) );
  FA_X1 U1655 ( .A(n1499), .B(n1498), .CI(n1497), .CO(n1371), .S(n1739) );
  FA_X1 U1656 ( .A(n1502), .B(n1501), .CI(n1500), .CO(n1735), .S(n1738) );
  FA_X1 U1657 ( .A(n1505), .B(n1504), .CI(n1503), .CO(n1740), .S(n1533) );
  FA_X1 U1658 ( .A(n1508), .B(n1507), .CI(n1506), .CO(n1524), .S(n1563) );
  FA_X1 U1659 ( .A(n1511), .B(n1510), .CI(n1509), .CO(n1523), .S(n1562) );
  XNOR2_X1 U1660 ( .A(n2103), .B(n1612), .ZN(n1568) );
  OAI22_X1 U1661 ( .A1(n1568), .A2(n1778), .B1(n1512), .B2(n1777), .ZN(n1600)
         );
  XNOR2_X1 U1662 ( .A(n1825), .B(n1808), .ZN(n1565) );
  OAI22_X1 U1663 ( .A1(n1565), .A2(n1901), .B1(n1513), .B2(n1903), .ZN(n1599)
         );
  INV_X1 U1664 ( .A(n2233), .ZN(n1514) );
  AND2_X1 U1665 ( .A1(n1126), .A2(n1514), .ZN(n1598) );
  XNOR2_X1 U1666 ( .A(n2109), .B(n16), .ZN(n1571) );
  OAI22_X1 U1667 ( .A1(n1890), .A2(n1571), .B1(n1515), .B2(n1889), .ZN(n1574)
         );
  XNOR2_X1 U1668 ( .A(n1812), .B(n1785), .ZN(n1570) );
  OAI22_X1 U1669 ( .A1(n1516), .A2(n2079), .B1(n1570), .B2(n2080), .ZN(n1573)
         );
  HA_X1 U1670 ( .A(n1518), .B(n1517), .CO(n1521), .S(n1572) );
  FA_X1 U1671 ( .A(n1521), .B(n1520), .CI(n1519), .CO(n1551), .S(n1578) );
  FA_X1 U1672 ( .A(n1524), .B(n1523), .CI(n1522), .CO(n1504), .S(n1556) );
  FA_X1 U1673 ( .A(n1527), .B(n1526), .CI(n1525), .CO(n1503), .S(n1555) );
  FA_X1 U1674 ( .A(n1530), .B(n1529), .CI(n1528), .CO(n1749), .S(n1531) );
  NOR2_X1 U1675 ( .A1(n1729), .A2(n1728), .ZN(n5443) );
  FA_X1 U1676 ( .A(n1533), .B(n1532), .CI(n1531), .CO(n1728), .S(n1727) );
  FA_X1 U1677 ( .A(n1536), .B(n1535), .CI(n1534), .CO(n1528), .S(n1560) );
  FA_X1 U1678 ( .A(n1539), .B(n1538), .CI(n1537), .CO(n1553), .S(n1589) );
  FA_X1 U1679 ( .A(n1542), .B(n1541), .CI(n1540), .CO(n1549), .S(n1588) );
  XNOR2_X1 U1680 ( .A(n58), .B(n1781), .ZN(n1566) );
  OAI22_X1 U1681 ( .A1(n2113), .A2(n1566), .B1(n1543), .B2(n2112), .ZN(n1603)
         );
  XNOR2_X1 U1682 ( .A(n1819), .B(n69), .ZN(n1564) );
  OAI22_X1 U1683 ( .A1(n1931), .A2(n1564), .B1(n6122), .B2(n1544), .ZN(n1602)
         );
  INV_X1 U1684 ( .A(n2079), .ZN(n1545) );
  AND2_X1 U1685 ( .A1(n1093), .A2(n1545), .ZN(n1595) );
  INV_X1 U1686 ( .A(dot_op_b_i[20]), .ZN(n1546) );
  INV_X1 U1687 ( .A(dot_op_c_i[4]), .ZN(n2457) );
  OAI22_X1 U1688 ( .A1(n1131), .A2(n1546), .B1(n1661), .B2(n2457), .ZN(n1594)
         );
  INV_X1 U1689 ( .A(dot_op_b_i[21]), .ZN(n1547) );
  INV_X1 U1690 ( .A(dot_op_c_i[5]), .ZN(n2446) );
  OAI22_X1 U1691 ( .A1(n1131), .A2(n1547), .B1(n1661), .B2(n2446), .ZN(n1685)
         );
  OR2_X1 U1692 ( .A1(n1093), .A2(n3015), .ZN(n1548) );
  OAI22_X1 U1693 ( .A1(n1548), .A2(n2079), .B1(n2080), .B2(n3015), .ZN(n1684)
         );
  FA_X1 U1694 ( .A(n1551), .B(n1550), .CI(n1549), .CO(n1535), .S(n1582) );
  FA_X1 U1695 ( .A(n1554), .B(n1553), .CI(n1552), .CO(n1536), .S(n1581) );
  FA_X1 U1696 ( .A(n1557), .B(n1556), .CI(n1555), .CO(n1532), .S(n1558) );
  NOR2_X1 U1697 ( .A1(n1727), .A2(n1726), .ZN(n5441) );
  NOR2_X1 U1698 ( .A1(n5443), .A2(n5441), .ZN(n1731) );
  FA_X1 U1699 ( .A(n1560), .B(n1559), .CI(n1558), .CO(n1726), .S(n1722) );
  FA_X1 U1700 ( .A(n1563), .B(n1562), .CI(n1561), .CO(n1557), .S(n1586) );
  XNOR2_X1 U1701 ( .A(n1905), .B(n69), .ZN(n1597) );
  OAI22_X1 U1702 ( .A1(n1931), .A2(n1597), .B1(n6122), .B2(n1564), .ZN(n1689)
         );
  XNOR2_X1 U1703 ( .A(n1770), .B(n1808), .ZN(n1590) );
  OAI22_X1 U1704 ( .A1(n1590), .A2(n1901), .B1(n1565), .B2(n1903), .ZN(n1688)
         );
  XNOR2_X1 U1705 ( .A(n58), .B(n1126), .ZN(n1567) );
  OAI22_X1 U1706 ( .A1(n2113), .A2(n1567), .B1(n1566), .B2(n50), .ZN(n1687) );
  XNOR2_X1 U1707 ( .A(n1804), .B(n1612), .ZN(n1591) );
  OAI22_X1 U1708 ( .A1(n1591), .A2(n1778), .B1(n1568), .B2(n1777), .ZN(n1683)
         );
  XNOR2_X1 U1709 ( .A(n1093), .B(n1785), .ZN(n1569) );
  OAI22_X1 U1710 ( .A1(n1570), .A2(n2079), .B1(n1569), .B2(n2080), .ZN(n1682)
         );
  XNOR2_X1 U1711 ( .A(n1784), .B(n16), .ZN(n1596) );
  OAI22_X1 U1712 ( .A1(n1890), .A2(n1596), .B1(n1571), .B2(n1889), .ZN(n1681)
         );
  FA_X1 U1713 ( .A(n1574), .B(n1573), .CI(n1572), .CO(n1579), .S(n1696) );
  FA_X1 U1714 ( .A(n1577), .B(n1576), .CI(n1575), .CO(n1554), .S(n1605) );
  FA_X1 U1715 ( .A(n1580), .B(n1579), .CI(n1578), .CO(n1561), .S(n1604) );
  FA_X1 U1716 ( .A(n1583), .B(n1582), .CI(n1581), .CO(n1559), .S(n1584) );
  OR2_X1 U1717 ( .A1(n1722), .A2(n1721), .ZN(n5414) );
  FA_X1 U1718 ( .A(n1586), .B(n1585), .CI(n1584), .CO(n1721), .S(n1720) );
  FA_X1 U1719 ( .A(n1589), .B(n1588), .CI(n1587), .CO(n1583), .S(n1712) );
  XNOR2_X1 U1720 ( .A(n1812), .B(n1808), .ZN(n1622) );
  OAI22_X1 U1721 ( .A1(n1590), .A2(n1903), .B1(n1622), .B2(n1901), .ZN(n1643)
         );
  AND2_X1 U1722 ( .A1(n1126), .A2(n49), .ZN(n1642) );
  XNOR2_X1 U1723 ( .A(n1825), .B(n1612), .ZN(n1618) );
  OAI22_X1 U1724 ( .A1(n1618), .A2(n1778), .B1(n1591), .B2(n1777), .ZN(n1641)
         );
  INV_X1 U1725 ( .A(n58), .ZN(n1593) );
  OR2_X1 U1726 ( .A1(n1126), .A2(n1593), .ZN(n1592) );
  OAI22_X1 U1727 ( .A1(n2113), .A2(n1593), .B1(n1592), .B2(n50), .ZN(n1676) );
  HA_X1 U1728 ( .A(n1595), .B(n1594), .CO(n1686), .S(n1617) );
  XNOR2_X1 U1729 ( .A(n1819), .B(n16), .ZN(n1623) );
  OAI22_X1 U1730 ( .A1(n1890), .A2(n1623), .B1(n1596), .B2(n1889), .ZN(n1616)
         );
  XNOR2_X1 U1731 ( .A(n1781), .B(n69), .ZN(n1609) );
  OAI22_X1 U1732 ( .A1(n1931), .A2(n1609), .B1(n6122), .B2(n1597), .ZN(n1615)
         );
  FA_X1 U1733 ( .A(n1600), .B(n1599), .CI(n1598), .CO(n1580), .S(n1703) );
  FA_X1 U1734 ( .A(n1603), .B(n1602), .CI(n1601), .CO(n1587), .S(n1702) );
  FA_X1 U1735 ( .A(n1606), .B(n1605), .CI(n1604), .CO(n1585), .S(n1710) );
  OR2_X1 U1736 ( .A1(n1720), .A2(n1719), .ZN(n5411) );
  NAND2_X1 U1737 ( .A1(n5414), .A2(n5411), .ZN(n1725) );
  INV_X1 U1738 ( .A(n1916), .ZN(n1608) );
  OR2_X1 U1739 ( .A1(n1126), .A2(n1608), .ZN(n1607) );
  OAI22_X1 U1740 ( .A1(n1931), .A2(n1608), .B1(n6122), .B2(n1607), .ZN(n1649)
         );
  XNOR2_X1 U1741 ( .A(n1126), .B(n69), .ZN(n1610) );
  OAI22_X1 U1742 ( .A1(n1931), .A2(n1610), .B1(n6122), .B2(n1609), .ZN(n1648)
         );
  INV_X1 U1743 ( .A(n1932), .ZN(n1611) );
  AND2_X1 U1744 ( .A1(n1126), .A2(n1611), .ZN(n1655) );
  XNOR2_X1 U1745 ( .A(n1770), .B(n1612), .ZN(n1619) );
  XNOR2_X1 U1746 ( .A(n1812), .B(n1612), .ZN(n1633) );
  OAI22_X1 U1747 ( .A1(n1619), .A2(n1777), .B1(n1633), .B2(n1778), .ZN(n1654)
         );
  INV_X1 U1748 ( .A(n1903), .ZN(n1613) );
  AND2_X1 U1749 ( .A1(n1093), .A2(n1613), .ZN(n1625) );
  INV_X1 U1750 ( .A(dot_op_b_i[18]), .ZN(n1614) );
  INV_X1 U1751 ( .A(dot_op_c_i[2]), .ZN(n2466) );
  OAI22_X1 U1752 ( .A1(n12), .A2(n1614), .B1(n1661), .B2(n2466), .ZN(n1624) );
  FA_X1 U1753 ( .A(n1617), .B(n1616), .CI(n1615), .CO(n1675), .S(n1691) );
  OAI22_X1 U1754 ( .A1(n1619), .A2(n1778), .B1(n1618), .B2(n1777), .ZN(n1637)
         );
  XNOR2_X1 U1755 ( .A(n1093), .B(n1808), .ZN(n1621) );
  OAI22_X1 U1756 ( .A1(n1622), .A2(n1903), .B1(n1621), .B2(n1901), .ZN(n1636)
         );
  XNOR2_X1 U1757 ( .A(n1905), .B(n16), .ZN(n1630) );
  OAI22_X1 U1758 ( .A1(n1890), .A2(n1630), .B1(n1623), .B2(n1889), .ZN(n1635)
         );
  HA_X1 U1759 ( .A(n1625), .B(n1624), .CO(n1640), .S(n1653) );
  INV_X1 U1760 ( .A(dot_op_b_i[19]), .ZN(n1626) );
  INV_X1 U1761 ( .A(dot_op_c_i[3]), .ZN(n2468) );
  OAI22_X1 U1762 ( .A1(n12), .A2(n1626), .B1(n1661), .B2(n2468), .ZN(n1639) );
  OR2_X1 U1763 ( .A1(n1093), .A2(n3078), .ZN(n1627) );
  OAI22_X1 U1764 ( .A1(n1627), .A2(n1903), .B1(n1901), .B2(n3078), .ZN(n1638)
         );
  OR2_X1 U1765 ( .A1(n1093), .A2(n1628), .ZN(n1629) );
  NAND2_X1 U1766 ( .A1(n1778), .A2(n1629), .ZN(n1660) );
  INV_X1 U1767 ( .A(dot_op_c_i[1]), .ZN(n2526) );
  OAI22_X1 U1768 ( .A1(n12), .A2(n2511), .B1(n1661), .B2(n2526), .ZN(n1659) );
  XNOR2_X1 U1769 ( .A(n1781), .B(n16), .ZN(n1634) );
  OAI22_X1 U1770 ( .A1(n1890), .A2(n1634), .B1(n1630), .B2(n1889), .ZN(n1651)
         );
  INV_X1 U1771 ( .A(n16), .ZN(n1631) );
  OR2_X1 U1772 ( .A1(n1126), .A2(n1631), .ZN(n1632) );
  NAND2_X1 U1773 ( .A1(n1632), .A2(n1890), .ZN(n1658) );
  OAI22_X1 U1774 ( .A1(n1633), .A2(n1777), .B1(n1093), .B2(n1778), .ZN(n1657)
         );
  OAI22_X1 U1775 ( .A1(n1890), .A2(n1126), .B1(n1634), .B2(n1889), .ZN(n1656)
         );
  FA_X1 U1776 ( .A(n1637), .B(n1636), .CI(n1635), .CO(n1680), .S(n1646) );
  FA_X1 U1777 ( .A(n1640), .B(n1639), .CI(n1638), .CO(n1679), .S(n1645) );
  FA_X1 U1778 ( .A(n1643), .B(n1642), .CI(n1641), .CO(n1677), .S(n1678) );
  NOR2_X1 U1779 ( .A1(n1674), .A2(n1673), .ZN(n2813) );
  FA_X1 U1780 ( .A(n1646), .B(n1645), .CI(n1644), .CO(n1690), .S(n1671) );
  FA_X1 U1781 ( .A(n1649), .B(n1648), .CI(n1647), .CO(n1692), .S(n1670) );
  OR2_X1 U1782 ( .A1(n1671), .A2(n1670), .ZN(n2749) );
  FA_X1 U1783 ( .A(n1652), .B(n1651), .CI(n1650), .CO(n1644), .S(n1669) );
  FA_X1 U1784 ( .A(n1655), .B(n1654), .CI(n1653), .CO(n1647), .S(n1668) );
  NOR2_X1 U1785 ( .A1(n1669), .A2(n1668), .ZN(n5316) );
  FA_X1 U1786 ( .A(n1658), .B(n1657), .CI(n1656), .CO(n1650), .S(n1665) );
  HA_X1 U1787 ( .A(n1660), .B(n1659), .CO(n1652), .S(n1664) );
  NOR2_X1 U1788 ( .A1(n1665), .A2(n1664), .ZN(n5278) );
  AND2_X1 U1789 ( .A1(n1093), .A2(dot_op_a_i[0]), .ZN(n5240) );
  INV_X1 U1790 ( .A(dot_op_b_i[16]), .ZN(n1662) );
  INV_X1 U1791 ( .A(dot_op_c_i[0]), .ZN(n2523) );
  OAI22_X1 U1792 ( .A1(n12), .A2(n1662), .B1(n1661), .B2(n2523), .ZN(n5239) );
  AND2_X1 U1793 ( .A1(n1126), .A2(n1663), .ZN(n5238) );
  INV_X1 U1794 ( .A(n5281), .ZN(n1666) );
  NAND2_X1 U1795 ( .A1(n1665), .A2(n1664), .ZN(n5279) );
  OAI21_X1 U1796 ( .B1(n5278), .B2(n1666), .A(n5279), .ZN(n1667) );
  INV_X1 U1797 ( .A(n1667), .ZN(n5319) );
  NAND2_X1 U1798 ( .A1(n1669), .A2(n1668), .ZN(n5317) );
  OAI21_X1 U1799 ( .B1(n5316), .B2(n5319), .A(n5317), .ZN(n2750) );
  NAND2_X1 U1800 ( .A1(n1671), .A2(n1670), .ZN(n2748) );
  INV_X1 U1801 ( .A(n2748), .ZN(n1672) );
  AOI21_X1 U1802 ( .B1(n2749), .B2(n2750), .A(n1672), .ZN(n2816) );
  NAND2_X1 U1803 ( .A1(n1674), .A2(n1673), .ZN(n2814) );
  OAI21_X1 U1804 ( .B1(n2813), .B2(n2816), .A(n2814), .ZN(n2656) );
  FA_X1 U1805 ( .A(n1677), .B(n1676), .CI(n1675), .CO(n1704), .S(n1707) );
  FA_X1 U1806 ( .A(n1680), .B(n1679), .CI(n1678), .CO(n1706), .S(n1673) );
  FA_X1 U1807 ( .A(n1683), .B(n1682), .CI(n1681), .CO(n1697), .S(n1701) );
  FA_X1 U1808 ( .A(n1686), .B(n1685), .CI(n1684), .CO(n1601), .S(n1700) );
  FA_X1 U1809 ( .A(n1689), .B(n1688), .CI(n1687), .CO(n1698), .S(n1699) );
  FA_X1 U1810 ( .A(n1692), .B(n1691), .CI(n1690), .CO(n1693), .S(n1674) );
  OR2_X1 U1811 ( .A1(n1694), .A2(n1693), .ZN(n2655) );
  NAND2_X1 U1812 ( .A1(n1694), .A2(n1693), .ZN(n2654) );
  INV_X1 U1813 ( .A(n2654), .ZN(n1695) );
  AOI21_X1 U1814 ( .B1(n2656), .B2(n2655), .A(n1695), .ZN(n5362) );
  FA_X1 U1815 ( .A(n1698), .B(n1697), .CI(n1696), .CO(n1606), .S(n1715) );
  FA_X1 U1816 ( .A(n1701), .B(n1700), .CI(n1699), .CO(n1714), .S(n1705) );
  FA_X1 U1817 ( .A(n1704), .B(n1703), .CI(n1702), .CO(n1711), .S(n1713) );
  FA_X1 U1818 ( .A(n1707), .B(n1706), .CI(n1705), .CO(n1708), .S(n1694) );
  NOR2_X1 U1819 ( .A1(n1709), .A2(n1708), .ZN(n5359) );
  NAND2_X1 U1820 ( .A1(n1709), .A2(n1708), .ZN(n5360) );
  OAI21_X1 U1821 ( .B1(n5362), .B2(n5359), .A(n5360), .ZN(n5048) );
  FA_X1 U1822 ( .A(n1712), .B(n1711), .CI(n1710), .CO(n1719), .S(n1717) );
  FA_X1 U1823 ( .A(n1715), .B(n1714), .CI(n1713), .CO(n1716), .S(n1709) );
  OR2_X1 U1824 ( .A1(n1717), .A2(n1716), .ZN(n5047) );
  NAND2_X1 U1825 ( .A1(n1717), .A2(n1716), .ZN(n5046) );
  INV_X1 U1826 ( .A(n5046), .ZN(n1718) );
  AOI21_X1 U1827 ( .B1(n5048), .B2(n5047), .A(n1718), .ZN(n5394) );
  NAND2_X1 U1828 ( .A1(n1720), .A2(n1719), .ZN(n5393) );
  INV_X1 U1829 ( .A(n5393), .ZN(n5410) );
  NAND2_X1 U1830 ( .A1(n1722), .A2(n1721), .ZN(n5413) );
  INV_X1 U1831 ( .A(n5413), .ZN(n1723) );
  AOI21_X1 U1832 ( .B1(n5414), .B2(n5410), .A(n1723), .ZN(n1724) );
  OAI21_X1 U1833 ( .B1(n1725), .B2(n5394), .A(n1724), .ZN(n4994) );
  NAND2_X1 U1834 ( .A1(n1727), .A2(n1726), .ZN(n5440) );
  NAND2_X1 U1835 ( .A1(n1729), .A2(n1728), .ZN(n5444) );
  OAI21_X1 U1836 ( .B1(n5443), .B2(n5440), .A(n5444), .ZN(n1730) );
  AOI21_X1 U1837 ( .B1(n1731), .B2(n4994), .A(n1730), .ZN(n5470) );
  FA_X1 U1838 ( .A(n1734), .B(n1733), .CI(n1732), .CO(n1760), .S(n1753) );
  FA_X1 U1839 ( .A(n1737), .B(n1736), .CI(n1735), .CO(n1376), .S(n1746) );
  FA_X1 U1840 ( .A(n1740), .B(n1739), .CI(n1738), .CO(n1745), .S(n1747) );
  FA_X1 U1841 ( .A(n1743), .B(n1742), .CI(n1741), .CO(n1733), .S(n1744) );
  OR2_X1 U1842 ( .A1(n1753), .A2(n1752), .ZN(n5503) );
  FA_X1 U1843 ( .A(n1746), .B(n1745), .CI(n1744), .CO(n1752), .S(n1751) );
  FA_X1 U1844 ( .A(n1749), .B(n1748), .CI(n1747), .CO(n1750), .S(n1729) );
  OR2_X1 U1845 ( .A1(n1751), .A2(n1750), .ZN(n5500) );
  NAND2_X1 U1846 ( .A1(n5503), .A2(n5500), .ZN(n1756) );
  NAND2_X1 U1847 ( .A1(n1751), .A2(n1750), .ZN(n5471) );
  INV_X1 U1848 ( .A(n5471), .ZN(n5499) );
  NAND2_X1 U1849 ( .A1(n1753), .A2(n1752), .ZN(n5502) );
  INV_X1 U1850 ( .A(n5502), .ZN(n1754) );
  AOI21_X1 U1851 ( .B1(n5503), .B2(n5499), .A(n1754), .ZN(n1755) );
  OAI21_X1 U1852 ( .B1(n5470), .B2(n1756), .A(n1755), .ZN(n4912) );
  NAND2_X1 U1853 ( .A1(n1757), .A2(n4912), .ZN(n1767) );
  NAND2_X1 U1854 ( .A1(n1759), .A2(n1758), .ZN(n4916) );
  NAND2_X1 U1855 ( .A1(n1761), .A2(n1760), .ZN(n5531) );
  INV_X1 U1856 ( .A(n5531), .ZN(n1765) );
  NAND2_X1 U1857 ( .A1(n1763), .A2(n1762), .ZN(n5160) );
  INV_X1 U1858 ( .A(n5160), .ZN(n1764) );
  AOI21_X1 U1859 ( .B1(n5161), .B2(n1765), .A(n1764), .ZN(n4913) );
  XNOR2_X1 U1860 ( .A(n1784), .B(n15), .ZN(n1768) );
  NOR2_X1 U1861 ( .A1(n1768), .A2(n5109), .ZN(n2117) );
  INV_X1 U1862 ( .A(n1804), .ZN(n1769) );
  NOR2_X1 U1863 ( .A1(n1769), .A2(n5116), .ZN(n2116) );
  XNOR2_X1 U1864 ( .A(n5085), .B(n1785), .ZN(n2078) );
  XNOR2_X1 U1865 ( .A(n5115), .B(n1785), .ZN(n1933) );
  OAI22_X1 U1866 ( .A1(n2078), .A2(n2079), .B1(n1933), .B2(n2080), .ZN(n2115)
         );
  XNOR2_X1 U1867 ( .A(n2109), .B(n17), .ZN(n1831) );
  XNOR2_X1 U1868 ( .A(n2153), .B(n17), .ZN(n2100) );
  OAI22_X1 U1869 ( .A1(n5113), .A2(n1831), .B1(n2100), .B2(n6114), .ZN(n2093)
         );
  XNOR2_X1 U1870 ( .A(n4742), .B(n1307), .ZN(n1837) );
  XNOR2_X1 U1871 ( .A(n4795), .B(n1307), .ZN(n2108) );
  OAI22_X1 U1872 ( .A1(n1837), .A2(n4630), .B1(n2108), .B2(n4629), .ZN(n2092)
         );
  XNOR2_X1 U1873 ( .A(n2226), .B(n6111), .ZN(n1835) );
  XNOR2_X1 U1874 ( .A(n4590), .B(n6111), .ZN(n2102) );
  OAI22_X1 U1875 ( .A1(n6125), .A2(n1835), .B1(n6123), .B2(n2102), .ZN(n2091)
         );
  XNOR2_X1 U1876 ( .A(n4683), .B(n4657), .ZN(n1821) );
  XNOR2_X1 U1877 ( .A(n4683), .B(n4681), .ZN(n2076) );
  OAI22_X1 U1878 ( .A1(n4732), .A2(n1821), .B1(n2076), .B2(n4731), .ZN(n2120)
         );
  XNOR2_X1 U1879 ( .A(n4740), .B(n4587), .ZN(n1772) );
  XNOR2_X1 U1880 ( .A(n4780), .B(n4587), .ZN(n2077) );
  OAI22_X1 U1881 ( .A1(n4661), .A2(n1772), .B1(n4660), .B2(n2077), .ZN(n2119)
         );
  XNOR2_X1 U1882 ( .A(n58), .B(n5107), .ZN(n1818) );
  XNOR2_X1 U1883 ( .A(n5083), .B(n58), .ZN(n2111) );
  OAI22_X1 U1884 ( .A1(n2113), .A2(n1818), .B1(n2111), .B2(n50), .ZN(n2118) );
  INV_X1 U1885 ( .A(n1770), .ZN(n1771) );
  NOR2_X1 U1886 ( .A1(n1771), .A2(n5116), .ZN(n1811) );
  INV_X1 U1887 ( .A(dot_op_c_i[18]), .ZN(n5187) );
  OAI21_X1 U1888 ( .B1(n1661), .B2(n5187), .A(n5114), .ZN(n1810) );
  OR2_X1 U1889 ( .A1(n1811), .A2(n1810), .ZN(n1824) );
  XNOR2_X1 U1890 ( .A(n4681), .B(n4587), .ZN(n1914) );
  OAI22_X1 U1891 ( .A1(n4661), .A2(n1914), .B1(n4660), .B2(n1772), .ZN(n1823)
         );
  XNOR2_X1 U1892 ( .A(n5085), .B(n1808), .ZN(n1904) );
  AOI21_X1 U1893 ( .B1(n1901), .B2(n1903), .A(n1904), .ZN(n1773) );
  INV_X1 U1894 ( .A(n1773), .ZN(n1822) );
  XNOR2_X1 U1895 ( .A(n4839), .B(n28), .ZN(n1827) );
  XNOR2_X1 U1896 ( .A(n5076), .B(n28), .ZN(n2114) );
  OAI22_X1 U1897 ( .A1(n1827), .A2(n2247), .B1(n2114), .B2(n2246), .ZN(n2090)
         );
  INV_X1 U1898 ( .A(dot_op_c_i[20]), .ZN(n4243) );
  OAI21_X1 U1899 ( .B1(n1661), .B2(n4243), .A(n5114), .ZN(n2089) );
  XNOR2_X1 U1900 ( .A(n2214), .B(n30), .ZN(n1841) );
  XNOR2_X1 U1901 ( .A(n4592), .B(n30), .ZN(n2107) );
  OAI22_X1 U1902 ( .A1(n1841), .A2(n4830), .B1(n2107), .B2(n4829), .ZN(n2088)
         );
  XNOR2_X1 U1903 ( .A(n2103), .B(n1803), .ZN(n1839) );
  XNOR2_X1 U1904 ( .A(n2169), .B(n1803), .ZN(n2101) );
  OAI22_X1 U1905 ( .A1(n1839), .A2(n5124), .B1(n2101), .B2(n5123), .ZN(n2087)
         );
  XNOR2_X1 U1906 ( .A(n4655), .B(n4679), .ZN(n1833) );
  XNOR2_X1 U1907 ( .A(n4673), .B(n4679), .ZN(n2105) );
  OAI22_X1 U1908 ( .A1(n1833), .A2(n4746), .B1(n2105), .B2(n4745), .ZN(n2086)
         );
  XNOR2_X1 U1909 ( .A(n4841), .B(n2147), .ZN(n1829) );
  XNOR2_X1 U1910 ( .A(n5078), .B(n2147), .ZN(n2106) );
  OAI22_X1 U1911 ( .A1(n6130), .A2(n1829), .B1(n6128), .B2(n2106), .ZN(n2085)
         );
  XNOR2_X1 U1912 ( .A(n58), .B(n4841), .ZN(n1913) );
  OAI22_X1 U1913 ( .A1(n2113), .A2(n1774), .B1(n1913), .B2(n50), .ZN(n1867) );
  XNOR2_X1 U1914 ( .A(n4657), .B(n4587), .ZN(n1915) );
  OAI22_X1 U1915 ( .A1(n4661), .A2(n1775), .B1(n4660), .B2(n1915), .ZN(n1866)
         );
  AOI21_X1 U1916 ( .B1(n1778), .B2(n1777), .A(n1776), .ZN(n1779) );
  INV_X1 U1917 ( .A(n1779), .ZN(n1865) );
  XNOR2_X1 U1918 ( .A(n5107), .B(n69), .ZN(n1917) );
  OAI22_X1 U1919 ( .A1(n1931), .A2(n1780), .B1(n6122), .B2(n1917), .ZN(n1870)
         );
  XNOR2_X1 U1920 ( .A(n1781), .B(n15), .ZN(n1782) );
  NOR2_X1 U1921 ( .A1(n1782), .A2(n5109), .ZN(n1869) );
  XNOR2_X1 U1922 ( .A(n4683), .B(n2226), .ZN(n1908) );
  OAI22_X1 U1923 ( .A1(n4732), .A2(n1783), .B1(n1908), .B2(n4731), .ZN(n1868)
         );
  XNOR2_X1 U1924 ( .A(n1819), .B(n17), .ZN(n1816) );
  XNOR2_X1 U1925 ( .A(n1784), .B(n17), .ZN(n1832) );
  OAI22_X1 U1926 ( .A1(n5113), .A2(n1816), .B1(n1832), .B2(n6114), .ZN(n1802)
         );
  XNOR2_X1 U1927 ( .A(n4839), .B(n1785), .ZN(n1794) );
  XNOR2_X1 U1928 ( .A(n5076), .B(n1785), .ZN(n1934) );
  OAI22_X1 U1929 ( .A1(n1794), .A2(n2080), .B1(n1934), .B2(n2079), .ZN(n1801)
         );
  XNOR2_X1 U1930 ( .A(n2109), .B(n6111), .ZN(n1791) );
  XNOR2_X1 U1931 ( .A(n2153), .B(n6111), .ZN(n1836) );
  OAI22_X1 U1932 ( .A1(n6125), .A2(n1791), .B1(n6123), .B2(n1836), .ZN(n1800)
         );
  XNOR2_X1 U1933 ( .A(n1825), .B(n1803), .ZN(n1805) );
  OAI22_X1 U1934 ( .A1(n1786), .A2(n5124), .B1(n1805), .B2(n5123), .ZN(n1858)
         );
  XNOR2_X1 U1935 ( .A(n4742), .B(n28), .ZN(n1806) );
  OAI22_X1 U1936 ( .A1(n1787), .A2(n2247), .B1(n1806), .B2(n2246), .ZN(n1857)
         );
  XNOR2_X1 U1937 ( .A(n4740), .B(n2147), .ZN(n1807) );
  OAI22_X1 U1938 ( .A1(n6131), .A2(n1788), .B1(n6128), .B2(n1807), .ZN(n1856)
         );
  XNOR2_X1 U1939 ( .A(n2214), .B(n4679), .ZN(n1798) );
  OAI22_X1 U1940 ( .A1(n1789), .A2(n4746), .B1(n1798), .B2(n4745), .ZN(n1855)
         );
  XNOR2_X1 U1941 ( .A(n2103), .B(n30), .ZN(n1797) );
  OAI22_X1 U1942 ( .A1(n1790), .A2(n4830), .B1(n1797), .B2(n4829), .ZN(n1854)
         );
  OAI22_X1 U1943 ( .A1(n6125), .A2(n1792), .B1(n6123), .B2(n1791), .ZN(n1853)
         );
  XNOR2_X1 U1944 ( .A(n4655), .B(n1307), .ZN(n1799) );
  OAI22_X1 U1945 ( .A1(n1793), .A2(n4630), .B1(n1799), .B2(n4629), .ZN(n1861)
         );
  OAI22_X1 U1946 ( .A1(n1795), .A2(n2080), .B1(n1794), .B2(n2079), .ZN(n1860)
         );
  OR2_X1 U1947 ( .A1(n1126), .A2(n53), .ZN(n1796) );
  NOR2_X1 U1948 ( .A1(n1796), .A2(n5109), .ZN(n1859) );
  XNOR2_X1 U1949 ( .A(n2169), .B(n30), .ZN(n1842) );
  OAI22_X1 U1950 ( .A1(n1797), .A2(n4830), .B1(n1842), .B2(n4829), .ZN(n1897)
         );
  XNOR2_X1 U1951 ( .A(n4592), .B(n4679), .ZN(n1834) );
  OAI22_X1 U1952 ( .A1(n1798), .A2(n4746), .B1(n1834), .B2(n4745), .ZN(n1896)
         );
  XNOR2_X1 U1953 ( .A(n4673), .B(n1307), .ZN(n1838) );
  OAI22_X1 U1954 ( .A1(n1799), .A2(n4630), .B1(n1838), .B2(n4629), .ZN(n1895)
         );
  FA_X1 U1955 ( .A(n1802), .B(n1801), .CI(n1800), .CO(n1974), .S(n1877) );
  XNOR2_X1 U1956 ( .A(n1804), .B(n1803), .ZN(n1840) );
  OAI22_X1 U1957 ( .A1(n1805), .A2(n5124), .B1(n1840), .B2(n5123), .ZN(n1900)
         );
  XNOR2_X1 U1958 ( .A(n4795), .B(n28), .ZN(n1828) );
  OAI22_X1 U1959 ( .A1(n1806), .A2(n2247), .B1(n1828), .B2(n2246), .ZN(n1899)
         );
  XNOR2_X1 U1960 ( .A(n4780), .B(n2147), .ZN(n1830) );
  OAI22_X1 U1961 ( .A1(n6131), .A2(n1807), .B1(n6128), .B2(n1830), .ZN(n1898)
         );
  INV_X1 U1962 ( .A(dot_op_c_i[17]), .ZN(n4923) );
  OAI21_X1 U1963 ( .B1(n1661), .B2(n4923), .A(n5114), .ZN(n1849) );
  XNOR2_X1 U1964 ( .A(n5115), .B(n1808), .ZN(n1902) );
  OAI22_X1 U1965 ( .A1(n1809), .A2(n1901), .B1(n1902), .B2(n1903), .ZN(n1848)
         );
  XNOR2_X1 U1966 ( .A(n1811), .B(n1810), .ZN(n1844) );
  INV_X1 U1967 ( .A(n1812), .ZN(n1813) );
  NOR2_X1 U1968 ( .A1(n1813), .A2(n5116), .ZN(n1852) );
  HA_X1 U1969 ( .A(n1815), .B(n1814), .CO(n1851), .S(n1918) );
  OAI22_X1 U1970 ( .A1(n5113), .A2(n1817), .B1(n1816), .B2(n6114), .ZN(n1850)
         );
  XNOR2_X1 U1971 ( .A(n58), .B(n5078), .ZN(n1912) );
  OAI22_X1 U1972 ( .A1(n2113), .A2(n1912), .B1(n1818), .B2(n50), .ZN(n1990) );
  XNOR2_X1 U1973 ( .A(n1819), .B(n15), .ZN(n1820) );
  NOR2_X1 U1974 ( .A1(n1820), .A2(n5109), .ZN(n1989) );
  XNOR2_X1 U1975 ( .A(n4683), .B(n4590), .ZN(n1907) );
  OAI22_X1 U1976 ( .A1(n4732), .A2(n1907), .B1(n1821), .B2(n4731), .ZN(n1988)
         );
  FA_X1 U1977 ( .A(n1824), .B(n1823), .CI(n1822), .CO(n2096), .S(n1994) );
  INV_X1 U1978 ( .A(n1825), .ZN(n1826) );
  NOR2_X1 U1979 ( .A1(n1826), .A2(n5116), .ZN(n1987) );
  OAI22_X1 U1980 ( .A1(n1828), .A2(n2247), .B1(n1827), .B2(n2246), .ZN(n1986)
         );
  OAI22_X1 U1981 ( .A1(n6131), .A2(n1830), .B1(n6128), .B2(n1829), .ZN(n1985)
         );
  OAI22_X1 U1982 ( .A1(n5113), .A2(n1832), .B1(n1831), .B2(n6114), .ZN(n1981)
         );
  OAI22_X1 U1983 ( .A1(n1834), .A2(n4746), .B1(n1833), .B2(n4745), .ZN(n1980)
         );
  OAI22_X1 U1984 ( .A1(n6125), .A2(n1836), .B1(n6123), .B2(n1835), .ZN(n1979)
         );
  OAI22_X1 U1985 ( .A1(n1838), .A2(n4630), .B1(n1837), .B2(n4629), .ZN(n1984)
         );
  OAI22_X1 U1986 ( .A1(n1840), .A2(n5124), .B1(n1839), .B2(n5123), .ZN(n1983)
         );
  OAI22_X1 U1987 ( .A1(n1842), .A2(n4830), .B1(n1841), .B2(n4829), .ZN(n1982)
         );
  FA_X1 U1988 ( .A(n97), .B(n1844), .CI(n1843), .CO(n1996), .S(n1949) );
  FA_X1 U1989 ( .A(n1847), .B(n1846), .CI(n1845), .CO(n1957), .S(n1950) );
  FA_X1 U1990 ( .A(n1852), .B(n1851), .CI(n1850), .CO(n1843), .S(n1956) );
  FA_X1 U1991 ( .A(n1855), .B(n1854), .CI(n1853), .CO(n1875), .S(n1963) );
  FA_X1 U1992 ( .A(n1858), .B(n1857), .CI(n1856), .CO(n1876), .S(n1962) );
  FA_X1 U1993 ( .A(n1861), .B(n1860), .CI(n1859), .CO(n1874), .S(n1961) );
  FA_X1 U1994 ( .A(n1864), .B(n1863), .CI(n1862), .CO(n2124), .S(n2015) );
  FA_X1 U1995 ( .A(n1867), .B(n1866), .CI(n1865), .CO(n1879), .S(n1966) );
  FA_X1 U1996 ( .A(n1870), .B(n1869), .CI(n1868), .CO(n1878), .S(n1965) );
  FA_X1 U1997 ( .A(n1873), .B(n1872), .CI(n1871), .CO(n1964), .S(n2008) );
  FA_X1 U1998 ( .A(n1876), .B(n1875), .CI(n1874), .CO(n1863), .S(n2002) );
  FA_X1 U1999 ( .A(n1879), .B(n1878), .CI(n1877), .CO(n1864), .S(n2001) );
  FA_X1 U2000 ( .A(n1882), .B(n1881), .CI(n1880), .CO(n2006), .S(n2012) );
  FA_X1 U2001 ( .A(n1885), .B(n1884), .CI(n1883), .CO(n2005), .S(n2007) );
  AOI21_X1 U2002 ( .B1(n1890), .B2(n1889), .A(n1888), .ZN(n1891) );
  INV_X1 U2003 ( .A(n1891), .ZN(n1910) );
  FA_X1 U2004 ( .A(n1894), .B(n1893), .CI(n1892), .CO(n1909), .S(n1880) );
  FA_X1 U2005 ( .A(n1897), .B(n1896), .CI(n1895), .CO(n1975), .S(n1943) );
  FA_X1 U2006 ( .A(n1900), .B(n1899), .CI(n1898), .CO(n1973), .S(n1942) );
  OAI22_X1 U2007 ( .A1(n1904), .A2(n1903), .B1(n1902), .B2(n1901), .ZN(n1937)
         );
  XNOR2_X1 U2008 ( .A(n1905), .B(n15), .ZN(n1906) );
  NOR2_X1 U2009 ( .A1(n1906), .A2(n5109), .ZN(n1936) );
  OAI22_X1 U2010 ( .A1(n4732), .A2(n1908), .B1(n1907), .B2(n4731), .ZN(n1935)
         );
  FA_X1 U2011 ( .A(n1911), .B(n1910), .CI(n1909), .CO(n1946), .S(n2004) );
  OAI22_X1 U2012 ( .A1(n2113), .A2(n1913), .B1(n1912), .B2(n50), .ZN(n1940) );
  OAI22_X1 U2013 ( .A1(n4661), .A2(n1915), .B1(n4660), .B2(n1914), .ZN(n1939)
         );
  XNOR2_X1 U2014 ( .A(n5083), .B(n69), .ZN(n1930) );
  OAI22_X1 U2015 ( .A1(n1930), .A2(n6122), .B1(n1931), .B2(n1917), .ZN(n1938)
         );
  FA_X1 U2016 ( .A(n1920), .B(n1919), .CI(n1918), .CO(n1955), .S(n1951) );
  FA_X1 U2017 ( .A(n1923), .B(n1922), .CI(n1921), .CO(n1954), .S(n1882) );
  FA_X1 U2018 ( .A(n1926), .B(n1925), .CI(n1924), .CO(n1953), .S(n1952) );
  FA_X1 U2019 ( .A(n1929), .B(n1928), .CI(n1927), .CO(n2068), .S(n2018) );
  INV_X1 U2020 ( .A(dot_op_c_i[19]), .ZN(n2996) );
  OAI21_X1 U2021 ( .B1(n1661), .B2(n2996), .A(n5114), .ZN(n1977) );
  AOI21_X1 U2022 ( .B1(n1932), .B2(n1931), .A(n1930), .ZN(n1978) );
  OAI22_X1 U2023 ( .A1(n1934), .A2(n2080), .B1(n1933), .B2(n2079), .ZN(n1976)
         );
  FA_X1 U2024 ( .A(n1937), .B(n1936), .CI(n1935), .CO(n1971), .S(n1941) );
  FA_X1 U2025 ( .A(n1940), .B(n1939), .CI(n1938), .CO(n1970), .S(n1945) );
  FA_X1 U2026 ( .A(n1943), .B(n1942), .CI(n1941), .CO(n1968), .S(n1999) );
  FA_X1 U2027 ( .A(n1946), .B(n1945), .CI(n1944), .CO(n1967), .S(n1998) );
  FA_X1 U2028 ( .A(n1949), .B(n1948), .CI(n1947), .CO(n1927), .S(n2033) );
  FA_X1 U2029 ( .A(n1952), .B(n1951), .CI(n1950), .CO(n2027), .S(n2010) );
  FA_X1 U2030 ( .A(n1955), .B(n1954), .CI(n1953), .CO(n1944), .S(n2026) );
  FA_X1 U2031 ( .A(n1957), .B(n98), .CI(n1956), .CO(n1948), .S(n2025) );
  FA_X1 U2032 ( .A(n1960), .B(n1959), .CI(n1958), .CO(n2024), .S(n2030) );
  FA_X1 U2033 ( .A(n1963), .B(n1962), .CI(n1961), .CO(n1947), .S(n2023) );
  FA_X1 U2034 ( .A(n1966), .B(n1965), .CI(n1964), .CO(n2003), .S(n2022) );
  FA_X1 U2035 ( .A(n1969), .B(n1968), .CI(n1967), .CO(n2129), .S(n2017) );
  FA_X1 U2036 ( .A(n1972), .B(n1971), .CI(n1970), .CO(n2123), .S(n1969) );
  FA_X1 U2037 ( .A(n1975), .B(n1974), .CI(n1973), .CO(n2122), .S(n1862) );
  FA_X1 U2038 ( .A(n1977), .B(n1978), .CI(n1976), .CO(n2075), .S(n1972) );
  INV_X1 U2039 ( .A(n1978), .ZN(n2074) );
  FA_X1 U2040 ( .A(n1981), .B(n1980), .CI(n1979), .CO(n2073), .S(n1992) );
  FA_X1 U2041 ( .A(n1984), .B(n1983), .CI(n1982), .CO(n2084), .S(n1991) );
  FA_X1 U2042 ( .A(n1987), .B(n1986), .CI(n1985), .CO(n2083), .S(n1993) );
  FA_X1 U2043 ( .A(n1990), .B(n1989), .CI(n1988), .CO(n2082), .S(n1995) );
  FA_X1 U2044 ( .A(n1993), .B(n1992), .CI(n1991), .CO(n2071), .S(n1928) );
  FA_X1 U2045 ( .A(n1996), .B(n1995), .CI(n1994), .CO(n2070), .S(n1929) );
  FA_X1 U2046 ( .A(n2000), .B(n1999), .CI(n1998), .CO(n2013), .S(n2036) );
  FA_X1 U2047 ( .A(n2003), .B(n2002), .CI(n2001), .CO(n2014), .S(n2035) );
  FA_X1 U2048 ( .A(n2006), .B(n2005), .CI(n2004), .CO(n2000), .S(n2045) );
  FA_X1 U2049 ( .A(n2009), .B(n2008), .CI(n2007), .CO(n2044), .S(n2041) );
  FA_X1 U2050 ( .A(n2012), .B(n2011), .CI(n2010), .CO(n2043), .S(n2042) );
  FA_X1 U2051 ( .A(n2015), .B(n2014), .CI(n2013), .CO(n2067), .S(n2020) );
  FA_X1 U2052 ( .A(n2018), .B(n2017), .CI(n2016), .CO(n2135), .S(n2019) );
  NOR2_X1 U2053 ( .A1(n2062), .A2(n2061), .ZN(n2278) );
  FA_X1 U2054 ( .A(n2021), .B(n2020), .CI(n2019), .CO(n2061), .S(n2060) );
  FA_X1 U2055 ( .A(n2024), .B(n2023), .CI(n2022), .CO(n2031), .S(n2048) );
  FA_X1 U2056 ( .A(n2025), .B(n2026), .CI(n2027), .CO(n2032), .S(n2047) );
  FA_X1 U2057 ( .A(n2030), .B(n2029), .CI(n2028), .CO(n2046), .S(n2053) );
  FA_X1 U2058 ( .A(n2033), .B(n2032), .CI(n2031), .CO(n2016), .S(n2038) );
  FA_X1 U2059 ( .A(n2036), .B(n2035), .CI(n2034), .CO(n2021), .S(n2037) );
  NOR2_X1 U2060 ( .A1(n2278), .A2(n2775), .ZN(n2064) );
  FA_X1 U2061 ( .A(n2039), .B(n2038), .CI(n2037), .CO(n2059), .S(n2058) );
  FA_X1 U2062 ( .A(n2042), .B(n2041), .CI(n2040), .CO(n2051), .S(n2052) );
  FA_X1 U2063 ( .A(n2045), .B(n2043), .CI(n2044), .CO(n2034), .S(n2050) );
  FA_X1 U2064 ( .A(n2048), .B(n2047), .CI(n2046), .CO(n2039), .S(n2049) );
  FA_X1 U2065 ( .A(n2051), .B(n2050), .CI(n2049), .CO(n2057), .S(n2056) );
  FA_X1 U2066 ( .A(n2054), .B(n2053), .CI(n2052), .CO(n2055), .S(n1759) );
  NOR2_X1 U2067 ( .A1(n2056), .A2(n2055), .ZN(n2766) );
  NOR2_X1 U2068 ( .A1(n2768), .A2(n2766), .ZN(n2774) );
  NAND2_X1 U2069 ( .A1(n2064), .A2(n2774), .ZN(n2066) );
  NAND2_X1 U2070 ( .A1(n2056), .A2(n2055), .ZN(n4908) );
  NAND2_X1 U2071 ( .A1(n2058), .A2(n2057), .ZN(n2769) );
  OAI21_X1 U2072 ( .B1(n2768), .B2(n4908), .A(n2769), .ZN(n2773) );
  NAND2_X1 U2073 ( .A1(n2060), .A2(n2059), .ZN(n2776) );
  NAND2_X1 U2074 ( .A1(n2062), .A2(n2061), .ZN(n2279) );
  OAI21_X1 U2075 ( .B1(n2278), .B2(n2776), .A(n2279), .ZN(n2063) );
  AOI21_X1 U2076 ( .B1(n2064), .B2(n2773), .A(n2063), .ZN(n2065) );
  FA_X1 U2077 ( .A(n2069), .B(n2068), .CI(n2067), .CO(n2197), .S(n2133) );
  FA_X1 U2078 ( .A(n2072), .B(n2071), .CI(n2070), .CO(n2194), .S(n2127) );
  FA_X1 U2079 ( .A(n2075), .B(n2074), .CI(n2073), .CO(n2188), .S(n2121) );
  XNOR2_X1 U2080 ( .A(n4683), .B(n4740), .ZN(n2150) );
  OAI22_X1 U2081 ( .A1(n4732), .A2(n2076), .B1(n2150), .B2(n4731), .ZN(n2173)
         );
  XNOR2_X1 U2082 ( .A(n4841), .B(n4587), .ZN(n2161) );
  OAI22_X1 U2083 ( .A1(n4661), .A2(n2077), .B1(n4660), .B2(n2161), .ZN(n2172)
         );
  AOI21_X1 U2084 ( .B1(n2080), .B2(n2079), .A(n2078), .ZN(n2081) );
  INV_X1 U2085 ( .A(n2081), .ZN(n2171) );
  FA_X1 U2086 ( .A(n2084), .B(n2083), .CI(n2082), .CO(n2186), .S(n2072) );
  FA_X1 U2087 ( .A(n2087), .B(n2086), .CI(n2085), .CO(n2157), .S(n2094) );
  FA_X1 U2088 ( .A(n2090), .B(n2089), .CI(n2088), .CO(n2156), .S(n2095) );
  FA_X1 U2089 ( .A(n2093), .B(n2092), .CI(n2091), .CO(n2155), .S(n2098) );
  FA_X1 U2090 ( .A(n2096), .B(n2095), .CI(n2094), .CO(n2145), .S(n2125) );
  FA_X1 U2091 ( .A(n2099), .B(n2098), .CI(n2097), .CO(n2144), .S(n2126) );
  XNOR2_X1 U2092 ( .A(n2226), .B(n17), .ZN(n2174) );
  OAI22_X1 U2093 ( .A1(n5113), .A2(n2100), .B1(n2174), .B2(n6114), .ZN(n2182)
         );
  XNOR2_X1 U2094 ( .A(n2214), .B(n1803), .ZN(n2151) );
  OAI22_X1 U2095 ( .A1(n2101), .A2(n5124), .B1(n2151), .B2(n5123), .ZN(n2181)
         );
  XNOR2_X1 U2096 ( .A(n4657), .B(n6111), .ZN(n2176) );
  OAI22_X1 U2097 ( .A1(n6125), .A2(n2102), .B1(n6123), .B2(n2176), .ZN(n2180)
         );
  INV_X1 U2098 ( .A(n2103), .ZN(n2104) );
  NOR2_X1 U2099 ( .A1(n2104), .A2(n5116), .ZN(n2179) );
  XNOR2_X1 U2100 ( .A(n4742), .B(n4679), .ZN(n2175) );
  OAI22_X1 U2101 ( .A1(n2105), .A2(n4746), .B1(n2175), .B2(n4745), .ZN(n2178)
         );
  XNOR2_X1 U2102 ( .A(n5107), .B(n2147), .ZN(n2148) );
  OAI22_X1 U2103 ( .A1(n6131), .A2(n2106), .B1(n6128), .B2(n2148), .ZN(n2177)
         );
  XNOR2_X1 U2104 ( .A(n4655), .B(n30), .ZN(n2152) );
  OAI22_X1 U2105 ( .A1(n2107), .A2(n4830), .B1(n2152), .B2(n4829), .ZN(n2185)
         );
  XNOR2_X1 U2106 ( .A(n4839), .B(n1307), .ZN(n2168) );
  OAI22_X1 U2107 ( .A1(n2108), .A2(n4630), .B1(n2168), .B2(n4629), .ZN(n2184)
         );
  XNOR2_X1 U2108 ( .A(n2109), .B(n15), .ZN(n2110) );
  NOR2_X1 U2109 ( .A1(n2110), .A2(n5109), .ZN(n2183) );
  INV_X1 U2110 ( .A(dot_op_c_i[21]), .ZN(n4087) );
  OAI21_X1 U2111 ( .B1(n1661), .B2(n4087), .A(n5114), .ZN(n2164) );
  AOI21_X1 U2112 ( .B1(n2113), .B2(n50), .A(n2111), .ZN(n2163) );
  XNOR2_X1 U2113 ( .A(n5115), .B(n28), .ZN(n2149) );
  OAI22_X1 U2114 ( .A1(n2114), .A2(n2247), .B1(n2149), .B2(n2246), .ZN(n2162)
         );
  FA_X1 U2115 ( .A(n2117), .B(n2116), .CI(n2115), .CO(n2159), .S(n2099) );
  FA_X1 U2116 ( .A(n2120), .B(n2119), .CI(n2118), .CO(n2158), .S(n2097) );
  FA_X1 U2117 ( .A(n2123), .B(n2122), .CI(n2121), .CO(n2189), .S(n2128) );
  FA_X1 U2118 ( .A(n2126), .B(n2125), .CI(n2124), .CO(n2142), .S(n2069) );
  FA_X1 U2119 ( .A(n2129), .B(n2128), .CI(n2127), .CO(n2141), .S(n2134) );
  NAND2_X1 U2120 ( .A1(n2131), .A2(n2130), .ZN(n2132) );
  NAND2_X1 U2121 ( .A1(n2133), .A2(n2132), .ZN(n2137) );
  NAND2_X1 U2122 ( .A1(n2135), .A2(n2134), .ZN(n2136) );
  NAND2_X1 U2123 ( .A1(n2137), .A2(n2136), .ZN(n2138) );
  NOR2_X1 U2124 ( .A1(n2139), .A2(n2138), .ZN(n2203) );
  INV_X1 U2125 ( .A(n2203), .ZN(n2270) );
  NAND2_X1 U2126 ( .A1(n2139), .A2(n2138), .ZN(n2269) );
  INV_X1 U2127 ( .A(n2269), .ZN(n2140) );
  AOI21_X1 U2128 ( .B1(n6127), .B2(n2270), .A(n2140), .ZN(n2202) );
  FA_X1 U2129 ( .A(n2143), .B(n2142), .CI(n2141), .CO(n2263), .S(n2195) );
  FA_X1 U2130 ( .A(n2146), .B(n2145), .CI(n2144), .CO(n2260), .S(n2192) );
  XNOR2_X1 U2131 ( .A(n5083), .B(n2147), .ZN(n2232) );
  OAI22_X1 U2132 ( .A1(n2232), .A2(n6128), .B1(n6130), .B2(n2148), .ZN(n2241)
         );
  XNOR2_X1 U2133 ( .A(n5085), .B(n28), .ZN(n2245) );
  OAI22_X1 U2134 ( .A1(n2245), .A2(n2246), .B1(n2149), .B2(n2247), .ZN(n2240)
         );
  XNOR2_X1 U2135 ( .A(n4683), .B(n4780), .ZN(n2228) );
  OAI22_X1 U2136 ( .A1(n4732), .A2(n2150), .B1(n2228), .B2(n4731), .ZN(n2239)
         );
  XNOR2_X1 U2137 ( .A(n4592), .B(n1803), .ZN(n2213) );
  OAI22_X1 U2138 ( .A1(n2151), .A2(n5124), .B1(n2213), .B2(n5123), .ZN(n2238)
         );
  XNOR2_X1 U2139 ( .A(n4673), .B(n30), .ZN(n2217) );
  OAI22_X1 U2140 ( .A1(n2152), .A2(n4830), .B1(n2217), .B2(n4829), .ZN(n2237)
         );
  XNOR2_X1 U2141 ( .A(n2153), .B(n15), .ZN(n2154) );
  NOR2_X1 U2142 ( .A1(n2154), .A2(n5109), .ZN(n2236) );
  FA_X1 U2143 ( .A(n2157), .B(n2156), .CI(n2155), .CO(n2252), .S(n2146) );
  FA_X1 U2144 ( .A(n2160), .B(n2159), .CI(n2158), .CO(n2211), .S(n2190) );
  INV_X1 U2145 ( .A(n2163), .ZN(n2221) );
  XNOR2_X1 U2146 ( .A(n5078), .B(n4587), .ZN(n2225) );
  OAI22_X1 U2147 ( .A1(n4661), .A2(n2161), .B1(n4660), .B2(n2225), .ZN(n2220)
         );
  FA_X1 U2148 ( .A(n2164), .B(n2163), .CI(n2162), .CO(n2219), .S(n2160) );
  FA_X1 U2149 ( .A(n2167), .B(n2166), .CI(n2165), .CO(n2209), .S(n2191) );
  XNOR2_X1 U2150 ( .A(n5076), .B(n1307), .ZN(n2235) );
  OAI22_X1 U2151 ( .A1(n2168), .A2(n4630), .B1(n2235), .B2(n4629), .ZN(n2244)
         );
  INV_X1 U2152 ( .A(dot_op_c_i[22]), .ZN(n4083) );
  OAI21_X1 U2153 ( .B1(n1661), .B2(n4083), .A(n5114), .ZN(n2243) );
  INV_X1 U2154 ( .A(n2169), .ZN(n2170) );
  NOR2_X1 U2155 ( .A1(n2170), .A2(n5116), .ZN(n2242) );
  FA_X1 U2156 ( .A(n2173), .B(n2172), .CI(n2171), .CO(n2230), .S(n2187) );
  XNOR2_X1 U2157 ( .A(n4590), .B(n17), .ZN(n2216) );
  OAI22_X1 U2158 ( .A1(n5113), .A2(n2174), .B1(n2216), .B2(n6114), .ZN(n2251)
         );
  XNOR2_X1 U2159 ( .A(n4795), .B(n4679), .ZN(n2212) );
  OAI22_X1 U2160 ( .A1(n2175), .A2(n4746), .B1(n2212), .B2(n4745), .ZN(n2250)
         );
  XNOR2_X1 U2161 ( .A(n4681), .B(n6111), .ZN(n2218) );
  OAI22_X1 U2162 ( .A1(n6125), .A2(n2176), .B1(n6123), .B2(n2218), .ZN(n2249)
         );
  FA_X1 U2163 ( .A(n2179), .B(n2178), .CI(n2177), .CO(n2224), .S(n2166) );
  FA_X1 U2164 ( .A(n2182), .B(n2181), .CI(n2180), .CO(n2223), .S(n2167) );
  FA_X1 U2165 ( .A(n2185), .B(n2184), .CI(n2183), .CO(n2222), .S(n2165) );
  FA_X1 U2166 ( .A(n2188), .B(n2187), .CI(n2186), .CO(n2255), .S(n2193) );
  FA_X1 U2167 ( .A(n2191), .B(n2190), .CI(n2189), .CO(n2207), .S(n2143) );
  FA_X1 U2168 ( .A(n2194), .B(n2193), .CI(n2192), .CO(n2206), .S(n2196) );
  FA_X1 U2169 ( .A(n2197), .B(n2196), .CI(n2195), .CO(n2198), .S(n2139) );
  NOR2_X1 U2170 ( .A1(n2199), .A2(n2198), .ZN(n2205) );
  INV_X1 U2171 ( .A(n2205), .ZN(n2200) );
  NAND2_X1 U2172 ( .A1(n2199), .A2(n2198), .ZN(n2204) );
  NAND2_X1 U2173 ( .A1(n2200), .A2(n2204), .ZN(n2201) );
  XOR2_X1 U2174 ( .A(n2202), .B(n2201), .Z(n5588) );
  NOR2_X1 U2175 ( .A1(n2203), .A2(n2205), .ZN(n5024) );
  OAI21_X1 U2176 ( .B1(n2205), .B2(n2269), .A(n2204), .ZN(n5026) );
  AOI21_X1 U2177 ( .B1(n6127), .B2(n5024), .A(n5026), .ZN(n2268) );
  FA_X1 U2178 ( .A(n2208), .B(n2207), .CI(n2206), .CO(n4621), .S(n2261) );
  FA_X1 U2179 ( .A(n2211), .B(n2210), .CI(n2209), .CO(n4618), .S(n2258) );
  XNOR2_X1 U2180 ( .A(n4839), .B(n4679), .ZN(n4579) );
  OAI22_X1 U2181 ( .A1(n2212), .A2(n4746), .B1(n4579), .B2(n4745), .ZN(n4606)
         );
  XNOR2_X1 U2182 ( .A(n4655), .B(n1803), .ZN(n4580) );
  OAI22_X1 U2183 ( .A1(n2213), .A2(n5124), .B1(n4580), .B2(n5123), .ZN(n4605)
         );
  INV_X1 U2184 ( .A(n2214), .ZN(n2215) );
  NOR2_X1 U2185 ( .A1(n2215), .A2(n5116), .ZN(n4604) );
  XNOR2_X1 U2186 ( .A(n4657), .B(n17), .ZN(n4584) );
  OAI22_X1 U2187 ( .A1(n5113), .A2(n2216), .B1(n4584), .B2(n6114), .ZN(n4600)
         );
  XNOR2_X1 U2188 ( .A(n4742), .B(n30), .ZN(n4585) );
  OAI22_X1 U2189 ( .A1(n2217), .A2(n4830), .B1(n4585), .B2(n4829), .ZN(n4599)
         );
  XNOR2_X1 U2190 ( .A(n4740), .B(n6111), .ZN(n4586) );
  OAI22_X1 U2191 ( .A1(n6125), .A2(n2218), .B1(n6123), .B2(n4586), .ZN(n4598)
         );
  FA_X1 U2192 ( .A(n2221), .B(n2220), .CI(n2219), .CO(n4610), .S(n2210) );
  FA_X1 U2193 ( .A(n2224), .B(n2223), .CI(n2222), .CO(n4578), .S(n2256) );
  XNOR2_X1 U2194 ( .A(n5107), .B(n1128), .ZN(n4588) );
  OAI22_X1 U2195 ( .A1(n4661), .A2(n2225), .B1(n4660), .B2(n4588), .ZN(n4583)
         );
  XNOR2_X1 U2196 ( .A(n2226), .B(n15), .ZN(n2227) );
  NOR2_X1 U2197 ( .A1(n2227), .A2(n5109), .ZN(n4582) );
  XNOR2_X1 U2198 ( .A(n4683), .B(n4841), .ZN(n4589) );
  OAI22_X1 U2199 ( .A1(n4732), .A2(n2228), .B1(n4589), .B2(n4731), .ZN(n4581)
         );
  FA_X1 U2200 ( .A(n2231), .B(n2230), .CI(n2229), .CO(n4576), .S(n2257) );
  INV_X1 U2201 ( .A(dot_op_c_i[23]), .ZN(n4226) );
  OAI21_X1 U2202 ( .B1(n1661), .B2(n4226), .A(n5114), .ZN(n4603) );
  AOI21_X1 U2203 ( .B1(n6130), .B2(n6128), .A(n2232), .ZN(n4602) );
  XNOR2_X1 U2204 ( .A(n5115), .B(n1307), .ZN(n4594) );
  OAI22_X1 U2205 ( .A1(n2235), .A2(n4630), .B1(n4594), .B2(n4629), .ZN(n4601)
         );
  FA_X1 U2206 ( .A(n2238), .B(n2237), .CI(n2236), .CO(n4608), .S(n2253) );
  FA_X1 U2207 ( .A(n2241), .B(n2240), .CI(n2239), .CO(n4607), .S(n2254) );
  FA_X1 U2208 ( .A(n2244), .B(n2243), .CI(n2242), .CO(n4597), .S(n2231) );
  AOI21_X1 U2209 ( .B1(n2247), .B2(n2246), .A(n2245), .ZN(n2248) );
  INV_X1 U2210 ( .A(n2248), .ZN(n4596) );
  FA_X1 U2211 ( .A(n2251), .B(n2250), .CI(n2249), .CO(n4595), .S(n2229) );
  FA_X1 U2212 ( .A(n2254), .B(n2253), .CI(n2252), .CO(n4613), .S(n2259) );
  FA_X1 U2213 ( .A(n2257), .B(n2256), .CI(n2255), .CO(n4574), .S(n2208) );
  FA_X1 U2214 ( .A(n2260), .B(n2259), .CI(n2258), .CO(n4573), .S(n2262) );
  FA_X1 U2215 ( .A(n2263), .B(n2262), .CI(n2261), .CO(n2264), .S(n2199) );
  NOR2_X1 U2216 ( .A1(n2265), .A2(n2264), .ZN(n5028) );
  INV_X1 U2217 ( .A(n5028), .ZN(n2266) );
  NAND2_X1 U2218 ( .A1(n2265), .A2(n2264), .ZN(n5027) );
  NAND2_X1 U2219 ( .A1(n2266), .A2(n5027), .ZN(n2267) );
  XOR2_X1 U2220 ( .A(n2268), .B(n2267), .Z(n5602) );
  AND2_X1 U2221 ( .A1(clpx_shift_i[0]), .A2(clpx_shift_i[1]), .ZN(n5490) );
  INV_X1 U2222 ( .A(n5490), .ZN(n5192) );
  NAND2_X1 U2223 ( .A1(n2270), .A2(n2269), .ZN(n2271) );
  XNOR2_X1 U2224 ( .A(n5032), .B(n2271), .ZN(n5573) );
  INV_X1 U2225 ( .A(clpx_shift_i[0]), .ZN(n2272) );
  INV_X1 U2226 ( .A(n2273), .ZN(n4911) );
  INV_X1 U2227 ( .A(n2774), .ZN(n2274) );
  NOR2_X1 U2228 ( .A1(n2274), .A2(n2775), .ZN(n2277) );
  INV_X1 U2229 ( .A(n2773), .ZN(n2275) );
  OAI21_X1 U2230 ( .B1(n2275), .B2(n2775), .A(n2776), .ZN(n2276) );
  AOI21_X1 U2231 ( .B1(n4911), .B2(n2277), .A(n2276), .ZN(n2282) );
  INV_X1 U2232 ( .A(n2278), .ZN(n2280) );
  NAND2_X1 U2233 ( .A1(n2280), .A2(n2279), .ZN(n2281) );
  XOR2_X1 U2234 ( .A(n2282), .B(n2281), .Z(n5183) );
  AOI22_X1 U2235 ( .A1(n5573), .A2(n5519), .B1(n5521), .B2(n5183), .ZN(n2283)
         );
  NOR2_X1 U2236 ( .A1(n2284), .A2(operator_i[1]), .ZN(n2659) );
  INV_X1 U2237 ( .A(n2659), .ZN(n2285) );
  INV_X1 U2238 ( .A(n38), .ZN(n5894) );
  AND2_X1 U2239 ( .A1(n2287), .A2(n2286), .ZN(n5622) );
  NAND2_X1 U2240 ( .A1(n5622), .A2(n2288), .ZN(n2347) );
  NOR2_X1 U2241 ( .A1(n2347), .A2(n2716), .ZN(n5158) );
  NAND2_X1 U2242 ( .A1(n2290), .A2(n2289), .ZN(n2291) );
  XNOR2_X1 U2243 ( .A(n2292), .B(n2291), .ZN(n5007) );
  NAND2_X1 U2244 ( .A1(n5007), .A2(n5008), .ZN(n2320) );
  INV_X1 U2245 ( .A(n2304), .ZN(n2293) );
  NOR2_X1 U2246 ( .A1(n2293), .A2(n2305), .ZN(n2297) );
  INV_X1 U2247 ( .A(n2294), .ZN(n2324) );
  INV_X1 U2248 ( .A(n2303), .ZN(n2295) );
  OAI21_X1 U2249 ( .B1(n2295), .B2(n2305), .A(n2306), .ZN(n2296) );
  AOI21_X1 U2250 ( .B1(n2297), .B2(n2324), .A(n2296), .ZN(n2302) );
  INV_X1 U2251 ( .A(n2298), .ZN(n2300) );
  NAND2_X1 U2252 ( .A1(n2300), .A2(n2299), .ZN(n2301) );
  XOR2_X1 U2253 ( .A(n2302), .B(n2301), .Z(n5011) );
  NAND2_X1 U2254 ( .A1(n5011), .A2(n5331), .ZN(n2319) );
  AOI21_X1 U2255 ( .B1(n2324), .B2(n2304), .A(n2303), .ZN(n2309) );
  INV_X1 U2256 ( .A(n2305), .ZN(n2307) );
  NAND2_X1 U2257 ( .A1(n2307), .A2(n2306), .ZN(n2308) );
  XOR2_X1 U2258 ( .A(n2309), .B(n2308), .Z(n5010) );
  NAND2_X1 U2259 ( .A1(n5010), .A2(n5304), .ZN(n2318) );
  INV_X1 U2260 ( .A(n2310), .ZN(n2322) );
  INV_X1 U2261 ( .A(n2321), .ZN(n2311) );
  AOI21_X1 U2262 ( .B1(n2324), .B2(n2322), .A(n2311), .ZN(n2316) );
  INV_X1 U2263 ( .A(n2312), .ZN(n2314) );
  NAND2_X1 U2264 ( .A1(n2314), .A2(n2313), .ZN(n2315) );
  XOR2_X1 U2265 ( .A(n2316), .B(n2315), .Z(n4985) );
  NAND2_X1 U2266 ( .A1(n4985), .A2(n5302), .ZN(n2317) );
  NAND4_X1 U2267 ( .A1(n2320), .A2(n2319), .A3(n2318), .A4(n2317), .ZN(n5507)
         );
  NAND2_X1 U2268 ( .A1(n2322), .A2(n2321), .ZN(n2323) );
  XNOR2_X1 U2269 ( .A(n2324), .B(n2323), .ZN(n4991) );
  INV_X1 U2270 ( .A(n2325), .ZN(n2341) );
  OAI21_X1 U2271 ( .B1(n2341), .B2(n2327), .A(n2326), .ZN(n2332) );
  INV_X1 U2272 ( .A(n2328), .ZN(n2330) );
  NAND2_X1 U2273 ( .A1(n2330), .A2(n2329), .ZN(n2331) );
  XNOR2_X1 U2274 ( .A(n2332), .B(n2331), .ZN(n4986) );
  NAND2_X1 U2275 ( .A1(n4986), .A2(n5331), .ZN(n2344) );
  OAI21_X1 U2276 ( .B1(n2341), .B2(n2333), .A(n2338), .ZN(n2337) );
  NAND2_X1 U2277 ( .A1(n2335), .A2(n2334), .ZN(n2336) );
  XNOR2_X1 U2278 ( .A(n2337), .B(n2336), .ZN(n4987) );
  NAND2_X1 U2279 ( .A1(n4987), .A2(n5304), .ZN(n2343) );
  NAND2_X1 U2280 ( .A1(n2339), .A2(n2338), .ZN(n2340) );
  XOR2_X1 U2281 ( .A(n2341), .B(n2340), .Z(n4999) );
  NAND2_X1 U2282 ( .A1(n4999), .A2(n5302), .ZN(n2342) );
  NAND3_X1 U2283 ( .A1(n2344), .A2(n2343), .A3(n2342), .ZN(n2345) );
  AOI21_X1 U2284 ( .B1(n5008), .B2(n4991), .A(n2345), .ZN(n5510) );
  INV_X1 U2285 ( .A(n2716), .ZN(n2346) );
  NOR2_X1 U2286 ( .A1(n2347), .A2(n2346), .ZN(n5529) );
  INV_X1 U2287 ( .A(n5529), .ZN(n5400) );
  NAND2_X1 U2288 ( .A1(n5622), .A2(n2830), .ZN(n2348) );
  NOR2_X1 U2289 ( .A1(n2348), .A2(n2716), .ZN(n5540) );
  INV_X1 U2290 ( .A(n2349), .ZN(n2368) );
  INV_X1 U2291 ( .A(n2350), .ZN(n2358) );
  INV_X1 U2292 ( .A(n2357), .ZN(n2351) );
  AOI21_X1 U2293 ( .B1(n2368), .B2(n2358), .A(n2351), .ZN(n2356) );
  INV_X1 U2294 ( .A(n2352), .ZN(n2354) );
  NAND2_X1 U2295 ( .A1(n2354), .A2(n2353), .ZN(n2355) );
  XOR2_X1 U2296 ( .A(n2356), .B(n2355), .Z(n5001) );
  INV_X1 U2297 ( .A(n5001), .ZN(n2375) );
  INV_X1 U2298 ( .A(n5331), .ZN(n5307) );
  NAND2_X1 U2299 ( .A1(n2358), .A2(n2357), .ZN(n2359) );
  XNOR2_X1 U2300 ( .A(n2368), .B(n2359), .ZN(n5000) );
  INV_X1 U2301 ( .A(n2360), .ZN(n2380) );
  OAI21_X1 U2302 ( .B1(n2380), .B2(n2376), .A(n2377), .ZN(n2365) );
  INV_X1 U2303 ( .A(n2361), .ZN(n2363) );
  NAND2_X1 U2304 ( .A1(n2363), .A2(n2362), .ZN(n2364) );
  XNOR2_X1 U2305 ( .A(n2365), .B(n2364), .ZN(n5310) );
  AOI22_X1 U2306 ( .A1(n5000), .A2(n5304), .B1(n5310), .B2(n5302), .ZN(n2374)
         );
  AOI21_X1 U2307 ( .B1(n2368), .B2(n2367), .A(n2366), .ZN(n2372) );
  NAND2_X1 U2308 ( .A1(n2370), .A2(n2369), .ZN(n2371) );
  XOR2_X1 U2309 ( .A(n2372), .B(n2371), .Z(n4998) );
  NAND2_X1 U2310 ( .A1(n4998), .A2(n5008), .ZN(n2373) );
  OAI211_X1 U2311 ( .C1(n2375), .C2(n5307), .A(n2374), .B(n2373), .ZN(n5418)
         );
  INV_X1 U2312 ( .A(n2376), .ZN(n2378) );
  NAND2_X1 U2313 ( .A1(n2378), .A2(n2377), .ZN(n2379) );
  XOR2_X1 U2314 ( .A(n2380), .B(n2379), .Z(n5301) );
  NAND2_X1 U2315 ( .A1(n2382), .A2(n2381), .ZN(n2386) );
  INV_X1 U2316 ( .A(n2383), .ZN(n2389) );
  AOI21_X1 U2317 ( .B1(n2389), .B2(n2388), .A(n2384), .ZN(n2385) );
  XOR2_X1 U2318 ( .A(n2386), .B(n2385), .Z(n5305) );
  INV_X1 U2319 ( .A(n5305), .ZN(n2396) );
  NAND2_X1 U2320 ( .A1(n2388), .A2(n2387), .ZN(n2390) );
  XNOR2_X1 U2321 ( .A(n2390), .B(n2389), .ZN(n5303) );
  NAND2_X1 U2322 ( .A1(n2392), .A2(n2391), .ZN(n2393) );
  XNOR2_X1 U2323 ( .A(n2394), .B(n2393), .ZN(n5335) );
  AOI22_X1 U2324 ( .A1(n5303), .A2(n5304), .B1(n5302), .B2(n5335), .ZN(n2395)
         );
  OAI21_X1 U2325 ( .B1(n2396), .B2(n5307), .A(n2395), .ZN(n2397) );
  AOI21_X1 U2326 ( .B1(n5311), .B2(n5301), .A(n2397), .ZN(n5293) );
  NAND2_X1 U2327 ( .A1(n5622), .A2(n5384), .ZN(n6095) );
  NOR2_X1 U2328 ( .A1(operator_i[2]), .A2(operator_i[1]), .ZN(n2840) );
  NAND2_X1 U2329 ( .A1(n2840), .A2(operator_i[0]), .ZN(n2866) );
  XNOR2_X1 U2330 ( .A(n2879), .B(op_a_i[0]), .ZN(n2621) );
  XNOR2_X1 U2331 ( .A(n6116), .B(n25), .ZN(n2399) );
  XOR2_X1 U2332 ( .A(op_b_i[4]), .B(n25), .Z(n2398) );
  INV_X1 U2333 ( .A(n2472), .ZN(n5811) );
  XOR2_X1 U2334 ( .A(op_b_i[4]), .B(n5811), .Z(n2865) );
  INV_X1 U2335 ( .A(n2865), .ZN(n6010) );
  XNOR2_X1 U2336 ( .A(n6002), .B(n25), .ZN(n3942) );
  INV_X1 U2337 ( .A(n2865), .ZN(n5809) );
  OAI22_X1 U2338 ( .A1(n2399), .A2(n2867), .B1(n3942), .B2(n5809), .ZN(n3965)
         );
  OR2_X1 U2339 ( .A1(n6116), .A2(n2442), .ZN(n2400) );
  OAI22_X1 U2340 ( .A1(n2400), .A2(n6010), .B1(n2867), .B2(n2442), .ZN(n3964)
         );
  INV_X1 U2341 ( .A(n2527), .ZN(n5985) );
  XNOR2_X1 U2342 ( .A(n22), .B(n5985), .ZN(n3899) );
  XNOR2_X1 U2343 ( .A(n55), .B(n5985), .ZN(n2475) );
  OAI22_X1 U2344 ( .A1(n3899), .A2(n5635), .B1(n2475), .B2(n3241), .ZN(n3940)
         );
  XNOR2_X1 U2345 ( .A(n2879), .B(op_a_i[3]), .ZN(n5976) );
  INV_X1 U2346 ( .A(n2472), .ZN(n6015) );
  XNOR2_X1 U2347 ( .A(n56), .B(n6015), .ZN(n3902) );
  INV_X1 U2348 ( .A(n2527), .ZN(n5856) );
  XNOR2_X1 U2349 ( .A(op_b_i[2]), .B(n5856), .ZN(n2401) );
  INV_X1 U2350 ( .A(n2401), .ZN(n4137) );
  XNOR2_X1 U2351 ( .A(n5848), .B(n6015), .ZN(n2476) );
  XOR2_X1 U2352 ( .A(op_b_i[2]), .B(n4342), .Z(n2402) );
  OAI22_X1 U2353 ( .A1(n3902), .A2(n10), .B1(n2476), .B2(n2585), .ZN(n3939) );
  XNOR2_X1 U2354 ( .A(dot_op_b_i[20]), .B(dot_op_b_i[19]), .ZN(n3719) );
  INV_X1 U2355 ( .A(n59), .ZN(n2403) );
  AND2_X1 U2356 ( .A1(dot_op_a_i[16]), .A2(n2403), .ZN(n2412) );
  INV_X1 U2357 ( .A(n3715), .ZN(n2404) );
  AND2_X1 U2358 ( .A1(dot_op_a_i[24]), .A2(n2404), .ZN(n2411) );
  NAND2_X1 U2359 ( .A1(dot_op_b_i[17]), .A2(n1662), .ZN(n3479) );
  XNOR2_X1 U2360 ( .A(dot_op_b_i[17]), .B(dot_op_a_i[19]), .ZN(n2481) );
  XNOR2_X1 U2361 ( .A(dot_op_b_i[17]), .B(dot_op_a_i[20]), .ZN(n2413) );
  OAI22_X1 U2362 ( .A1(n3479), .A2(n2481), .B1(n2413), .B2(n1662), .ZN(n2574)
         );
  XOR2_X1 U2363 ( .A(dot_op_b_i[26]), .B(dot_op_b_i[27]), .Z(n2405) );
  OR2_X1 U2364 ( .A1(dot_op_a_i[24]), .A2(n1226), .ZN(n2406) );
  OAI22_X1 U2365 ( .A1(n3713), .A2(n1226), .B1(n2406), .B2(n3711), .ZN(n2492)
         );
  XNOR2_X1 U2366 ( .A(dot_op_b_i[27]), .B(dot_op_a_i[24]), .ZN(n2407) );
  XNOR2_X1 U2367 ( .A(dot_op_b_i[27]), .B(dot_op_a_i[25]), .ZN(n2415) );
  OAI22_X1 U2368 ( .A1(n3713), .A2(n2407), .B1(n3711), .B2(n2415), .ZN(n2491)
         );
  NAND2_X1 U2369 ( .A1(dot_op_b_i[25]), .A2(n1312), .ZN(n3482) );
  XNOR2_X1 U2370 ( .A(dot_op_b_i[25]), .B(dot_op_a_i[26]), .ZN(n2484) );
  XNOR2_X1 U2371 ( .A(dot_op_b_i[25]), .B(dot_op_a_i[27]), .ZN(n2417) );
  OAI22_X1 U2372 ( .A1(n3482), .A2(n2484), .B1(n2417), .B2(n1312), .ZN(n2490)
         );
  XOR2_X1 U2373 ( .A(dot_op_b_i[20]), .B(dot_op_b_i[21]), .Z(n2408) );
  NAND2_X1 U2374 ( .A1(n2408), .A2(n3719), .ZN(n3721) );
  XNOR2_X1 U2375 ( .A(dot_op_b_i[21]), .B(dot_op_a_i[16]), .ZN(n2409) );
  XNOR2_X1 U2376 ( .A(dot_op_b_i[21]), .B(dot_op_a_i[17]), .ZN(n3720) );
  OAI22_X1 U2377 ( .A1(n3721), .A2(n2409), .B1(n59), .B2(n3720), .ZN(n3916) );
  XOR2_X1 U2378 ( .A(dot_op_b_i[18]), .B(dot_op_b_i[19]), .Z(n2410) );
  XNOR2_X1 U2379 ( .A(dot_op_b_i[18]), .B(dot_op_b_i[17]), .ZN(n3463) );
  NAND2_X1 U2380 ( .A1(n2410), .A2(n3463), .ZN(n3465) );
  XNOR2_X1 U2381 ( .A(dot_op_b_i[19]), .B(dot_op_a_i[18]), .ZN(n2418) );
  XNOR2_X1 U2382 ( .A(dot_op_b_i[19]), .B(dot_op_a_i[19]), .ZN(n3416) );
  OAI22_X1 U2383 ( .A1(n3465), .A2(n2418), .B1(n60), .B2(n3416), .ZN(n3915) );
  HA_X1 U2384 ( .A(n2412), .B(n2411), .CO(n3914), .S(n2575) );
  XNOR2_X1 U2385 ( .A(dot_op_b_i[25]), .B(dot_op_a_i[28]), .ZN(n2416) );
  XNOR2_X1 U2386 ( .A(dot_op_b_i[25]), .B(dot_op_a_i[29]), .ZN(n3415) );
  OAI22_X1 U2387 ( .A1(n3482), .A2(n2416), .B1(n3415), .B2(n1312), .ZN(n3846)
         );
  XNOR2_X1 U2388 ( .A(dot_op_b_i[17]), .B(dot_op_a_i[21]), .ZN(n3414) );
  OAI22_X1 U2389 ( .A1(n3479), .A2(n2413), .B1(n3414), .B2(n1662), .ZN(n3845)
         );
  OR2_X1 U2390 ( .A1(dot_op_a_i[16]), .A2(n1547), .ZN(n2414) );
  OAI22_X1 U2391 ( .A1(n3721), .A2(n1547), .B1(n2414), .B2(n59), .ZN(n3844) );
  XNOR2_X1 U2392 ( .A(dot_op_b_i[27]), .B(dot_op_a_i[26]), .ZN(n2422) );
  OAI22_X1 U2393 ( .A1(n3713), .A2(n2415), .B1(n3711), .B2(n2422), .ZN(n2479)
         );
  OAI22_X1 U2394 ( .A1(n3482), .A2(n2417), .B1(n2416), .B2(n1312), .ZN(n2478)
         );
  XNOR2_X1 U2395 ( .A(dot_op_b_i[19]), .B(dot_op_a_i[17]), .ZN(n2482) );
  OAI22_X1 U2396 ( .A1(n3465), .A2(n2482), .B1(n60), .B2(n2418), .ZN(n2477) );
  XOR2_X1 U2397 ( .A(dot_op_b_i[28]), .B(dot_op_b_i[29]), .Z(n2419) );
  OR2_X1 U2398 ( .A1(dot_op_a_i[24]), .A2(n1239), .ZN(n2420) );
  OAI22_X1 U2399 ( .A1(n3717), .A2(n1239), .B1(n2420), .B2(n3715), .ZN(n3841)
         );
  XNOR2_X1 U2400 ( .A(dot_op_b_i[29]), .B(dot_op_a_i[24]), .ZN(n2421) );
  XNOR2_X1 U2401 ( .A(dot_op_b_i[29]), .B(dot_op_a_i[25]), .ZN(n3716) );
  OAI22_X1 U2402 ( .A1(n3717), .A2(n2421), .B1(n3715), .B2(n3716), .ZN(n3840)
         );
  XNOR2_X1 U2403 ( .A(dot_op_b_i[27]), .B(dot_op_a_i[27]), .ZN(n3712) );
  OAI22_X1 U2404 ( .A1(n3713), .A2(n2422), .B1(n3711), .B2(n3712), .ZN(n3839)
         );
  MUX2_X1 U2406 ( .A(n2424), .B(n2423), .S(n6143), .Z(n3962) );
  XOR2_X1 U2407 ( .A(dot_op_b_i[10]), .B(dot_op_b_i[11]), .Z(n2425) );
  NAND2_X1 U2408 ( .A1(n2425), .A2(n3493), .ZN(n3496) );
  XNOR2_X1 U2409 ( .A(dot_op_a_i[9]), .B(dot_op_b_i[11]), .ZN(n2438) );
  XNOR2_X1 U2410 ( .A(dot_op_b_i[11]), .B(dot_op_a_i[10]), .ZN(n2557) );
  OAI22_X1 U2411 ( .A1(n3496), .A2(n2438), .B1(n3493), .B2(n2557), .ZN(n2552)
         );
  INV_X1 U2412 ( .A(dot_op_b_i[8]), .ZN(n3544) );
  NAND2_X1 U2413 ( .A1(dot_op_b_i[9]), .A2(n3544), .ZN(n3547) );
  XNOR2_X1 U2414 ( .A(dot_op_a_i[11]), .B(dot_op_b_i[9]), .ZN(n2440) );
  XNOR2_X1 U2415 ( .A(dot_op_b_i[9]), .B(dot_op_a_i[12]), .ZN(n2546) );
  OAI22_X1 U2416 ( .A1(n3547), .A2(n2440), .B1(n2546), .B2(n3544), .ZN(n2551)
         );
  XOR2_X1 U2417 ( .A(dot_op_b_i[2]), .B(dot_op_b_i[3]), .Z(n2426) );
  NAND2_X1 U2418 ( .A1(n2426), .A2(n3549), .ZN(n3551) );
  XNOR2_X1 U2419 ( .A(dot_op_a_i[1]), .B(dot_op_b_i[3]), .ZN(n2429) );
  XNOR2_X1 U2420 ( .A(dot_op_b_i[3]), .B(dot_op_a_i[2]), .ZN(n2543) );
  OAI22_X1 U2421 ( .A1(n3551), .A2(n2429), .B1(n3549), .B2(n2543), .ZN(n2550)
         );
  INV_X1 U2422 ( .A(dot_op_b_i[3]), .ZN(n2428) );
  OR2_X1 U2423 ( .A1(dot_op_a_i[0]), .A2(n2428), .ZN(n2427) );
  OAI22_X1 U2424 ( .A1(n3551), .A2(n2428), .B1(n2427), .B2(n3549), .ZN(n2471)
         );
  INV_X1 U2425 ( .A(dot_op_b_i[0]), .ZN(n3540) );
  NAND2_X1 U2426 ( .A1(dot_op_b_i[1]), .A2(n3540), .ZN(n3543) );
  XNOR2_X1 U2427 ( .A(dot_op_b_i[1]), .B(dot_op_a_i[2]), .ZN(n2431) );
  XNOR2_X1 U2428 ( .A(dot_op_a_i[3]), .B(dot_op_b_i[1]), .ZN(n2449) );
  OAI22_X1 U2429 ( .A1(n3543), .A2(n2431), .B1(n2449), .B2(n3540), .ZN(n2470)
         );
  XNOR2_X1 U2430 ( .A(dot_op_b_i[3]), .B(dot_op_a_i[0]), .ZN(n2430) );
  OAI22_X1 U2431 ( .A1(n3551), .A2(n2430), .B1(n2429), .B2(n3549), .ZN(n2469)
         );
  XNOR2_X1 U2432 ( .A(dot_op_a_i[9]), .B(dot_op_b_i[9]), .ZN(n2459) );
  XNOR2_X1 U2433 ( .A(dot_op_b_i[9]), .B(dot_op_a_i[10]), .ZN(n2441) );
  OAI22_X1 U2434 ( .A1(n3547), .A2(n2459), .B1(n2441), .B2(n3544), .ZN(n2534)
         );
  XNOR2_X1 U2435 ( .A(dot_op_a_i[1]), .B(dot_op_b_i[1]), .ZN(n2458) );
  OAI22_X1 U2436 ( .A1(n3543), .A2(n2458), .B1(n2431), .B2(n3540), .ZN(n2533)
         );
  INV_X1 U2437 ( .A(n3549), .ZN(n2432) );
  AND2_X1 U2438 ( .A1(dot_op_a_i[0]), .A2(n2432), .ZN(n2435) );
  INV_X1 U2439 ( .A(n3493), .ZN(n2433) );
  AND2_X1 U2440 ( .A1(dot_op_a_i[8]), .A2(n2433), .ZN(n2434) );
  HA_X1 U2441 ( .A(n2435), .B(n2434), .CO(n2582), .S(n2532) );
  INV_X1 U2442 ( .A(dot_op_b_i[11]), .ZN(n2437) );
  OR2_X1 U2443 ( .A1(dot_op_a_i[8]), .A2(n2437), .ZN(n2436) );
  OAI22_X1 U2444 ( .A1(n3496), .A2(n2437), .B1(n2436), .B2(n3493), .ZN(n2452)
         );
  XNOR2_X1 U2445 ( .A(dot_op_b_i[11]), .B(dot_op_a_i[8]), .ZN(n2439) );
  OAI22_X1 U2446 ( .A1(n3496), .A2(n2439), .B1(n2438), .B2(n3493), .ZN(n2451)
         );
  OAI22_X1 U2447 ( .A1(n3547), .A2(n2441), .B1(n2440), .B2(n3544), .ZN(n2450)
         );
  INV_X1 U2448 ( .A(op_b_i[5]), .ZN(n2442) );
  NOR2_X1 U2449 ( .A1(n6119), .A2(n2442), .ZN(n2443) );
  MUX2_X1 U2450 ( .A(n2444), .B(n2443), .S(n29), .Z(n3973) );
  INV_X1 U2451 ( .A(op_c_i[5]), .ZN(n2445) );
  OAI22_X1 U2452 ( .A1(n6112), .A2(n2446), .B1(n2525), .B2(n2445), .ZN(n3972)
         );
  INV_X1 U2453 ( .A(n3536), .ZN(n2447) );
  AND2_X1 U2454 ( .A1(dot_op_a_i[0]), .A2(n2447), .ZN(n2545) );
  INV_X1 U2455 ( .A(n3511), .ZN(n2448) );
  AND2_X1 U2456 ( .A1(dot_op_a_i[8]), .A2(n2448), .ZN(n2544) );
  XNOR2_X1 U2457 ( .A(dot_op_b_i[1]), .B(dot_op_a_i[4]), .ZN(n2547) );
  OAI22_X1 U2458 ( .A1(n3543), .A2(n2449), .B1(n2547), .B2(n3540), .ZN(n2539)
         );
  FA_X1 U2459 ( .A(n2452), .B(n2451), .CI(n2450), .CO(n2538), .S(n2581) );
  INV_X1 U2460 ( .A(op_b_i[4]), .ZN(n2453) );
  NOR2_X1 U2461 ( .A1(n6118), .A2(n2453), .ZN(n2454) );
  MUX2_X1 U2462 ( .A(n2455), .B(n2454), .S(n29), .Z(n2497) );
  INV_X1 U2463 ( .A(op_c_i[4]), .ZN(n2456) );
  OAI22_X1 U2464 ( .A1(n6112), .A2(n2457), .B1(n2525), .B2(n2456), .ZN(n2496)
         );
  OAI22_X1 U2465 ( .A1(n3543), .A2(dot_op_a_i[0]), .B1(n2458), .B2(n3540), 
        .ZN(n2613) );
  OAI22_X1 U2466 ( .A1(n3547), .A2(dot_op_a_i[8]), .B1(n2459), .B2(n3544), 
        .ZN(n2612) );
  INV_X1 U2467 ( .A(dot_op_b_i[1]), .ZN(n2460) );
  OR2_X1 U2468 ( .A1(dot_op_a_i[0]), .A2(n2460), .ZN(n2461) );
  NAND2_X1 U2469 ( .A1(n2461), .A2(n3543), .ZN(n2611) );
  INV_X1 U2470 ( .A(op_b_i[2]), .ZN(n2462) );
  NOR2_X1 U2471 ( .A1(n6119), .A2(n2462), .ZN(n2463) );
  MUX2_X1 U2472 ( .A(n2464), .B(n2463), .S(n29), .Z(n2537) );
  INV_X1 U2473 ( .A(op_c_i[2]), .ZN(n2465) );
  OAI22_X1 U2474 ( .A1(n6112), .A2(n2466), .B1(n2525), .B2(n2465), .ZN(n2536)
         );
  INV_X1 U2475 ( .A(op_c_i[3]), .ZN(n2467) );
  OAI22_X1 U2476 ( .A1(n6112), .A2(n2468), .B1(n2525), .B2(n2467), .ZN(n2506)
         );
  FA_X1 U2477 ( .A(n2471), .B(n2470), .CI(n2469), .CO(n2568), .S(n2474) );
  INV_X1 U2478 ( .A(op_b_i[3]), .ZN(n2472) );
  NOR2_X1 U2479 ( .A1(n6119), .A2(n2472), .ZN(n2473) );
  MUX2_X1 U2480 ( .A(n2474), .B(n2473), .S(n29), .Z(n2505) );
  XNOR2_X1 U2481 ( .A(n56), .B(n5985), .ZN(n2499) );
  OAI22_X1 U2482 ( .A1(n2499), .A2(n3241), .B1(n2475), .B2(n5635), .ZN(n2561)
         );
  AND2_X1 U2483 ( .A1(n6116), .A2(n2865), .ZN(n2560) );
  XNOR2_X1 U2484 ( .A(n6002), .B(n6015), .ZN(n2586) );
  OAI22_X1 U2485 ( .A1(n2586), .A2(n2585), .B1(n2476), .B2(n10), .ZN(n2559) );
  FA_X1 U2486 ( .A(n2479), .B(n2478), .CI(n2477), .CO(n3947), .S(n2564) );
  OR2_X1 U2487 ( .A1(dot_op_a_i[16]), .A2(n1626), .ZN(n2480) );
  OAI22_X1 U2488 ( .A1(n3465), .A2(n1626), .B1(n2480), .B2(n60), .ZN(n2590) );
  XNOR2_X1 U2489 ( .A(dot_op_b_i[17]), .B(dot_op_a_i[18]), .ZN(n2485) );
  OAI22_X1 U2490 ( .A1(n3479), .A2(n2485), .B1(n2481), .B2(n1662), .ZN(n2589)
         );
  XNOR2_X1 U2491 ( .A(dot_op_b_i[19]), .B(dot_op_a_i[16]), .ZN(n2483) );
  OAI22_X1 U2492 ( .A1(n3465), .A2(n2483), .B1(n60), .B2(n2482), .ZN(n2588) );
  XNOR2_X1 U2493 ( .A(dot_op_b_i[25]), .B(dot_op_a_i[25]), .ZN(n2510) );
  OAI22_X1 U2494 ( .A1(n3482), .A2(n2510), .B1(n2484), .B2(n1312), .ZN(n2517)
         );
  XNOR2_X1 U2495 ( .A(dot_op_b_i[17]), .B(dot_op_a_i[17]), .ZN(n2509) );
  OAI22_X1 U2496 ( .A1(n3479), .A2(n2509), .B1(n2485), .B2(n1662), .ZN(n2516)
         );
  INV_X1 U2497 ( .A(n3463), .ZN(n2486) );
  AND2_X1 U2498 ( .A1(dot_op_a_i[16]), .A2(n2486), .ZN(n2489) );
  INV_X1 U2499 ( .A(n3711), .ZN(n2487) );
  AND2_X1 U2500 ( .A1(dot_op_a_i[24]), .A2(n2487), .ZN(n2488) );
  HA_X1 U2501 ( .A(n2489), .B(n2488), .CO(n2501), .S(n2515) );
  FA_X1 U2502 ( .A(n2492), .B(n2491), .CI(n2490), .CO(n2573), .S(n2500) );
  MUX2_X1 U2503 ( .A(n2494), .B(n2493), .S(n6117), .Z(n2598) );
  FA_X1 U2504 ( .A(n2497), .B(n2496), .CI(n2495), .CO(n3971), .S(n2597) );
  OR2_X1 U2505 ( .A1(n6116), .A2(n2472), .ZN(n2498) );
  OAI22_X1 U2506 ( .A1(n2498), .A2(n10), .B1(n2585), .B2(n2472), .ZN(n2572) );
  XNOR2_X1 U2507 ( .A(n5848), .B(n5985), .ZN(n2508) );
  OAI22_X1 U2508 ( .A1(n2499), .A2(n5635), .B1(n2508), .B2(n3241), .ZN(n2571)
         );
  FA_X1 U2509 ( .A(n2502), .B(n2501), .CI(n2500), .CO(n2562), .S(n2503) );
  MUX2_X1 U2510 ( .A(n2504), .B(n2503), .S(n6143), .Z(n2604) );
  FA_X1 U2511 ( .A(n2507), .B(n2506), .CI(n2505), .CO(n2495), .S(n2603) );
  XNOR2_X1 U2512 ( .A(n6002), .B(n5985), .ZN(n2622) );
  OAI22_X1 U2513 ( .A1(n2622), .A2(n3241), .B1(n2508), .B2(n5635), .ZN(n2514)
         );
  OAI22_X1 U2514 ( .A1(n3479), .A2(dot_op_a_i[16]), .B1(n2509), .B2(n1662), 
        .ZN(n2618) );
  OAI22_X1 U2515 ( .A1(n3482), .A2(dot_op_a_i[24]), .B1(n2510), .B2(n1312), 
        .ZN(n2617) );
  INV_X1 U2516 ( .A(dot_op_b_i[17]), .ZN(n2511) );
  OR2_X1 U2517 ( .A1(dot_op_a_i[16]), .A2(n2511), .ZN(n2512) );
  NAND2_X1 U2518 ( .A1(n2512), .A2(n3479), .ZN(n2616) );
  MUX2_X1 U2519 ( .A(n2514), .B(n2513), .S(n6142), .Z(n2639) );
  AND2_X1 U2520 ( .A1(n6116), .A2(n4137), .ZN(n2519) );
  FA_X1 U2521 ( .A(n2517), .B(n2516), .CI(n2515), .CO(n2502), .S(n2518) );
  MUX2_X1 U2522 ( .A(n2519), .B(n2518), .S(n6117), .Z(n2638) );
  AND2_X1 U2523 ( .A1(dot_op_a_i[16]), .A2(dot_op_b_i[16]), .ZN(n2520) );
  AND2_X1 U2524 ( .A1(n2520), .A2(n6140), .ZN(n2629) );
  AND2_X1 U2525 ( .A1(dot_op_a_i[0]), .A2(dot_op_b_i[0]), .ZN(n2521) );
  AND2_X1 U2526 ( .A1(n2521), .A2(n2591), .ZN(n2628) );
  INV_X1 U2527 ( .A(op_c_i[0]), .ZN(n2522) );
  OAI22_X1 U2528 ( .A1(n6112), .A2(n2523), .B1(n2525), .B2(n2522), .ZN(n2627)
         );
  INV_X1 U2529 ( .A(op_c_i[1]), .ZN(n2524) );
  OAI22_X1 U2530 ( .A1(n6112), .A2(n2526), .B1(n2525), .B2(n2524), .ZN(n2609)
         );
  INV_X1 U2531 ( .A(op_b_i[1]), .ZN(n2527) );
  NOR2_X1 U2532 ( .A1(n6119), .A2(n2527), .ZN(n2531) );
  INV_X1 U2533 ( .A(dot_op_b_i[9]), .ZN(n2528) );
  OR2_X1 U2534 ( .A1(dot_op_a_i[8]), .A2(n2528), .ZN(n2529) );
  NAND2_X1 U2535 ( .A1(n2529), .A2(n3547), .ZN(n2530) );
  MUX2_X1 U2536 ( .A(n2531), .B(n2530), .S(n6140), .Z(n2608) );
  FA_X1 U2537 ( .A(n2534), .B(n2533), .CI(n2532), .CO(n2583), .S(n2535) );
  AND2_X1 U2538 ( .A1(n2535), .A2(n6117), .ZN(n2579) );
  HA_X1 U2539 ( .A(n2537), .B(n2536), .CO(n2507), .S(n2578) );
  FA_X1 U2540 ( .A(n2540), .B(n2539), .CI(n2538), .CO(n3976), .S(n2455) );
  XOR2_X1 U2541 ( .A(dot_op_b_i[4]), .B(dot_op_b_i[5]), .Z(n2541) );
  NAND2_X1 U2542 ( .A1(n2541), .A2(n3536), .ZN(n3539) );
  XNOR2_X1 U2543 ( .A(dot_op_b_i[5]), .B(dot_op_a_i[0]), .ZN(n2542) );
  XNOR2_X1 U2544 ( .A(dot_op_a_i[1]), .B(dot_op_b_i[5]), .ZN(n3492) );
  OAI22_X1 U2545 ( .A1(n3539), .A2(n2542), .B1(n3492), .B2(n3536), .ZN(n3810)
         );
  XNOR2_X1 U2546 ( .A(dot_op_a_i[3]), .B(dot_op_b_i[3]), .ZN(n3550) );
  OAI22_X1 U2547 ( .A1(n3551), .A2(n2543), .B1(n3550), .B2(n3549), .ZN(n3809)
         );
  HA_X1 U2548 ( .A(n2545), .B(n2544), .CO(n3808), .S(n2540) );
  XNOR2_X1 U2549 ( .A(dot_op_a_i[13]), .B(dot_op_b_i[9]), .ZN(n3546) );
  OAI22_X1 U2550 ( .A1(n3547), .A2(n2546), .B1(n3546), .B2(n3544), .ZN(n3679)
         );
  XNOR2_X1 U2551 ( .A(dot_op_a_i[5]), .B(dot_op_b_i[1]), .ZN(n3542) );
  OAI22_X1 U2552 ( .A1(n3543), .A2(n2547), .B1(n3542), .B2(n3540), .ZN(n3678)
         );
  INV_X1 U2553 ( .A(dot_op_b_i[5]), .ZN(n2549) );
  OR2_X1 U2554 ( .A1(dot_op_a_i[0]), .A2(n2549), .ZN(n2548) );
  OAI22_X1 U2555 ( .A1(n3539), .A2(n2549), .B1(n2548), .B2(n3536), .ZN(n3677)
         );
  FA_X1 U2556 ( .A(n2552), .B(n2551), .CI(n2550), .CO(n3881), .S(n2569) );
  XOR2_X1 U2557 ( .A(dot_op_b_i[12]), .B(dot_op_b_i[13]), .Z(n2553) );
  INV_X1 U2558 ( .A(dot_op_b_i[13]), .ZN(n2555) );
  OR2_X1 U2559 ( .A1(dot_op_a_i[8]), .A2(n2555), .ZN(n2554) );
  OAI22_X1 U2560 ( .A1(n3514), .A2(n2555), .B1(n2554), .B2(n3511), .ZN(n3674)
         );
  XNOR2_X1 U2561 ( .A(dot_op_b_i[13]), .B(dot_op_a_i[8]), .ZN(n2556) );
  XNOR2_X1 U2562 ( .A(dot_op_a_i[9]), .B(dot_op_b_i[13]), .ZN(n3491) );
  OAI22_X1 U2563 ( .A1(n3514), .A2(n2556), .B1(n3491), .B2(n3511), .ZN(n3673)
         );
  XNOR2_X1 U2564 ( .A(dot_op_a_i[11]), .B(dot_op_b_i[11]), .ZN(n3490) );
  OAI22_X1 U2565 ( .A1(n3496), .A2(n2557), .B1(n3490), .B2(n3493), .ZN(n3672)
         );
  AND2_X1 U2566 ( .A1(n2558), .A2(n6145), .ZN(n3959) );
  FA_X1 U2567 ( .A(n2561), .B(n2560), .CI(n2559), .CO(n2566), .S(n2494) );
  FA_X1 U2568 ( .A(n2564), .B(n2563), .CI(n2562), .CO(n2565), .S(n2493) );
  MUX2_X1 U2569 ( .A(n2566), .B(n2565), .S(n6117), .Z(n3958) );
  FA_X1 U2570 ( .A(n2569), .B(n2568), .CI(n2567), .CO(n2444), .S(n2570) );
  AND2_X1 U2571 ( .A1(n2570), .A2(n6142), .ZN(n2601) );
  HA_X1 U2572 ( .A(n2572), .B(n2571), .CO(n2577), .S(n2504) );
  FA_X1 U2573 ( .A(n2575), .B(n2574), .CI(n2573), .CO(n3968), .S(n2576) );
  MUX2_X1 U2574 ( .A(n2577), .B(n2576), .S(n6141), .Z(n2600) );
  FA_X1 U2575 ( .A(n2580), .B(n2579), .CI(n2578), .CO(n2607), .S(n2637) );
  FA_X1 U2576 ( .A(n2583), .B(n2582), .CI(n2581), .CO(n2567), .S(n2584) );
  AND2_X1 U2577 ( .A1(n2584), .A2(n6142), .ZN(n2606) );
  XNOR2_X1 U2578 ( .A(n6116), .B(n6015), .ZN(n2587) );
  OAI22_X1 U2579 ( .A1(n2587), .A2(n2585), .B1(n2586), .B2(n10), .ZN(n2593) );
  FA_X1 U2580 ( .A(n2590), .B(n2589), .CI(n2588), .CO(n2563), .S(n2592) );
  MUX2_X1 U2581 ( .A(n2593), .B(n2592), .S(n6141), .Z(n2605) );
  OR2_X1 U2582 ( .A1(n2595), .A2(n2594), .ZN(n3989) );
  NAND2_X1 U2583 ( .A1(n2595), .A2(n2594), .ZN(n3986) );
  NAND2_X1 U2584 ( .A1(n3989), .A2(n3986), .ZN(n2651) );
  FA_X1 U2585 ( .A(n2598), .B(n2597), .CI(n2596), .CO(n3960), .S(n2650) );
  FA_X1 U2586 ( .A(n2601), .B(n2600), .CI(n2599), .CO(n3957), .S(n2649) );
  NOR2_X1 U2587 ( .A1(n2650), .A2(n2649), .ZN(n2805) );
  FA_X1 U2588 ( .A(n2604), .B(n2603), .CI(n2602), .CO(n2596), .S(n2647) );
  FA_X1 U2589 ( .A(n2607), .B(n2606), .CI(n2605), .CO(n2599), .S(n2646) );
  NOR2_X1 U2590 ( .A1(n2647), .A2(n2646), .ZN(n2753) );
  FA_X1 U2591 ( .A(n2610), .B(n2609), .CI(n2608), .CO(n2580), .S(n2642) );
  FA_X1 U2592 ( .A(n2613), .B(n2612), .CI(n2611), .CO(n2464), .S(n2614) );
  AND2_X1 U2593 ( .A1(n2614), .A2(n6142), .ZN(n2641) );
  OR2_X1 U2594 ( .A1(n6116), .A2(n2527), .ZN(n2615) );
  NAND2_X1 U2595 ( .A1(n3241), .A2(n2615), .ZN(n2620) );
  FA_X1 U2596 ( .A(n2618), .B(n2617), .CI(n2616), .CO(n2513), .S(n2619) );
  MUX2_X1 U2597 ( .A(n2620), .B(n2619), .S(n6117), .Z(n2640) );
  OAI22_X1 U2598 ( .A1(n6116), .A2(n3241), .B1(n2622), .B2(n5635), .ZN(n2626)
         );
  INV_X1 U2599 ( .A(dot_op_b_i[25]), .ZN(n2623) );
  OR2_X1 U2600 ( .A1(dot_op_a_i[24]), .A2(n2623), .ZN(n2624) );
  NAND2_X1 U2601 ( .A1(n2624), .A2(n3482), .ZN(n2625) );
  MUX2_X1 U2602 ( .A(n2626), .B(n2625), .S(n6117), .Z(n2634) );
  NOR2_X1 U2603 ( .A1(n2635), .A2(n2634), .ZN(n5284) );
  FA_X1 U2604 ( .A(n2629), .B(n2628), .CI(n2627), .CO(n2610), .S(n5237) );
  NOR2_X1 U2605 ( .A1(n6118), .A2(n5635), .ZN(n2631) );
  AND2_X1 U2606 ( .A1(dot_op_a_i[8]), .A2(dot_op_b_i[8]), .ZN(n2630) );
  MUX2_X1 U2607 ( .A(n2631), .B(n2630), .S(n6141), .Z(n5236) );
  AND2_X1 U2608 ( .A1(n6116), .A2(op_b_i[0]), .ZN(n2633) );
  AND2_X1 U2609 ( .A1(dot_op_a_i[24]), .A2(dot_op_b_i[24]), .ZN(n2632) );
  MUX2_X1 U2610 ( .A(n2633), .B(n2632), .S(n6143), .Z(n5235) );
  INV_X1 U2611 ( .A(n5287), .ZN(n2636) );
  NAND2_X1 U2612 ( .A1(n2635), .A2(n2634), .ZN(n5285) );
  OAI21_X1 U2613 ( .B1(n5284), .B2(n2636), .A(n5285), .ZN(n5314) );
  FA_X1 U2614 ( .A(n2639), .B(n2638), .CI(n2637), .CO(n2602), .S(n2644) );
  FA_X1 U2615 ( .A(n2642), .B(n2641), .CI(n2640), .CO(n2643), .S(n2635) );
  OR2_X1 U2616 ( .A1(n2644), .A2(n2643), .ZN(n5313) );
  NAND2_X1 U2617 ( .A1(n2644), .A2(n2643), .ZN(n5312) );
  INV_X1 U2618 ( .A(n5312), .ZN(n2645) );
  AOI21_X1 U2619 ( .B1(n5314), .B2(n5313), .A(n2645), .ZN(n2756) );
  NAND2_X1 U2620 ( .A1(n2647), .A2(n2646), .ZN(n2754) );
  OAI21_X1 U2621 ( .B1(n2753), .B2(n2756), .A(n2754), .ZN(n2648) );
  INV_X1 U2622 ( .A(n2648), .ZN(n2808) );
  NAND2_X1 U2623 ( .A1(n2650), .A2(n2649), .ZN(n2806) );
  OAI21_X1 U2624 ( .B1(n2805), .B2(n2808), .A(n2806), .ZN(n3988) );
  XNOR2_X1 U2625 ( .A(n2651), .B(n3988), .ZN(n2653) );
  NAND2_X1 U2626 ( .A1(n2653), .A2(n5615), .ZN(n2662) );
  NAND2_X1 U2627 ( .A1(n2655), .A2(n2654), .ZN(n2657) );
  XNOR2_X1 U2628 ( .A(n2657), .B(n2656), .ZN(n2660) );
  NAND2_X1 U2629 ( .A1(n2659), .A2(n2658), .ZN(n6101) );
  NAND2_X1 U2630 ( .A1(n2659), .A2(n1087), .ZN(n6106) );
  INV_X1 U2631 ( .A(n6106), .ZN(n5605) );
  AOI22_X1 U2632 ( .A1(n2660), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[5]), 
        .ZN(n2661) );
  OAI211_X1 U2633 ( .C1(n5293), .C2(n6095), .A(n2662), .B(n2661), .ZN(n2663)
         );
  AOI21_X1 U2634 ( .B1(n5540), .B2(n5418), .A(n2663), .ZN(n2664) );
  OAI21_X1 U2635 ( .B1(n5510), .B2(n5400), .A(n2664), .ZN(n2665) );
  AOI21_X1 U2636 ( .B1(n5158), .B2(n5507), .A(n2665), .ZN(n2666) );
  INV_X1 U2637 ( .A(n2667), .ZN(n2668) );
  NAND2_X1 U2638 ( .A1(n2669), .A2(n2668), .ZN(result_o[5]) );
  NOR2_X1 U2639 ( .A1(n2670), .A2(n2686), .ZN(n2688) );
  NAND2_X1 U2640 ( .A1(n2671), .A2(n2688), .ZN(n2691) );
  NOR2_X1 U2641 ( .A1(n2691), .A2(n2672), .ZN(n5220) );
  INV_X1 U2642 ( .A(n2673), .ZN(n2674) );
  NOR2_X1 U2643 ( .A1(n2675), .A2(n2674), .ZN(n2704) );
  MUX2_X1 U2644 ( .A(mulh_carry_q), .B(op_c_i[31]), .S(n2713), .Z(n2676) );
  INV_X1 U2645 ( .A(n2676), .ZN(n2706) );
  HA_X1 U2646 ( .A(op_c_i[31]), .B(op_c_i[30]), .CO(n2705), .S(n2678) );
  FA_X1 U2647 ( .A(n2679), .B(n2678), .CI(n2677), .CO(n2702), .S(n2680) );
  FA_X1 U2648 ( .A(n2682), .B(n2681), .CI(n2680), .CO(n2693), .S(n998) );
  OR2_X1 U2649 ( .A1(n2694), .A2(n2693), .ZN(n5223) );
  NAND2_X1 U2650 ( .A1(n5220), .A2(n5223), .ZN(n2697) );
  NOR2_X1 U2651 ( .A1(n2683), .A2(n2697), .ZN(n2700) );
  OAI21_X1 U2652 ( .B1(n2686), .B2(n2685), .A(n2684), .ZN(n2687) );
  AOI21_X1 U2653 ( .B1(n2689), .B2(n2688), .A(n2687), .ZN(n2690) );
  OAI21_X1 U2654 ( .B1(n2692), .B2(n2691), .A(n2690), .ZN(n5219) );
  NAND2_X1 U2655 ( .A1(n2694), .A2(n2693), .ZN(n5222) );
  INV_X1 U2656 ( .A(n5222), .ZN(n2695) );
  AOI21_X1 U2657 ( .B1(n5219), .B2(n5223), .A(n2695), .ZN(n2696) );
  OAI21_X1 U2658 ( .B1(n979), .B2(n2697), .A(n2696), .ZN(n2699) );
  AOI21_X1 U2659 ( .B1(n1002), .B2(n2700), .A(n2699), .ZN(n2701) );
  INV_X1 U2660 ( .A(n2701), .ZN(n2712) );
  FA_X1 U2661 ( .A(n2704), .B(n2703), .CI(n2702), .CO(n2710), .S(n2694) );
  INV_X1 U2662 ( .A(n2704), .ZN(n2708) );
  HA_X1 U2663 ( .A(n2706), .B(n2705), .CO(n2707), .S(n2703) );
  XOR2_X1 U2664 ( .A(n2708), .B(n2707), .Z(n2709) );
  XOR2_X1 U2665 ( .A(n2710), .B(n2709), .Z(n2711) );
  XOR2_X1 U2666 ( .A(n2712), .B(n2711), .Z(n2714) );
  NOR2_X1 U2667 ( .A1(n2714), .A2(n2713), .ZN(n2715) );
  NOR2_X1 U2668 ( .A1(n2829), .A2(n2715), .ZN(n4880) );
  INV_X1 U2670 ( .A(n2831), .ZN(n5171) );
  OR2_X1 U2671 ( .A1(n2716), .A2(n2830), .ZN(n5261) );
  AOI22_X1 U2672 ( .A1(n4956), .A2(n5304), .B1(n4958), .B2(n5331), .ZN(n2718)
         );
  AOI22_X1 U2673 ( .A1(n4963), .A2(n5008), .B1(n4959), .B2(n5302), .ZN(n2717)
         );
  NAND2_X1 U2674 ( .A1(n2718), .A2(n2717), .ZN(n5157) );
  INV_X1 U2675 ( .A(n5157), .ZN(n2725) );
  AOI22_X1 U2676 ( .A1(n4974), .A2(n5331), .B1(n4975), .B2(n5302), .ZN(n2720)
         );
  AOI22_X1 U2677 ( .A1(n5304), .A2(n4976), .B1(n4957), .B2(n5008), .ZN(n2719)
         );
  NAND2_X1 U2678 ( .A1(n2720), .A2(n2719), .ZN(n5431) );
  AOI22_X1 U2679 ( .A1(n5007), .A2(n5304), .B1(n5011), .B2(n5302), .ZN(n2722)
         );
  NAND2_X1 U2680 ( .A1(n4977), .A2(n5311), .ZN(n2721) );
  OAI211_X1 U2681 ( .C1(n2723), .C2(n5307), .A(n2722), .B(n2721), .ZN(n5164)
         );
  OAI22_X1 U2682 ( .A1(n5431), .A2(n5386), .B1(n5164), .B2(n5344), .ZN(n2724)
         );
  AOI21_X1 U2683 ( .B1(n5264), .B2(n2725), .A(n2724), .ZN(n2726) );
  OAI21_X1 U2684 ( .B1(n5171), .B2(n5261), .A(n2726), .ZN(n4940) );
  INV_X1 U2685 ( .A(n4985), .ZN(n2729) );
  AOI22_X1 U2686 ( .A1(n4991), .A2(n5304), .B1(n5302), .B2(n4986), .ZN(n2728)
         );
  NAND2_X1 U2687 ( .A1(n5010), .A2(n5311), .ZN(n2727) );
  OAI211_X1 U2688 ( .C1(n2729), .C2(n5307), .A(n2728), .B(n2727), .ZN(n5439)
         );
  NAND2_X1 U2689 ( .A1(n4987), .A2(n5311), .ZN(n2732) );
  AOI22_X1 U2690 ( .A1(n5302), .A2(n5001), .B1(n4998), .B2(n5304), .ZN(n2731)
         );
  NAND2_X1 U2691 ( .A1(n4999), .A2(n5331), .ZN(n2730) );
  NAND3_X1 U2692 ( .A1(n2732), .A2(n2731), .A3(n2730), .ZN(n5449) );
  INV_X1 U2693 ( .A(n5449), .ZN(n2764) );
  NAND2_X1 U2694 ( .A1(n5000), .A2(n5311), .ZN(n2735) );
  AOI22_X1 U2695 ( .A1(n5301), .A2(n5304), .B1(n5302), .B2(n5305), .ZN(n2734)
         );
  NAND2_X1 U2696 ( .A1(n5310), .A2(n5331), .ZN(n2733) );
  NAND3_X1 U2697 ( .A1(n2735), .A2(n2734), .A3(n2733), .ZN(n5045) );
  INV_X1 U2698 ( .A(n2736), .ZN(n2738) );
  NAND2_X1 U2699 ( .A1(n2738), .A2(n2737), .ZN(n2740) );
  XOR2_X1 U2700 ( .A(n2740), .B(n2739), .Z(n5277) );
  INV_X1 U2701 ( .A(n5277), .ZN(n5332) );
  NAND2_X1 U2702 ( .A1(n2742), .A2(n2741), .ZN(n2744) );
  XNOR2_X1 U2703 ( .A(n2744), .B(n2743), .ZN(n5328) );
  INV_X1 U2704 ( .A(n6095), .ZN(n5898) );
  OAI21_X1 U2705 ( .B1(n5328), .B2(n5325), .A(n5898), .ZN(n2746) );
  NOR2_X1 U2706 ( .A1(n5335), .A2(n5307), .ZN(n2745) );
  AOI211_X1 U2707 ( .C1(n5304), .C2(n5332), .A(n2746), .B(n2745), .ZN(n2747)
         );
  OAI21_X1 U2708 ( .B1(n5303), .B2(n5334), .A(n2747), .ZN(n2761) );
  NAND2_X1 U2709 ( .A1(n2749), .A2(n2748), .ZN(n2751) );
  XNOR2_X1 U2710 ( .A(n2751), .B(n2750), .ZN(n2752) );
  AOI22_X1 U2711 ( .A1(n2752), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[3]), 
        .ZN(n2760) );
  INV_X1 U2712 ( .A(n2753), .ZN(n2755) );
  NAND2_X1 U2713 ( .A1(n2755), .A2(n2754), .ZN(n2757) );
  XOR2_X1 U2714 ( .A(n2757), .B(n2756), .Z(n2758) );
  NAND2_X1 U2715 ( .A1(n2758), .A2(n5615), .ZN(n2759) );
  NAND3_X1 U2716 ( .A1(n2761), .A2(n2760), .A3(n2759), .ZN(n2762) );
  AOI21_X1 U2717 ( .B1(n5045), .B2(n5540), .A(n2762), .ZN(n2763) );
  OAI21_X1 U2718 ( .B1(n2764), .B2(n5400), .A(n2763), .ZN(n2765) );
  INV_X1 U2719 ( .A(n5521), .ZN(n5376) );
  INV_X1 U2720 ( .A(n2766), .ZN(n4909) );
  INV_X1 U2721 ( .A(n4908), .ZN(n2767) );
  AOI21_X1 U2722 ( .B1(n4911), .B2(n4909), .A(n2767), .ZN(n2772) );
  INV_X1 U2723 ( .A(n2768), .ZN(n2770) );
  NAND2_X1 U2724 ( .A1(n2770), .A2(n2769), .ZN(n2771) );
  XOR2_X1 U2725 ( .A(n2772), .B(n2771), .Z(n4907) );
  INV_X1 U2726 ( .A(n4907), .ZN(n5188) );
  AOI21_X1 U2727 ( .B1(n4911), .B2(n2774), .A(n2773), .ZN(n2779) );
  INV_X1 U2728 ( .A(n2775), .ZN(n2777) );
  NAND2_X1 U2729 ( .A1(n2777), .A2(n2776), .ZN(n2778) );
  XOR2_X1 U2730 ( .A(n2779), .B(n2778), .Z(n4934) );
  INV_X1 U2731 ( .A(n4934), .ZN(n4922) );
  INV_X1 U2732 ( .A(n5519), .ZN(n5465) );
  OAI22_X1 U2733 ( .A1(n5376), .A2(n5188), .B1(n4922), .B2(n5465), .ZN(n2781)
         );
  AOI211_X1 U2734 ( .C1(n5183), .C2(n5463), .A(n2781), .B(n2780), .ZN(n4936)
         );
  OR2_X1 U2735 ( .A1(n4936), .A2(n5894), .ZN(n2782) );
  OAI211_X1 U2736 ( .C1(n4940), .C2(n5553), .A(n2783), .B(n2782), .ZN(
        result_o[3]) );
  AOI22_X1 U2737 ( .A1(n5331), .A2(n4963), .B1(n4962), .B2(n5008), .ZN(n2785)
         );
  AOI22_X1 U2738 ( .A1(n5302), .A2(n4956), .B1(n4958), .B2(n5304), .ZN(n2784)
         );
  AND2_X1 U2739 ( .A1(n2785), .A2(n2784), .ZN(n5700) );
  INV_X1 U2740 ( .A(n5700), .ZN(n2791) );
  AOI22_X1 U2741 ( .A1(n4974), .A2(n5304), .B1(n4959), .B2(n5008), .ZN(n2787)
         );
  AOI22_X1 U2742 ( .A1(n5302), .A2(n4976), .B1(n4957), .B2(n5331), .ZN(n2786)
         );
  NAND2_X1 U2743 ( .A1(n2787), .A2(n2786), .ZN(n5383) );
  INV_X1 U2744 ( .A(n5383), .ZN(n5482) );
  AOI22_X1 U2745 ( .A1(n5331), .A2(n4977), .B1(n4975), .B2(n5008), .ZN(n2789)
         );
  AOI22_X1 U2746 ( .A1(n5009), .A2(n5304), .B1(n5302), .B2(n5007), .ZN(n2788)
         );
  AND2_X1 U2747 ( .A1(n2789), .A2(n2788), .ZN(n5481) );
  AOI22_X1 U2748 ( .A1(n5482), .A2(n5257), .B1(n5384), .B2(n5481), .ZN(n2790)
         );
  OAI211_X1 U2749 ( .C1(n2792), .C2(n2791), .A(n79), .B(n2790), .ZN(n4893) );
  INV_X1 U2750 ( .A(n5573), .ZN(n2794) );
  INV_X1 U2751 ( .A(n5463), .ZN(n5488) );
  AOI22_X1 U2752 ( .A1(n5183), .A2(n5519), .B1(n4934), .B2(n5521), .ZN(n2793)
         );
  OAI21_X1 U2753 ( .B1(n2794), .B2(n5488), .A(n2793), .ZN(n2795) );
  AOI22_X1 U2754 ( .A1(n5311), .A2(n5011), .B1(n5010), .B2(n5331), .ZN(n2798)
         );
  AOI22_X1 U2755 ( .A1(n4985), .A2(n5304), .B1(n5302), .B2(n4991), .ZN(n2797)
         );
  AND2_X1 U2756 ( .A1(n2798), .A2(n2797), .ZN(n5551) );
  INV_X1 U2757 ( .A(n5551), .ZN(n2825) );
  NAND2_X1 U2758 ( .A1(n5001), .A2(n5311), .ZN(n2802) );
  AOI22_X1 U2759 ( .A1(n5310), .A2(n5304), .B1(n5301), .B2(n5302), .ZN(n2800)
         );
  NAND2_X1 U2760 ( .A1(n5000), .A2(n5331), .ZN(n2799) );
  AND2_X1 U2761 ( .A1(n2800), .A2(n2799), .ZN(n2801) );
  AND2_X1 U2762 ( .A1(n2802), .A2(n2801), .ZN(n5399) );
  INV_X1 U2763 ( .A(n5540), .ZN(n5477) );
  AOI22_X1 U2764 ( .A1(n5331), .A2(n4987), .B1(n4986), .B2(n5008), .ZN(n2804)
         );
  AOI22_X1 U2765 ( .A1(n4999), .A2(n5304), .B1(n5302), .B2(n4998), .ZN(n2803)
         );
  NAND2_X1 U2766 ( .A1(n2804), .A2(n2803), .ZN(n5474) );
  NAND2_X1 U2767 ( .A1(n5474), .A2(n5529), .ZN(n2823) );
  INV_X1 U2768 ( .A(n2805), .ZN(n2807) );
  NAND2_X1 U2769 ( .A1(n2807), .A2(n2806), .ZN(n2809) );
  XOR2_X1 U2770 ( .A(n2809), .B(n2808), .Z(n2821) );
  INV_X1 U2771 ( .A(n5303), .ZN(n2811) );
  AOI22_X1 U2772 ( .A1(n5335), .A2(n5304), .B1(n5277), .B2(n5302), .ZN(n2810)
         );
  OAI21_X1 U2773 ( .B1(n2811), .B2(n5307), .A(n2810), .ZN(n2812) );
  AOI21_X1 U2774 ( .B1(n5008), .B2(n5305), .A(n2812), .ZN(n5258) );
  INV_X1 U2775 ( .A(n2813), .ZN(n2815) );
  NAND2_X1 U2776 ( .A1(n2815), .A2(n2814), .ZN(n2817) );
  XOR2_X1 U2777 ( .A(n2817), .B(n2816), .Z(n2818) );
  AOI22_X1 U2778 ( .A1(n2818), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[4]), 
        .ZN(n2819) );
  OAI21_X1 U2779 ( .B1(n5258), .B2(n6095), .A(n2819), .ZN(n2820) );
  AOI21_X1 U2780 ( .B1(n2821), .B2(n5615), .A(n2820), .ZN(n2822) );
  OAI211_X1 U2781 ( .C1(n5399), .C2(n5477), .A(n2823), .B(n2822), .ZN(n2824)
         );
  OAI21_X1 U2782 ( .B1(n5215), .B2(mulh_CS[1]), .A(n5210), .ZN(n2828) );
  INV_X1 U2783 ( .A(n2828), .ZN(n465) );
  NOR2_X1 U2784 ( .A1(n2829), .A2(n2830), .ZN(n5382) );
  NOR2_X1 U2785 ( .A1(n2831), .A2(n5386), .ZN(n2832) );
  AOI211_X1 U2786 ( .C1(n5384), .C2(n5157), .A(n5382), .B(n2832), .ZN(n5461)
         );
  INV_X1 U2787 ( .A(n5622), .ZN(n5703) );
  INV_X1 U2788 ( .A(n3312), .ZN(n2835) );
  INV_X1 U2789 ( .A(dot_op_b_i[15]), .ZN(n2833) );
  INV_X1 U2790 ( .A(dot_signed_i[0]), .ZN(n2928) );
  NOR2_X1 U2791 ( .A1(n2833), .A2(n2928), .ZN(n2834) );
  XNOR2_X1 U2792 ( .A(n2834), .B(dot_op_b_i[15]), .ZN(n3500) );
  NOR2_X1 U2793 ( .A1(n2835), .A2(n3500), .ZN(n2845) );
  INV_X1 U2794 ( .A(n2845), .ZN(n2861) );
  AND2_X1 U2795 ( .A1(dot_op_a_i[7]), .A2(dot_signed_i[1]), .ZN(n3314) );
  INV_X1 U2796 ( .A(n3314), .ZN(n2838) );
  INV_X1 U2797 ( .A(dot_op_b_i[7]), .ZN(n2836) );
  NOR2_X1 U2798 ( .A1(n2836), .A2(n2928), .ZN(n2837) );
  XNOR2_X1 U2799 ( .A(n2837), .B(dot_op_b_i[7]), .ZN(n3316) );
  NOR2_X1 U2800 ( .A1(n2838), .A2(n3316), .ZN(n2860) );
  XOR2_X1 U2801 ( .A(dot_op_b_i[7]), .B(dot_op_b_i[6]), .Z(n2839) );
  XNOR2_X1 U2802 ( .A(dot_op_b_i[6]), .B(dot_op_b_i[5]), .ZN(n3532) );
  NAND2_X1 U2803 ( .A1(n2839), .A2(n3532), .ZN(n3489) );
  XNOR2_X1 U2804 ( .A(n3314), .B(dot_op_b_i[7]), .ZN(n2850) );
  AOI21_X1 U2805 ( .B1(n3489), .B2(n63), .A(n2850), .ZN(n3022) );
  INV_X1 U2806 ( .A(n3022), .ZN(n2846) );
  NOR2_X1 U2807 ( .A1(n6119), .A2(n2874), .ZN(n2841) );
  MUX2_X1 U2808 ( .A(n2842), .B(n2841), .S(n29), .Z(n3038) );
  INV_X1 U2809 ( .A(op_c_i[17]), .ZN(n2844) );
  OAI22_X1 U2810 ( .A1(n6146), .A2(n4923), .B1(n2525), .B2(n2844), .ZN(n3037)
         );
  FA_X1 U2811 ( .A(n2860), .B(n2846), .CI(n2845), .CO(n2859), .S(n3032) );
  INV_X1 U2812 ( .A(dot_op_a_i[7]), .ZN(n2847) );
  NOR2_X1 U2813 ( .A1(n2847), .A2(n3316), .ZN(n3023) );
  INV_X1 U2814 ( .A(dot_op_a_i[15]), .ZN(n2848) );
  NOR2_X1 U2815 ( .A1(n2848), .A2(n3500), .ZN(n3021) );
  XNOR2_X1 U2816 ( .A(n3312), .B(dot_op_b_i[15]), .ZN(n2851) );
  XOR2_X1 U2817 ( .A(dot_op_b_i[15]), .B(dot_op_b_i[14]), .Z(n2849) );
  XNOR2_X1 U2818 ( .A(dot_op_a_i[15]), .B(dot_op_b_i[15]), .ZN(n2856) );
  OAI22_X1 U2819 ( .A1(n2851), .A2(n3534), .B1(n3510), .B2(n2856), .ZN(n3014)
         );
  XNOR2_X1 U2820 ( .A(dot_op_a_i[7]), .B(dot_op_b_i[7]), .ZN(n2855) );
  OAI22_X1 U2821 ( .A1(n2850), .A2(n63), .B1(n3489), .B2(n2855), .ZN(n3013) );
  XNOR2_X1 U2822 ( .A(n3314), .B(dot_op_b_i[5]), .ZN(n3091) );
  AOI21_X1 U2823 ( .B1(n3536), .B2(n3539), .A(n3091), .ZN(n3102) );
  INV_X1 U2824 ( .A(n3102), .ZN(n3012) );
  AOI21_X1 U2825 ( .B1(n3510), .B2(n3534), .A(n2851), .ZN(n2852) );
  INV_X1 U2826 ( .A(n2852), .ZN(n3025) );
  INV_X1 U2827 ( .A(dot_op_a_i[14]), .ZN(n2853) );
  NOR2_X1 U2828 ( .A1(n2853), .A2(n3500), .ZN(n3020) );
  INV_X1 U2829 ( .A(dot_op_a_i[6]), .ZN(n2854) );
  NOR2_X1 U2830 ( .A1(n2854), .A2(n3316), .ZN(n3019) );
  XNOR2_X1 U2831 ( .A(dot_op_b_i[7]), .B(dot_op_a_i[6]), .ZN(n3088) );
  OAI22_X1 U2832 ( .A1(n3489), .A2(n3088), .B1(n2855), .B2(n63), .ZN(n3103) );
  XNOR2_X1 U2833 ( .A(dot_op_b_i[15]), .B(dot_op_a_i[14]), .ZN(n3086) );
  OAI22_X1 U2834 ( .A1(n3510), .A2(n3086), .B1(n2856), .B2(n3534), .ZN(n3101)
         );
  AND2_X1 U2835 ( .A1(n2857), .A2(n6144), .ZN(n3036) );
  INV_X1 U2836 ( .A(n2860), .ZN(n2858) );
  AND2_X1 U2837 ( .A1(n2858), .A2(n6144), .ZN(n2993) );
  OAI22_X1 U2838 ( .A1(n6146), .A2(n5187), .B1(n2525), .B2(n251), .ZN(n2992)
         );
  FA_X1 U2839 ( .A(n2861), .B(n2860), .CI(n2859), .CO(n2864), .S(n2842) );
  INV_X1 U2840 ( .A(op_b_i[18]), .ZN(n2862) );
  NOR2_X1 U2841 ( .A1(n6118), .A2(n2862), .ZN(n2863) );
  MUX2_X1 U2842 ( .A(n2864), .B(n2863), .S(n29), .Z(n2991) );
  XNOR2_X1 U2843 ( .A(n6118), .B(op_a_i[13]), .ZN(n6031) );
  XNOR2_X1 U2844 ( .A(n66), .B(n25), .ZN(n2961) );
  XNOR2_X1 U2845 ( .A(n6121), .B(n25), .ZN(n2908) );
  OAI22_X1 U2846 ( .A1(n2961), .A2(n5809), .B1(n2908), .B2(n2867), .ZN(n2943)
         );
  XNOR2_X1 U2847 ( .A(n22), .B(op_b_i[13]), .ZN(n2952) );
  XNOR2_X1 U2848 ( .A(op_b_i[12]), .B(op_b_i[11]), .ZN(n5936) );
  XNOR2_X1 U2849 ( .A(n55), .B(op_b_i[13]), .ZN(n2904) );
  XOR2_X1 U2850 ( .A(op_b_i[12]), .B(op_b_i[13]), .Z(n2868) );
  OAI22_X1 U2851 ( .A1(n2952), .A2(n72), .B1(n2904), .B2(n5934), .ZN(n2942) );
  XNOR2_X1 U2852 ( .A(n6116), .B(op_b_i[17]), .ZN(n2870) );
  XOR2_X1 U2853 ( .A(op_b_i[16]), .B(op_b_i[17]), .Z(n2869) );
  NAND2_X1 U2854 ( .A1(n2869), .A2(n5917), .ZN(n5915) );
  XNOR2_X1 U2855 ( .A(n6002), .B(op_b_i[17]), .ZN(n2950) );
  OAI22_X1 U2856 ( .A1(n2870), .A2(n5915), .B1(n2950), .B2(n5917), .ZN(n2941)
         );
  INV_X1 U2857 ( .A(op_b_i[9]), .ZN(n3386) );
  XNOR2_X1 U2858 ( .A(n21), .B(n27), .ZN(n2951) );
  XNOR2_X1 U2859 ( .A(op_b_i[8]), .B(op_b_i[7]), .ZN(n2871) );
  INV_X1 U2860 ( .A(n2871), .ZN(n3388) );
  INV_X1 U2861 ( .A(n3388), .ZN(n4546) );
  XNOR2_X1 U2862 ( .A(n20), .B(n27), .ZN(n2900) );
  XOR2_X1 U2863 ( .A(op_b_i[8]), .B(n27), .Z(n2872) );
  OAI22_X1 U2864 ( .A1(n2951), .A2(n4546), .B1(n2900), .B2(n5822), .ZN(n2949)
         );
  XNOR2_X1 U2865 ( .A(n5976), .B(n4123), .ZN(n2944) );
  XNOR2_X1 U2866 ( .A(n5848), .B(n4123), .ZN(n2902) );
  XOR2_X1 U2867 ( .A(op_b_i[14]), .B(n4123), .Z(n2873) );
  NAND2_X1 U2868 ( .A1(n2873), .A2(n5927), .ZN(n5925) );
  OAI22_X1 U2869 ( .A1(n2944), .A2(n5927), .B1(n2902), .B2(n5925), .ZN(n2948)
         );
  INV_X1 U2870 ( .A(op_b_i[17]), .ZN(n2874) );
  OR2_X1 U2871 ( .A1(n6116), .A2(n2874), .ZN(n2875) );
  OAI22_X1 U2872 ( .A1(n2875), .A2(n5917), .B1(n5915), .B2(n2874), .ZN(n2947)
         );
  XNOR2_X1 U2873 ( .A(n51), .B(n25), .ZN(n2909) );
  XNOR2_X1 U2874 ( .A(n52), .B(n25), .ZN(n2882) );
  OAI22_X1 U2875 ( .A1(n2909), .A2(n5809), .B1(n2882), .B2(n2867), .ZN(n3051)
         );
  XNOR2_X1 U2876 ( .A(n21), .B(n5919), .ZN(n2907) );
  INV_X1 U2877 ( .A(n2442), .ZN(n5807) );
  XOR2_X1 U2878 ( .A(op_b_i[6]), .B(n5807), .Z(n3900) );
  XNOR2_X1 U2879 ( .A(n20), .B(n5919), .ZN(n2881) );
  INV_X1 U2880 ( .A(n3889), .ZN(n4383) );
  XOR2_X1 U2881 ( .A(op_b_i[6]), .B(n4383), .Z(n2876) );
  OAI22_X1 U2882 ( .A1(n2907), .A2(n5922), .B1(n2881), .B2(n3128), .ZN(n3050)
         );
  XNOR2_X1 U2883 ( .A(n6116), .B(n4123), .ZN(n2877) );
  XNOR2_X1 U2884 ( .A(n6002), .B(n4123), .ZN(n2903) );
  OAI22_X1 U2885 ( .A1(n2877), .A2(n5925), .B1(n2903), .B2(n5927), .ZN(n3049)
         );
  XNOR2_X1 U2886 ( .A(n22), .B(n5941), .ZN(n2899) );
  XOR2_X1 U2887 ( .A(op_b_i[10]), .B(op_b_i[9]), .Z(n3402) );
  XNOR2_X1 U2888 ( .A(n55), .B(op_b_i[11]), .ZN(n2892) );
  XOR2_X1 U2889 ( .A(op_b_i[10]), .B(n5941), .Z(n2878) );
  NAND2_X1 U2890 ( .A1(n2878), .A2(n26), .ZN(n5943) );
  OAI22_X1 U2891 ( .A1(n2899), .A2(n26), .B1(n2892), .B2(n5943), .ZN(n2891) );
  XNOR2_X1 U2892 ( .A(n56), .B(op_b_i[13]), .ZN(n2905) );
  XNOR2_X1 U2893 ( .A(n5848), .B(op_b_i[13]), .ZN(n2883) );
  OAI22_X1 U2894 ( .A1(n2905), .A2(n72), .B1(n2883), .B2(n5934), .ZN(n2890) );
  XNOR2_X1 U2895 ( .A(n2879), .B(op_a_i[7]), .ZN(n5992) );
  XNOR2_X1 U2896 ( .A(n54), .B(n27), .ZN(n2901) );
  XNOR2_X1 U2897 ( .A(n19), .B(n27), .ZN(n2886) );
  OAI22_X1 U2898 ( .A1(n2901), .A2(n2871), .B1(n2886), .B2(n5822), .ZN(n2889)
         );
  XNOR2_X1 U2899 ( .A(n65), .B(n6015), .ZN(n2910) );
  XNOR2_X1 U2900 ( .A(n6121), .B(n6015), .ZN(n2884) );
  OAI22_X1 U2901 ( .A1(n2910), .A2(n10), .B1(n2884), .B2(n2585), .ZN(n2888) );
  OR2_X1 U2902 ( .A1(n6116), .A2(n3107), .ZN(n2880) );
  OAI22_X1 U2903 ( .A1(n2880), .A2(n5927), .B1(n5925), .B2(n3107), .ZN(n2887)
         );
  XNOR2_X1 U2904 ( .A(n54), .B(n5919), .ZN(n3040) );
  OAI22_X1 U2905 ( .A1(n3040), .A2(n3128), .B1(n2881), .B2(n5922), .ZN(n3118)
         );
  XNOR2_X1 U2906 ( .A(n21), .B(n25), .ZN(n3042) );
  OAI22_X1 U2907 ( .A1(n3042), .A2(n2867), .B1(n2882), .B2(n5809), .ZN(n3117)
         );
  XNOR2_X1 U2908 ( .A(n51), .B(n6015), .ZN(n2885) );
  XNOR2_X1 U2909 ( .A(n52), .B(n6015), .ZN(n3127) );
  OAI22_X1 U2910 ( .A1(n2885), .A2(n10), .B1(n3127), .B2(n2585), .ZN(n3125) );
  XNOR2_X1 U2911 ( .A(n66), .B(n5985), .ZN(n2895) );
  XNOR2_X1 U2912 ( .A(n6120), .B(n5985), .ZN(n3123) );
  OAI22_X1 U2913 ( .A1(n2895), .A2(n5635), .B1(n3123), .B2(n3241), .ZN(n3124)
         );
  XNOR2_X1 U2914 ( .A(n6002), .B(op_b_i[13]), .ZN(n3044) );
  OAI22_X1 U2915 ( .A1(n3044), .A2(n5934), .B1(n2883), .B2(n72), .ZN(n3121) );
  OAI22_X1 U2916 ( .A1(n2885), .A2(n2585), .B1(n2884), .B2(n10), .ZN(n3120) );
  XNOR2_X1 U2917 ( .A(n22), .B(n27), .ZN(n3039) );
  OAI22_X1 U2918 ( .A1(n3039), .A2(n5822), .B1(n2886), .B2(n4546), .ZN(n3119)
         );
  FA_X1 U2919 ( .A(n2889), .B(n2888), .CI(n2887), .CO(n2896), .S(n3113) );
  HA_X1 U2920 ( .A(n2891), .B(n2890), .CO(n2897), .S(n3054) );
  XNOR2_X1 U2921 ( .A(n5914), .B(n5985), .ZN(n2911) );
  XNOR2_X1 U2922 ( .A(n5844), .B(n5985), .ZN(n2894) );
  OAI22_X1 U2923 ( .A1(n2911), .A2(n5635), .B1(n2894), .B2(n3241), .ZN(n3053)
         );
  XNOR2_X1 U2924 ( .A(n56), .B(op_b_i[11]), .ZN(n3043) );
  OAI22_X1 U2925 ( .A1(n3043), .A2(n5943), .B1(n2892), .B2(n26), .ZN(n3048) );
  INV_X1 U2926 ( .A(n5927), .ZN(n2893) );
  AND2_X1 U2927 ( .A1(n6116), .A2(n2893), .ZN(n3047) );
  OAI22_X1 U2928 ( .A1(n2895), .A2(n3241), .B1(n2894), .B2(n5635), .ZN(n3046)
         );
  FA_X1 U2929 ( .A(n2898), .B(n2897), .CI(n2896), .CO(n2935), .S(n3058) );
  XNOR2_X1 U2930 ( .A(n19), .B(n5941), .ZN(n2914) );
  OAI22_X1 U2931 ( .A1(n2899), .A2(n5943), .B1(n2914), .B2(n26), .ZN(n2918) );
  OAI22_X1 U2932 ( .A1(n2901), .A2(n5822), .B1(n2900), .B2(n4546), .ZN(n2917)
         );
  OAI22_X1 U2933 ( .A1(n2903), .A2(n5925), .B1(n2902), .B2(n5927), .ZN(n2916)
         );
  OAI22_X1 U2934 ( .A1(n2905), .A2(n5934), .B1(n2904), .B2(n5936), .ZN(n2921)
         );
  INV_X1 U2935 ( .A(n5917), .ZN(n2906) );
  AND2_X1 U2936 ( .A1(n6116), .A2(n2906), .ZN(n2920) );
  XNOR2_X1 U2937 ( .A(n52), .B(n5919), .ZN(n2915) );
  OAI22_X1 U2938 ( .A1(n2907), .A2(n3128), .B1(n2915), .B2(n5922), .ZN(n2919)
         );
  OAI22_X1 U2939 ( .A1(n2909), .A2(n2867), .B1(n2908), .B2(n5809), .ZN(n2924)
         );
  XNOR2_X1 U2940 ( .A(n5844), .B(n6015), .ZN(n2912) );
  OAI22_X1 U2941 ( .A1(n2910), .A2(n2585), .B1(n2912), .B2(n10), .ZN(n2923) );
  XNOR2_X1 U2942 ( .A(n2866), .B(op_a_i[16]), .ZN(n5819) );
  XNOR2_X1 U2943 ( .A(n5819), .B(n5985), .ZN(n2913) );
  OAI22_X1 U2944 ( .A1(n2911), .A2(n3241), .B1(n2913), .B2(n5635), .ZN(n2922)
         );
  XNOR2_X1 U2945 ( .A(n5914), .B(n6015), .ZN(n2940) );
  OAI22_X1 U2946 ( .A1(n2940), .A2(n10), .B1(n2912), .B2(n2585), .ZN(n2967) );
  XNOR2_X1 U2947 ( .A(n2866), .B(op_a_i[17]), .ZN(n5924) );
  XNOR2_X1 U2948 ( .A(n5924), .B(n5985), .ZN(n2964) );
  OAI22_X1 U2949 ( .A1(n2964), .A2(n5635), .B1(n2913), .B2(n3241), .ZN(n2966)
         );
  XNOR2_X1 U2950 ( .A(n54), .B(op_b_i[11]), .ZN(n2962) );
  OAI22_X1 U2951 ( .A1(n2962), .A2(n26), .B1(n2914), .B2(n5943), .ZN(n2939) );
  XNOR2_X1 U2952 ( .A(n51), .B(n5919), .ZN(n2946) );
  OAI22_X1 U2953 ( .A1(n2946), .A2(n5922), .B1(n2915), .B2(n3128), .ZN(n2938)
         );
  FA_X1 U2954 ( .A(n2918), .B(n2917), .CI(n2916), .CO(n2970), .S(n3057) );
  FA_X1 U2955 ( .A(n2921), .B(n2920), .CI(n2919), .CO(n2969), .S(n3056) );
  FA_X1 U2956 ( .A(n2924), .B(n2923), .CI(n2922), .CO(n2968), .S(n3055) );
  INV_X1 U2957 ( .A(n3407), .ZN(n2927) );
  NOR2_X1 U2958 ( .A1(n2925), .A2(n2928), .ZN(n2926) );
  XNOR2_X1 U2959 ( .A(n2926), .B(dot_op_b_i[31]), .ZN(n3430) );
  NOR2_X1 U2960 ( .A1(n2927), .A2(n3430), .ZN(n3133) );
  INV_X1 U2961 ( .A(n3133), .ZN(n3062) );
  AND2_X1 U2962 ( .A1(dot_op_a_i[23]), .A2(dot_signed_i[1]), .ZN(n3405) );
  INV_X1 U2963 ( .A(n3405), .ZN(n2931) );
  NOR2_X1 U2964 ( .A1(n2929), .A2(n2928), .ZN(n2930) );
  XNOR2_X1 U2965 ( .A(n2930), .B(dot_op_b_i[23]), .ZN(n3448) );
  NOR2_X1 U2966 ( .A1(n2931), .A2(n3448), .ZN(n3135) );
  XOR2_X1 U2967 ( .A(dot_op_b_i[22]), .B(dot_op_b_i[23]), .Z(n2932) );
  XNOR2_X1 U2968 ( .A(dot_op_b_i[22]), .B(dot_op_b_i[21]), .ZN(n3467) );
  NAND2_X1 U2969 ( .A1(n2932), .A2(n3467), .ZN(n3469) );
  XNOR2_X1 U2970 ( .A(n3405), .B(dot_op_b_i[23]), .ZN(n3140) );
  AOI21_X1 U2971 ( .B1(n3469), .B2(n61), .A(n3140), .ZN(n3143) );
  INV_X1 U2972 ( .A(n3143), .ZN(n3134) );
  MUX2_X1 U2973 ( .A(n2934), .B(n2933), .S(n6144), .Z(n3065) );
  FA_X1 U2974 ( .A(n2937), .B(n2936), .CI(n2935), .CO(n3005), .S(n3149) );
  HA_X1 U2975 ( .A(n2939), .B(n2938), .CO(n2955), .S(n2965) );
  XNOR2_X1 U2976 ( .A(n5819), .B(n6015), .ZN(n2956) );
  OAI22_X1 U2977 ( .A1(n2940), .A2(n2585), .B1(n2956), .B2(n10), .ZN(n2954) );
  FA_X1 U2978 ( .A(n2943), .B(n2942), .CI(n2941), .CO(n2953), .S(n2937) );
  XNOR2_X1 U2979 ( .A(n55), .B(n4123), .ZN(n2979) );
  OAI22_X1 U2980 ( .A1(n2944), .A2(n5925), .B1(n2979), .B2(n5927), .ZN(n2973)
         );
  INV_X1 U2981 ( .A(n6034), .ZN(n2945) );
  AND2_X1 U2982 ( .A1(n6116), .A2(n2945), .ZN(n2972) );
  XNOR2_X1 U2983 ( .A(n6121), .B(n5919), .ZN(n2975) );
  OAI22_X1 U2984 ( .A1(n2946), .A2(n3128), .B1(n2975), .B2(n5922), .ZN(n2971)
         );
  FA_X1 U2985 ( .A(n2949), .B(n2948), .CI(n2947), .CO(n2958), .S(n2936) );
  XNOR2_X1 U2986 ( .A(n5848), .B(op_b_i[17]), .ZN(n2980) );
  OAI22_X1 U2987 ( .A1(n2950), .A2(n5915), .B1(n2980), .B2(n5917), .ZN(n2978)
         );
  XNOR2_X1 U2988 ( .A(n52), .B(n27), .ZN(n2987) );
  OAI22_X1 U2989 ( .A1(n2951), .A2(n5822), .B1(n2987), .B2(n4546), .ZN(n2977)
         );
  XNOR2_X1 U2990 ( .A(n19), .B(op_b_i[13]), .ZN(n2974) );
  OAI22_X1 U2991 ( .A1(n2952), .A2(n5934), .B1(n2974), .B2(n72), .ZN(n2976) );
  FA_X1 U2992 ( .A(n2955), .B(n2954), .CI(n2953), .CO(n4107), .S(n3004) );
  XNOR2_X1 U2993 ( .A(n5914), .B(n25), .ZN(n4136) );
  XNOR2_X1 U2994 ( .A(n5844), .B(n25), .ZN(n2960) );
  OAI22_X1 U2995 ( .A1(n4136), .A2(n5809), .B1(n2960), .B2(n2867), .ZN(n4104)
         );
  XNOR2_X1 U2996 ( .A(n6118), .B(op_a_i[19]), .ZN(n5933) );
  XNOR2_X1 U2997 ( .A(n5933), .B(n5985), .ZN(n4095) );
  XNOR2_X1 U2998 ( .A(n6118), .B(op_a_i[18]), .ZN(n5824) );
  XNOR2_X1 U2999 ( .A(n5824), .B(n5985), .ZN(n2963) );
  OAI22_X1 U3000 ( .A1(n4095), .A2(n5635), .B1(n2963), .B2(n3241), .ZN(n4103)
         );
  XNOR2_X1 U3001 ( .A(n5924), .B(n6015), .ZN(n4139) );
  OAI22_X1 U3002 ( .A1(n4139), .A2(n10), .B1(n2956), .B2(n2585), .ZN(n4102) );
  FA_X1 U3003 ( .A(n2959), .B(n2958), .CI(n2957), .CO(n4105), .S(n3003) );
  OAI22_X1 U3004 ( .A1(n2961), .A2(n2867), .B1(n2960), .B2(n5809), .ZN(n2986)
         );
  XNOR2_X1 U3005 ( .A(n20), .B(n5941), .ZN(n2988) );
  OAI22_X1 U3006 ( .A1(n2962), .A2(n5943), .B1(n2988), .B2(n26), .ZN(n2985) );
  OAI22_X1 U3007 ( .A1(n2964), .A2(n3241), .B1(n2963), .B2(n5635), .ZN(n2984)
         );
  FA_X1 U3008 ( .A(n2967), .B(n2966), .CI(n2965), .CO(n3001), .S(n2998) );
  FA_X1 U3009 ( .A(n2970), .B(n2969), .CI(n2968), .CO(n3000), .S(n2997) );
  FA_X1 U3010 ( .A(n2973), .B(n2972), .CI(n2971), .CO(n4144), .S(n2959) );
  XNOR2_X1 U3011 ( .A(n54), .B(op_b_i[13]), .ZN(n4093) );
  OAI22_X1 U3012 ( .A1(n4093), .A2(n5936), .B1(n2974), .B2(n5934), .ZN(n4141)
         );
  XNOR2_X1 U3013 ( .A(n6031), .B(n5919), .ZN(n4094) );
  OAI22_X1 U3014 ( .A1(n4094), .A2(n5922), .B1(n2975), .B2(n3128), .ZN(n4140)
         );
  FA_X1 U3015 ( .A(n2978), .B(n2977), .CI(n2976), .CO(n4142), .S(n2957) );
  XNOR2_X1 U3016 ( .A(n22), .B(n4123), .ZN(n4090) );
  OAI22_X1 U3017 ( .A1(n4090), .A2(n5927), .B1(n2979), .B2(n5925), .ZN(n4098)
         );
  XNOR2_X1 U3018 ( .A(n56), .B(op_b_i[17]), .ZN(n4088) );
  OAI22_X1 U3019 ( .A1(n4088), .A2(n5917), .B1(n2980), .B2(n5915), .ZN(n4097)
         );
  INV_X1 U3020 ( .A(op_b_i[19]), .ZN(n2982) );
  OR2_X1 U3021 ( .A1(n6116), .A2(n2982), .ZN(n2983) );
  XOR2_X1 U3022 ( .A(op_b_i[18]), .B(op_b_i[19]), .Z(n2981) );
  OAI22_X1 U3023 ( .A1(n2983), .A2(n6034), .B1(n6032), .B2(n2982), .ZN(n4096)
         );
  FA_X1 U3024 ( .A(n2986), .B(n2985), .CI(n2984), .CO(n4149), .S(n3002) );
  XNOR2_X1 U3025 ( .A(n51), .B(n27), .ZN(n4092) );
  OAI22_X1 U3026 ( .A1(n4092), .A2(n2871), .B1(n2987), .B2(n5822), .ZN(n4101)
         );
  XNOR2_X1 U3027 ( .A(n21), .B(n5941), .ZN(n4089) );
  OAI22_X1 U3028 ( .A1(n4089), .A2(n26), .B1(n2988), .B2(n5943), .ZN(n4100) );
  XNOR2_X1 U3029 ( .A(n6116), .B(op_b_i[19]), .ZN(n2989) );
  XNOR2_X1 U3030 ( .A(n6002), .B(op_b_i[19]), .ZN(n4091) );
  OAI22_X1 U3031 ( .A1(n2989), .A2(n6032), .B1(n4091), .B2(n6034), .ZN(n4099)
         );
  AND2_X1 U3032 ( .A1(n2990), .A2(n29), .ZN(n4296) );
  FA_X1 U3033 ( .A(n2993), .B(n2992), .CI(n2991), .CO(n4284), .S(n3066) );
  NOR2_X1 U3034 ( .A1(n6118), .A2(n2982), .ZN(n2994) );
  OR2_X1 U3035 ( .A1(n2994), .A2(n6145), .ZN(n4267) );
  INV_X1 U3036 ( .A(op_c_i[19]), .ZN(n2995) );
  OAI22_X1 U3037 ( .A1(n6146), .A2(n2996), .B1(n2525), .B2(n2995), .ZN(n4266)
         );
  FA_X1 U3038 ( .A(n2999), .B(n2998), .CI(n2997), .CO(n3009), .S(n3147) );
  FA_X1 U3039 ( .A(n3002), .B(n3001), .CI(n3000), .CO(n4246), .S(n3008) );
  FA_X1 U3040 ( .A(n3005), .B(n3004), .CI(n3003), .CO(n4270), .S(n3007) );
  OR2_X1 U3041 ( .A1(n3006), .A2(n6145), .ZN(n4282) );
  FA_X1 U3042 ( .A(n3009), .B(n3008), .CI(n3007), .CO(n3006), .S(n3011) );
  INV_X1 U3043 ( .A(n3135), .ZN(n3010) );
  MUX2_X1 U3044 ( .A(n3011), .B(n3010), .S(n6117), .Z(n3070) );
  FA_X1 U3045 ( .A(n3014), .B(n3013), .CI(n3012), .CO(n3026), .S(n3106) );
  INV_X1 U3046 ( .A(dot_op_a_i[5]), .ZN(n3015) );
  NOR2_X1 U3047 ( .A1(n3015), .A2(n3316), .ZN(n3081) );
  INV_X1 U3048 ( .A(dot_op_a_i[13]), .ZN(n3016) );
  NOR2_X1 U3049 ( .A1(n3016), .A2(n3500), .ZN(n3080) );
  XNOR2_X1 U3050 ( .A(n3312), .B(dot_op_b_i[13]), .ZN(n3093) );
  AOI21_X1 U3051 ( .B1(n3511), .B2(n3514), .A(n3093), .ZN(n3017) );
  INV_X1 U3052 ( .A(n3017), .ZN(n3079) );
  FA_X1 U3053 ( .A(n3020), .B(n3019), .CI(n3018), .CO(n3024), .S(n3104) );
  FA_X1 U3054 ( .A(n3023), .B(n3022), .CI(n3021), .CO(n3031), .S(n3072) );
  FA_X1 U3055 ( .A(n3026), .B(n3025), .CI(n3024), .CO(n3030), .S(n3071) );
  AND2_X1 U3056 ( .A1(n3027), .A2(n6145), .ZN(n3112) );
  INV_X1 U3057 ( .A(op_c_i[16]), .ZN(n3028) );
  OAI22_X1 U3058 ( .A1(n6146), .A2(n3029), .B1(n2525), .B2(n3028), .ZN(n3111)
         );
  FA_X1 U3059 ( .A(n3032), .B(n3031), .CI(n3030), .CO(n2857), .S(n3035) );
  INV_X1 U3060 ( .A(op_b_i[16]), .ZN(n3033) );
  NOR2_X1 U3061 ( .A1(n6119), .A2(n3033), .ZN(n3034) );
  MUX2_X1 U3062 ( .A(n3035), .B(n3034), .S(n29), .Z(n3110) );
  FA_X1 U3063 ( .A(n3038), .B(n3037), .CI(n3036), .CO(n3067), .S(n3156) );
  XNOR2_X1 U3064 ( .A(n55), .B(n27), .ZN(n3122) );
  OAI22_X1 U3065 ( .A1(n3039), .A2(n2871), .B1(n3122), .B2(n5822), .ZN(n3239)
         );
  XNOR2_X1 U3066 ( .A(n19), .B(n5919), .ZN(n3129) );
  OAI22_X1 U3067 ( .A1(n3040), .A2(n5922), .B1(n3129), .B2(n3128), .ZN(n3238)
         );
  OR2_X1 U3068 ( .A1(n6116), .A2(n3330), .ZN(n3041) );
  OAI22_X1 U3069 ( .A1(n3041), .A2(n72), .B1(n5934), .B2(n3330), .ZN(n3237) );
  XNOR2_X1 U3070 ( .A(n20), .B(n25), .ZN(n3243) );
  OAI22_X1 U3071 ( .A1(n3042), .A2(n6010), .B1(n3243), .B2(n2867), .ZN(n3236)
         );
  XNOR2_X1 U3072 ( .A(n5848), .B(n5941), .ZN(n3126) );
  OAI22_X1 U3073 ( .A1(n3043), .A2(n26), .B1(n3126), .B2(n5943), .ZN(n3235) );
  XNOR2_X1 U3074 ( .A(n6116), .B(op_b_i[13]), .ZN(n3045) );
  OAI22_X1 U3075 ( .A1(n3045), .A2(n5934), .B1(n3044), .B2(n72), .ZN(n3234) );
  FA_X1 U3076 ( .A(n3048), .B(n3047), .CI(n3046), .CO(n3052), .S(n3231) );
  FA_X1 U3077 ( .A(n3051), .B(n3050), .CI(n3049), .CO(n2898), .S(n3131) );
  FA_X1 U3078 ( .A(n3054), .B(n3053), .CI(n3052), .CO(n3059), .S(n3130) );
  FA_X1 U3079 ( .A(n3057), .B(n3056), .CI(n3055), .CO(n2999), .S(n3162) );
  FA_X1 U3080 ( .A(n3060), .B(n3059), .CI(n3058), .CO(n3148), .S(n3161) );
  FA_X1 U3081 ( .A(n3062), .B(n3135), .CI(n3061), .CO(n2933), .S(n3063) );
  MUX2_X1 U3082 ( .A(n3064), .B(n3063), .S(n6145), .Z(n3155) );
  FA_X1 U3083 ( .A(n3067), .B(n3066), .CI(n3065), .CO(n4297), .S(n3068) );
  NOR2_X1 U3084 ( .A1(n4075), .A2(n4074), .ZN(n4929) );
  FA_X1 U3085 ( .A(n3070), .B(n3069), .CI(n3068), .CO(n4074), .S(n4073) );
  FA_X1 U3086 ( .A(n3073), .B(n3072), .CI(n3071), .CO(n3027), .S(n3074) );
  AND2_X1 U3087 ( .A1(n3074), .A2(n6145), .ZN(n3189) );
  INV_X1 U3088 ( .A(op_c_i[15]), .ZN(n3075) );
  OAI22_X1 U3089 ( .A1(n6112), .A2(n3076), .B1(n2525), .B2(n3075), .ZN(n3188)
         );
  XNOR2_X1 U3090 ( .A(dot_op_b_i[5]), .B(dot_op_a_i[6]), .ZN(n3082) );
  XNOR2_X1 U3091 ( .A(dot_op_a_i[7]), .B(dot_op_b_i[5]), .ZN(n3090) );
  OAI22_X1 U3092 ( .A1(n3539), .A2(n3082), .B1(n3090), .B2(n3536), .ZN(n3201)
         );
  XNOR2_X1 U3093 ( .A(n3314), .B(dot_op_b_i[3]), .ZN(n3204) );
  AOI21_X1 U3094 ( .B1(n3549), .B2(n3551), .A(n3204), .ZN(n3200) );
  XNOR2_X1 U3095 ( .A(dot_op_b_i[7]), .B(dot_op_a_i[4]), .ZN(n3202) );
  XNOR2_X1 U3096 ( .A(dot_op_a_i[5]), .B(dot_op_b_i[7]), .ZN(n3089) );
  OAI22_X1 U3097 ( .A1(n3489), .A2(n3202), .B1(n3089), .B2(n63), .ZN(n3199) );
  INV_X1 U3098 ( .A(dot_op_a_i[12]), .ZN(n3077) );
  NOR2_X1 U3099 ( .A1(n3077), .A2(n3500), .ZN(n3197) );
  XNOR2_X1 U3100 ( .A(dot_op_b_i[13]), .B(dot_op_a_i[14]), .ZN(n3203) );
  XNOR2_X1 U3101 ( .A(dot_op_a_i[15]), .B(dot_op_b_i[13]), .ZN(n3092) );
  OAI22_X1 U3102 ( .A1(n3514), .A2(n3203), .B1(n3092), .B2(n3511), .ZN(n3218)
         );
  XNOR2_X1 U3103 ( .A(dot_op_b_i[15]), .B(dot_op_a_i[12]), .ZN(n3083) );
  XNOR2_X1 U3104 ( .A(dot_op_a_i[13]), .B(dot_op_b_i[15]), .ZN(n3087) );
  OAI22_X1 U3105 ( .A1(n3510), .A2(n3083), .B1(n3087), .B2(n3534), .ZN(n3217)
         );
  INV_X1 U3106 ( .A(dot_op_a_i[3]), .ZN(n3078) );
  NOR2_X1 U3107 ( .A1(n3078), .A2(n3316), .ZN(n3216) );
  FA_X1 U3108 ( .A(n3081), .B(n3080), .CI(n3079), .CO(n3105), .S(n3226) );
  XNOR2_X1 U3109 ( .A(dot_op_a_i[5]), .B(dot_op_b_i[5]), .ZN(n3214) );
  OAI22_X1 U3110 ( .A1(n3539), .A2(n3214), .B1(n3536), .B2(n3082), .ZN(n3212)
         );
  XNOR2_X1 U3111 ( .A(dot_op_a_i[11]), .B(dot_op_b_i[15]), .ZN(n3210) );
  OAI22_X1 U3112 ( .A1(n3510), .A2(n3210), .B1(n3083), .B2(n3534), .ZN(n3211)
         );
  OR2_X1 U3113 ( .A1(n3212), .A2(n3211), .ZN(n3221) );
  INV_X1 U3114 ( .A(dot_op_a_i[11]), .ZN(n3084) );
  NOR2_X1 U3115 ( .A1(n3084), .A2(n3500), .ZN(n3220) );
  XNOR2_X1 U3116 ( .A(n3312), .B(dot_op_b_i[11]), .ZN(n3206) );
  AOI21_X1 U3117 ( .B1(n3493), .B2(n3496), .A(n3206), .ZN(n3085) );
  INV_X1 U3118 ( .A(n3085), .ZN(n3219) );
  OAI22_X1 U3119 ( .A1(n3510), .A2(n3087), .B1(n3086), .B2(n3534), .ZN(n3100)
         );
  OAI22_X1 U3120 ( .A1(n3489), .A2(n3089), .B1(n3088), .B2(n63), .ZN(n3099) );
  OAI22_X1 U3121 ( .A1(n3091), .A2(n3536), .B1(n3539), .B2(n3090), .ZN(n3098)
         );
  INV_X1 U3122 ( .A(n3200), .ZN(n3097) );
  OAI22_X1 U3123 ( .A1(n3093), .A2(n3511), .B1(n3514), .B2(n3092), .ZN(n3096)
         );
  INV_X1 U3124 ( .A(dot_op_a_i[4]), .ZN(n3094) );
  NOR2_X1 U3125 ( .A1(n3094), .A2(n3316), .ZN(n3095) );
  FA_X1 U3126 ( .A(n3097), .B(n3096), .CI(n3095), .CO(n3224), .S(n3324) );
  FA_X1 U3127 ( .A(n3100), .B(n3099), .CI(n3098), .CO(n3223), .S(n3325) );
  FA_X1 U3128 ( .A(n3103), .B(n3102), .CI(n3101), .CO(n3018), .S(n3222) );
  FA_X1 U3129 ( .A(n3106), .B(n3105), .CI(n3104), .CO(n3073), .S(n3190) );
  INV_X1 U3130 ( .A(op_b_i[15]), .ZN(n3107) );
  NOR2_X1 U3131 ( .A1(n6119), .A2(n3107), .ZN(n3108) );
  MUX2_X1 U3132 ( .A(n3109), .B(n3108), .S(n29), .Z(n3187) );
  FA_X1 U3133 ( .A(n3112), .B(n3111), .CI(n3110), .CO(n3157), .S(n3279) );
  FA_X1 U3134 ( .A(n3115), .B(n3114), .CI(n3113), .CO(n3060), .S(n3286) );
  FA_X1 U3135 ( .A(n3118), .B(n3117), .CI(n3116), .CO(n3115), .S(n3250) );
  FA_X1 U3136 ( .A(n3121), .B(n3120), .CI(n3119), .CO(n3114), .S(n3249) );
  XNOR2_X1 U3137 ( .A(n56), .B(n27), .ZN(n3240) );
  OAI22_X1 U3138 ( .A1(n3240), .A2(n5822), .B1(n3122), .B2(n4546), .ZN(n3338)
         );
  AND2_X1 U3139 ( .A1(n6116), .A2(n71), .ZN(n3337) );
  XNOR2_X1 U3140 ( .A(n51), .B(n4337), .ZN(n3242) );
  OAI22_X1 U3141 ( .A1(n3242), .A2(n3241), .B1(n3123), .B2(n5635), .ZN(n3336)
         );
  HA_X1 U3142 ( .A(n3125), .B(n3124), .CO(n3116), .S(n3344) );
  XNOR2_X1 U3143 ( .A(n6002), .B(op_b_i[11]), .ZN(n3246) );
  OAI22_X1 U3144 ( .A1(n3246), .A2(n5943), .B1(n3126), .B2(n26), .ZN(n3335) );
  XNOR2_X1 U3145 ( .A(n21), .B(n6015), .ZN(n3340) );
  OAI22_X1 U3146 ( .A1(n3340), .A2(n2585), .B1(n3127), .B2(n10), .ZN(n3334) );
  XNOR2_X1 U3147 ( .A(n22), .B(n5919), .ZN(n3245) );
  OAI22_X1 U3148 ( .A1(n3245), .A2(n3128), .B1(n3129), .B2(n5922), .ZN(n3333)
         );
  FA_X1 U3149 ( .A(n3132), .B(n3131), .CI(n3130), .CO(n3163), .S(n3284) );
  FA_X1 U3150 ( .A(n3135), .B(n3134), .CI(n3133), .CO(n3061), .S(n3152) );
  XOR2_X1 U3151 ( .A(dot_op_b_i[30]), .B(dot_op_b_i[31]), .Z(n3136) );
  XNOR2_X1 U3152 ( .A(dot_op_b_i[30]), .B(dot_op_b_i[29]), .ZN(n3472) );
  NAND2_X1 U3153 ( .A1(n3136), .A2(n3472), .ZN(n3474) );
  XNOR2_X1 U3154 ( .A(n3407), .B(dot_op_b_i[31]), .ZN(n3139) );
  AOI21_X1 U3155 ( .B1(n3474), .B2(n62), .A(n3139), .ZN(n3137) );
  INV_X1 U3156 ( .A(n3137), .ZN(n3144) );
  INV_X1 U3157 ( .A(dot_op_a_i[23]), .ZN(n3138) );
  NOR2_X1 U3158 ( .A1(n3138), .A2(n3448), .ZN(n3142) );
  XNOR2_X1 U3159 ( .A(dot_op_b_i[31]), .B(dot_op_a_i[31]), .ZN(n3175) );
  OAI22_X1 U3160 ( .A1(n3474), .A2(n3175), .B1(n3139), .B2(n62), .ZN(n3166) );
  XNOR2_X1 U3161 ( .A(dot_op_b_i[23]), .B(dot_op_a_i[23]), .ZN(n3173) );
  OAI22_X1 U3162 ( .A1(n3469), .A2(n3173), .B1(n3140), .B2(n61), .ZN(n3165) );
  XNOR2_X1 U3163 ( .A(n3405), .B(dot_op_b_i[21]), .ZN(n3171) );
  AOI21_X1 U3164 ( .B1(n59), .B2(n3721), .A(n3171), .ZN(n3180) );
  INV_X1 U3165 ( .A(n3180), .ZN(n3164) );
  INV_X1 U3166 ( .A(dot_op_a_i[31]), .ZN(n3141) );
  NOR2_X1 U3167 ( .A1(n3141), .A2(n3430), .ZN(n3183) );
  FA_X1 U3168 ( .A(n3144), .B(n3143), .CI(n3142), .CO(n3151), .S(n3182) );
  MUX2_X1 U3169 ( .A(n3146), .B(n3145), .S(n6143), .Z(n3278) );
  FA_X1 U3170 ( .A(n3149), .B(n3148), .CI(n3147), .CO(n2934), .S(n3154) );
  FA_X1 U3171 ( .A(n3152), .B(n3151), .CI(n3150), .CO(n3153), .S(n3145) );
  MUX2_X1 U3172 ( .A(n3154), .B(n3153), .S(n6141), .Z(n3159) );
  FA_X1 U3173 ( .A(n3157), .B(n3156), .CI(n3155), .CO(n3069), .S(n3158) );
  NOR2_X1 U3174 ( .A1(n4073), .A2(n4072), .ZN(n5177) );
  NOR2_X1 U3175 ( .A1(n4929), .A2(n5177), .ZN(n4077) );
  FA_X1 U3176 ( .A(n3160), .B(n3159), .CI(n3158), .CO(n4072), .S(n4071) );
  FA_X1 U3177 ( .A(n3163), .B(n3162), .CI(n3161), .CO(n3064), .S(n3186) );
  FA_X1 U3178 ( .A(n3166), .B(n3165), .CI(n3164), .CO(n3184), .S(n3275) );
  INV_X1 U3179 ( .A(dot_op_a_i[21]), .ZN(n3167) );
  NOR2_X1 U3180 ( .A1(n3167), .A2(n3448), .ZN(n3259) );
  XNOR2_X1 U3181 ( .A(n3407), .B(dot_op_b_i[29]), .ZN(n3172) );
  AOI21_X1 U3182 ( .B1(n3717), .B2(n3715), .A(n3172), .ZN(n3168) );
  INV_X1 U3183 ( .A(n3168), .ZN(n3258) );
  INV_X1 U3184 ( .A(dot_op_a_i[29]), .ZN(n3169) );
  NOR2_X1 U3185 ( .A1(n3169), .A2(n3430), .ZN(n3257) );
  XNOR2_X1 U3186 ( .A(n3405), .B(dot_op_b_i[19]), .ZN(n3355) );
  AOI21_X1 U3187 ( .B1(n60), .B2(n3465), .A(n3355), .ZN(n3353) );
  INV_X1 U3188 ( .A(n3353), .ZN(n3269) );
  XNOR2_X1 U3189 ( .A(dot_op_b_i[31]), .B(dot_op_a_i[29]), .ZN(n3255) );
  XNOR2_X1 U3190 ( .A(dot_op_b_i[31]), .B(dot_op_a_i[30]), .ZN(n3176) );
  OAI22_X1 U3191 ( .A1(n3474), .A2(n3255), .B1(n62), .B2(n3176), .ZN(n3268) );
  INV_X1 U3192 ( .A(dot_op_a_i[28]), .ZN(n3170) );
  NOR2_X1 U3193 ( .A1(n3170), .A2(n3430), .ZN(n3267) );
  XNOR2_X1 U3194 ( .A(dot_op_b_i[21]), .B(dot_op_a_i[23]), .ZN(n3251) );
  OAI22_X1 U3195 ( .A1(n3721), .A2(n3251), .B1(n3171), .B2(n59), .ZN(n3262) );
  XNOR2_X1 U3196 ( .A(dot_op_b_i[23]), .B(dot_op_a_i[21]), .ZN(n3252) );
  XNOR2_X1 U3197 ( .A(dot_op_b_i[23]), .B(dot_op_a_i[22]), .ZN(n3174) );
  OAI22_X1 U3198 ( .A1(n3469), .A2(n3252), .B1(n61), .B2(n3174), .ZN(n3261) );
  XNOR2_X1 U3199 ( .A(dot_op_b_i[29]), .B(dot_op_a_i[31]), .ZN(n3254) );
  OAI22_X1 U3200 ( .A1(n3717), .A2(n3254), .B1(n3172), .B2(n3715), .ZN(n3260)
         );
  OAI22_X1 U3201 ( .A1(n3469), .A2(n3174), .B1(n61), .B2(n3173), .ZN(n3181) );
  OAI22_X1 U3202 ( .A1(n3474), .A2(n3176), .B1(n62), .B2(n3175), .ZN(n3179) );
  INV_X1 U3203 ( .A(dot_op_a_i[30]), .ZN(n3177) );
  NOR2_X1 U3204 ( .A1(n3177), .A2(n3430), .ZN(n3272) );
  INV_X1 U3205 ( .A(dot_op_a_i[22]), .ZN(n3178) );
  NOR2_X1 U3206 ( .A1(n3178), .A2(n3448), .ZN(n3271) );
  FA_X1 U3207 ( .A(n3181), .B(n3180), .CI(n3179), .CO(n3270), .S(n3375) );
  FA_X1 U3208 ( .A(n3184), .B(n3183), .CI(n3182), .CO(n3150), .S(n3287) );
  MUX2_X1 U3209 ( .A(n3186), .B(n3185), .S(n6117), .Z(n3283) );
  FA_X1 U3210 ( .A(n3189), .B(n3188), .CI(n3187), .CO(n3280), .S(n3385) );
  FA_X1 U3211 ( .A(n3192), .B(n3191), .CI(n3190), .CO(n3109), .S(n3193) );
  AND2_X1 U3212 ( .A1(n3193), .A2(n6145), .ZN(n3294) );
  INV_X1 U3213 ( .A(op_c_i[14]), .ZN(n3194) );
  OAI22_X1 U3214 ( .A1(n6112), .A2(n3195), .B1(n2525), .B2(n3194), .ZN(n3293)
         );
  FA_X1 U3215 ( .A(n3198), .B(n3197), .CI(n3196), .CO(n3227), .S(n3329) );
  FA_X1 U3216 ( .A(n3201), .B(n3200), .CI(n3199), .CO(n3198), .S(n3303) );
  XNOR2_X1 U3217 ( .A(dot_op_a_i[3]), .B(dot_op_b_i[7]), .ZN(n3209) );
  OAI22_X1 U3218 ( .A1(n3489), .A2(n3209), .B1(n3202), .B2(n63), .ZN(n3308) );
  XNOR2_X1 U3219 ( .A(dot_op_a_i[13]), .B(dot_op_b_i[13]), .ZN(n3213) );
  OAI22_X1 U3220 ( .A1(n3514), .A2(n3213), .B1(n3511), .B2(n3203), .ZN(n3307)
         );
  XNOR2_X1 U3221 ( .A(dot_op_a_i[7]), .B(dot_op_b_i[3]), .ZN(n3215) );
  OAI22_X1 U3222 ( .A1(n3204), .A2(n3549), .B1(n3551), .B2(n3215), .ZN(n3306)
         );
  INV_X1 U3223 ( .A(dot_op_a_i[2]), .ZN(n3205) );
  NOR2_X1 U3224 ( .A1(n3205), .A2(n3316), .ZN(n3320) );
  XNOR2_X1 U3225 ( .A(dot_op_a_i[15]), .B(dot_op_b_i[11]), .ZN(n3208) );
  OAI22_X1 U3226 ( .A1(n3206), .A2(n3493), .B1(n3496), .B2(n3208), .ZN(n3319)
         );
  INV_X1 U3227 ( .A(dot_op_a_i[10]), .ZN(n3207) );
  NOR2_X1 U3228 ( .A1(n3207), .A2(n3500), .ZN(n3318) );
  XNOR2_X1 U3229 ( .A(dot_op_b_i[11]), .B(dot_op_a_i[14]), .ZN(n3304) );
  OAI22_X1 U3230 ( .A1(n3496), .A2(n3304), .B1(n3208), .B2(n3493), .ZN(n3557)
         );
  XNOR2_X1 U3231 ( .A(dot_op_b_i[7]), .B(dot_op_a_i[2]), .ZN(n3311) );
  OAI22_X1 U3232 ( .A1(n3489), .A2(n3311), .B1(n3209), .B2(n63), .ZN(n3556) );
  XNOR2_X1 U3233 ( .A(dot_op_b_i[15]), .B(dot_op_a_i[10]), .ZN(n3305) );
  OAI22_X1 U3234 ( .A1(n3510), .A2(n3305), .B1(n3210), .B2(n3534), .ZN(n3555)
         );
  XNOR2_X1 U3235 ( .A(n3212), .B(n3211), .ZN(n3322) );
  XNOR2_X1 U3236 ( .A(dot_op_b_i[13]), .B(dot_op_a_i[12]), .ZN(n3309) );
  OAI22_X1 U3237 ( .A1(n3514), .A2(n3309), .B1(n3213), .B2(n3511), .ZN(n3560)
         );
  XNOR2_X1 U3238 ( .A(dot_op_b_i[5]), .B(dot_op_a_i[4]), .ZN(n3315) );
  OAI22_X1 U3239 ( .A1(n3539), .A2(n3315), .B1(n3214), .B2(n3536), .ZN(n3559)
         );
  XNOR2_X1 U3240 ( .A(dot_op_b_i[3]), .B(dot_op_a_i[6]), .ZN(n3310) );
  OAI22_X1 U3241 ( .A1(n3551), .A2(n3310), .B1(n3215), .B2(n3549), .ZN(n3558)
         );
  FA_X1 U3242 ( .A(n3218), .B(n3217), .CI(n3216), .CO(n3196), .S(n3644) );
  FA_X1 U3243 ( .A(n3221), .B(n3220), .CI(n3219), .CO(n3326), .S(n3643) );
  FA_X1 U3244 ( .A(n3224), .B(n3223), .CI(n3222), .CO(n3191), .S(n3296) );
  FA_X1 U3245 ( .A(n3227), .B(n3226), .CI(n3225), .CO(n3192), .S(n3295) );
  INV_X1 U3246 ( .A(op_b_i[14]), .ZN(n3228) );
  NOR2_X1 U3247 ( .A1(n6118), .A2(n3228), .ZN(n3229) );
  MUX2_X1 U3248 ( .A(n3230), .B(n3229), .S(n29), .Z(n3292) );
  FA_X1 U3249 ( .A(n3233), .B(n3232), .CI(n3231), .CO(n3132), .S(n3784) );
  FA_X1 U3250 ( .A(n3236), .B(n3235), .CI(n3234), .CO(n3232), .S(n3348) );
  FA_X1 U3251 ( .A(n3239), .B(n3238), .CI(n3237), .CO(n3233), .S(n3347) );
  XNOR2_X1 U3252 ( .A(n5848), .B(n27), .ZN(n3390) );
  OAI22_X1 U3253 ( .A1(n3240), .A2(n2871), .B1(n3390), .B2(n5822), .ZN(n3342)
         );
  XNOR2_X1 U3254 ( .A(n52), .B(n5985), .ZN(n3403) );
  OAI22_X1 U3255 ( .A1(n3242), .A2(n5635), .B1(n3403), .B2(n3241), .ZN(n3341)
         );
  XNOR2_X1 U3256 ( .A(n5992), .B(n25), .ZN(n3244) );
  OAI22_X1 U3257 ( .A1(n3244), .A2(n2867), .B1(n3243), .B2(n5809), .ZN(n3615)
         );
  XNOR2_X1 U3258 ( .A(n19), .B(n25), .ZN(n3393) );
  OAI22_X1 U3259 ( .A1(n3244), .A2(n6010), .B1(n3393), .B2(n2867), .ZN(n3598)
         );
  XNOR2_X1 U3260 ( .A(n55), .B(n5919), .ZN(n3400) );
  OAI22_X1 U3261 ( .A1(n3245), .A2(n5922), .B1(n3400), .B2(n3128), .ZN(n3597)
         );
  XNOR2_X1 U3262 ( .A(n6116), .B(op_b_i[11]), .ZN(n3247) );
  OAI22_X1 U3263 ( .A1(n3247), .A2(n5943), .B1(n3246), .B2(n26), .ZN(n3596) );
  FA_X1 U3264 ( .A(n3250), .B(n3249), .CI(n3248), .CO(n3285), .S(n3782) );
  XNOR2_X1 U3265 ( .A(dot_op_b_i[21]), .B(dot_op_a_i[22]), .ZN(n3265) );
  OAI22_X1 U3266 ( .A1(n3721), .A2(n3265), .B1(n59), .B2(n3251), .ZN(n3354) );
  XNOR2_X1 U3267 ( .A(dot_op_b_i[23]), .B(dot_op_a_i[20]), .ZN(n3359) );
  OAI22_X1 U3268 ( .A1(n3469), .A2(n3359), .B1(n61), .B2(n3252), .ZN(n3352) );
  INV_X1 U3269 ( .A(dot_op_a_i[20]), .ZN(n3253) );
  NOR2_X1 U3270 ( .A1(n3253), .A2(n3448), .ZN(n3350) );
  XNOR2_X1 U3271 ( .A(dot_op_b_i[29]), .B(dot_op_a_i[30]), .ZN(n3356) );
  OAI22_X1 U3272 ( .A1(n3717), .A2(n3356), .B1(n3715), .B2(n3254), .ZN(n3366)
         );
  XNOR2_X1 U3273 ( .A(dot_op_b_i[31]), .B(dot_op_a_i[28]), .ZN(n3266) );
  OAI22_X1 U3274 ( .A1(n3474), .A2(n3266), .B1(n62), .B2(n3255), .ZN(n3365) );
  XNOR2_X1 U3275 ( .A(n3407), .B(dot_op_b_i[27]), .ZN(n3357) );
  AOI21_X1 U3276 ( .B1(n3711), .B2(n3713), .A(n3357), .ZN(n3256) );
  INV_X1 U3277 ( .A(n3256), .ZN(n3364) );
  FA_X1 U3278 ( .A(n3259), .B(n3258), .CI(n3257), .CO(n3274), .S(n3379) );
  FA_X1 U3279 ( .A(n3262), .B(n3261), .CI(n3260), .CO(n3376), .S(n3627) );
  INV_X1 U3280 ( .A(dot_op_a_i[27]), .ZN(n3263) );
  NOR2_X1 U3281 ( .A1(n3263), .A2(n3430), .ZN(n3363) );
  INV_X1 U3282 ( .A(dot_op_a_i[19]), .ZN(n3264) );
  NOR2_X1 U3283 ( .A1(n3264), .A2(n3448), .ZN(n3362) );
  XNOR2_X1 U3284 ( .A(dot_op_b_i[21]), .B(dot_op_a_i[21]), .ZN(n3374) );
  OAI22_X1 U3285 ( .A1(n3721), .A2(n3374), .B1(n59), .B2(n3265), .ZN(n3371) );
  XNOR2_X1 U3286 ( .A(dot_op_b_i[31]), .B(dot_op_a_i[27]), .ZN(n3369) );
  OAI22_X1 U3287 ( .A1(n3474), .A2(n3369), .B1(n62), .B2(n3266), .ZN(n3370) );
  OR2_X1 U3288 ( .A1(n3371), .A2(n3370), .ZN(n3361) );
  FA_X1 U3289 ( .A(n3269), .B(n3268), .CI(n3267), .CO(n3377), .S(n3625) );
  FA_X1 U3290 ( .A(n3272), .B(n3271), .CI(n3270), .CO(n3288), .S(n3786) );
  FA_X1 U3291 ( .A(n3275), .B(n3274), .CI(n3273), .CO(n3289), .S(n3785) );
  MUX2_X1 U3292 ( .A(n3277), .B(n3276), .S(n6142), .Z(n3383) );
  FA_X1 U3293 ( .A(n3280), .B(n3279), .CI(n3278), .CO(n3160), .S(n3281) );
  NOR2_X1 U3294 ( .A1(n4071), .A2(n4070), .ZN(n4901) );
  FA_X1 U3295 ( .A(n3283), .B(n3282), .CI(n3281), .CO(n4070), .S(n4069) );
  FA_X1 U3296 ( .A(n3286), .B(n3285), .CI(n3284), .CO(n3146), .S(n3291) );
  FA_X1 U3297 ( .A(n3289), .B(n3288), .CI(n3287), .CO(n3185), .S(n3290) );
  MUX2_X1 U3298 ( .A(n3291), .B(n3290), .S(n6144), .Z(n3778) );
  FA_X1 U3299 ( .A(n3294), .B(n3293), .CI(n3292), .CO(n3384), .S(n3792) );
  FA_X1 U3300 ( .A(n3297), .B(n3296), .CI(n3295), .CO(n3230), .S(n3298) );
  AND2_X1 U3301 ( .A1(n3298), .A2(n6144), .ZN(n3761) );
  INV_X1 U3302 ( .A(op_c_i[13]), .ZN(n3299) );
  OAI22_X1 U3303 ( .A1(n6112), .A2(n3300), .B1(n2525), .B2(n3299), .ZN(n3760)
         );
  FA_X1 U3304 ( .A(n3303), .B(n3302), .CI(n3301), .CO(n3328), .S(n3647) );
  NOR2_X1 U3305 ( .A1(n1313), .A2(n3500), .ZN(n3520) );
  XNOR2_X1 U3306 ( .A(dot_op_a_i[13]), .B(dot_op_b_i[11]), .ZN(n3494) );
  OAI22_X1 U3307 ( .A1(n3496), .A2(n3494), .B1(n3493), .B2(n3304), .ZN(n3503)
         );
  XNOR2_X1 U3308 ( .A(dot_op_a_i[9]), .B(dot_op_b_i[15]), .ZN(n3508) );
  OAI22_X1 U3309 ( .A1(n3510), .A2(n3508), .B1(n3305), .B2(n3534), .ZN(n3502)
         );
  NOR2_X1 U3310 ( .A1(n1628), .A2(n3316), .ZN(n3518) );
  FA_X1 U3311 ( .A(n3308), .B(n3307), .CI(n3306), .CO(n3302), .S(n3581) );
  XNOR2_X1 U3312 ( .A(dot_op_a_i[11]), .B(dot_op_b_i[13]), .ZN(n3512) );
  OAI22_X1 U3313 ( .A1(n3514), .A2(n3512), .B1(n3511), .B2(n3309), .ZN(n3531)
         );
  XNOR2_X1 U3314 ( .A(dot_op_a_i[5]), .B(dot_op_b_i[3]), .ZN(n3486) );
  OAI22_X1 U3315 ( .A1(n3551), .A2(n3486), .B1(n3549), .B2(n3310), .ZN(n3530)
         );
  XNOR2_X1 U3316 ( .A(dot_op_a_i[1]), .B(dot_op_b_i[7]), .ZN(n3487) );
  OAI22_X1 U3317 ( .A1(n3489), .A2(n3487), .B1(n3311), .B2(n63), .ZN(n3529) );
  XNOR2_X1 U3318 ( .A(n3312), .B(dot_op_b_i[9]), .ZN(n3499) );
  AOI21_X1 U3319 ( .B1(n3547), .B2(n3544), .A(n3499), .ZN(n3313) );
  INV_X1 U3320 ( .A(n3313), .ZN(n3553) );
  XNOR2_X1 U3321 ( .A(n3314), .B(dot_op_b_i[1]), .ZN(n3521) );
  XNOR2_X1 U3322 ( .A(dot_op_a_i[7]), .B(dot_op_b_i[1]), .ZN(n3497) );
  OAI22_X1 U3323 ( .A1(n3521), .A2(n3540), .B1(n3543), .B2(n3497), .ZN(n3528)
         );
  XNOR2_X1 U3324 ( .A(dot_op_a_i[3]), .B(dot_op_b_i[5]), .ZN(n3537) );
  OAI22_X1 U3325 ( .A1(n3539), .A2(n3537), .B1(n3536), .B2(n3315), .ZN(n3527)
         );
  INV_X1 U3326 ( .A(n3316), .ZN(n3317) );
  AND2_X1 U3327 ( .A1(dot_op_a_i[0]), .A2(n3317), .ZN(n3526) );
  FA_X1 U3328 ( .A(n3320), .B(n3319), .CI(n3318), .CO(n3301), .S(n3573) );
  FA_X1 U3329 ( .A(n3323), .B(n3322), .CI(n3321), .CO(n3645), .S(n3572) );
  FA_X1 U3330 ( .A(n3326), .B(n3325), .CI(n3324), .CO(n3225), .S(n3658) );
  FA_X1 U3331 ( .A(n3329), .B(n3328), .CI(n3327), .CO(n3297), .S(n3657) );
  INV_X1 U3332 ( .A(op_b_i[13]), .ZN(n3330) );
  NOR2_X1 U3333 ( .A1(n6118), .A2(n3330), .ZN(n3331) );
  MUX2_X1 U3334 ( .A(n3332), .B(n3331), .S(n29), .Z(n3759) );
  FA_X1 U3335 ( .A(n3335), .B(n3334), .CI(n3333), .CO(n3343), .S(n3622) );
  FA_X1 U3336 ( .A(n3338), .B(n3337), .CI(n3336), .CO(n3345), .S(n3621) );
  OR2_X1 U3337 ( .A1(n6116), .A2(n3636), .ZN(n3339) );
  OAI22_X1 U3338 ( .A1(n3339), .A2(n26), .B1(n5943), .B2(n3636), .ZN(n3589) );
  XNOR2_X1 U3339 ( .A(n20), .B(n6015), .ZN(n3391) );
  OAI22_X1 U3340 ( .A1(n3340), .A2(n10), .B1(n3391), .B2(n2585), .ZN(n3588) );
  HA_X1 U3341 ( .A(n3342), .B(n3341), .CO(n3616), .S(n3587) );
  FA_X1 U3342 ( .A(n3345), .B(n3344), .CI(n3343), .CO(n3248), .S(n3752) );
  FA_X1 U3343 ( .A(n3348), .B(n3347), .CI(n3346), .CO(n3783), .S(n3751) );
  FA_X1 U3344 ( .A(n3351), .B(n3350), .CI(n3349), .CO(n3380), .S(n3630) );
  FA_X1 U3345 ( .A(n3354), .B(n3353), .CI(n3352), .CO(n3351), .S(n3606) );
  XNOR2_X1 U3346 ( .A(dot_op_b_i[19]), .B(dot_op_a_i[23]), .ZN(n3373) );
  OAI22_X1 U3347 ( .A1(n3465), .A2(n3373), .B1(n3355), .B2(n60), .ZN(n3452) );
  XNOR2_X1 U3348 ( .A(dot_op_b_i[29]), .B(dot_op_a_i[29]), .ZN(n3367) );
  OAI22_X1 U3349 ( .A1(n3717), .A2(n3367), .B1(n3715), .B2(n3356), .ZN(n3451)
         );
  XNOR2_X1 U3350 ( .A(dot_op_b_i[27]), .B(dot_op_a_i[31]), .ZN(n3372) );
  OAI22_X1 U3351 ( .A1(n3713), .A2(n3372), .B1(n3357), .B2(n3711), .ZN(n3450)
         );
  INV_X1 U3352 ( .A(dot_op_a_i[18]), .ZN(n3358) );
  NOR2_X1 U3353 ( .A1(n3358), .A2(n3448), .ZN(n3440) );
  XNOR2_X1 U3354 ( .A(dot_op_b_i[23]), .B(dot_op_a_i[19]), .ZN(n3368) );
  OAI22_X1 U3355 ( .A1(n3469), .A2(n3368), .B1(n61), .B2(n3359), .ZN(n3439) );
  INV_X1 U3356 ( .A(dot_op_a_i[26]), .ZN(n3360) );
  NOR2_X1 U3357 ( .A1(n3360), .A2(n3430), .ZN(n3438) );
  FA_X1 U3358 ( .A(n3363), .B(n3362), .CI(n3361), .CO(n3626), .S(n3603) );
  FA_X1 U3359 ( .A(n3366), .B(n3365), .CI(n3364), .CO(n3349), .S(n3602) );
  XNOR2_X1 U3360 ( .A(dot_op_b_i[29]), .B(dot_op_a_i[28]), .ZN(n3433) );
  OAI22_X1 U3361 ( .A1(n3717), .A2(n3433), .B1(n3715), .B2(n3367), .ZN(n3426)
         );
  XNOR2_X1 U3362 ( .A(dot_op_b_i[23]), .B(dot_op_a_i[18]), .ZN(n3409) );
  OAI22_X1 U3363 ( .A1(n3469), .A2(n3409), .B1(n61), .B2(n3368), .ZN(n3425) );
  XNOR2_X1 U3364 ( .A(dot_op_b_i[31]), .B(dot_op_a_i[26]), .ZN(n3434) );
  OAI22_X1 U3365 ( .A1(n3474), .A2(n3434), .B1(n62), .B2(n3369), .ZN(n3424) );
  XNOR2_X1 U3366 ( .A(n3371), .B(n3370), .ZN(n3442) );
  XNOR2_X1 U3367 ( .A(dot_op_b_i[27]), .B(dot_op_a_i[30]), .ZN(n3410) );
  OAI22_X1 U3368 ( .A1(n3713), .A2(n3410), .B1(n3711), .B2(n3372), .ZN(n3429)
         );
  XNOR2_X1 U3369 ( .A(dot_op_b_i[19]), .B(dot_op_a_i[22]), .ZN(n3406) );
  OAI22_X1 U3370 ( .A1(n3465), .A2(n3406), .B1(n60), .B2(n3373), .ZN(n3428) );
  XNOR2_X1 U3371 ( .A(dot_op_b_i[21]), .B(dot_op_a_i[20]), .ZN(n3408) );
  OAI22_X1 U3372 ( .A1(n3721), .A2(n3408), .B1(n59), .B2(n3374), .ZN(n3427) );
  FA_X1 U3373 ( .A(n3377), .B(n3376), .CI(n3375), .CO(n3273), .S(n3755) );
  FA_X1 U3374 ( .A(n3380), .B(n3379), .CI(n3378), .CO(n3787), .S(n3754) );
  MUX2_X1 U3375 ( .A(n3382), .B(n3381), .S(n6117), .Z(n3790) );
  FA_X1 U3376 ( .A(n3385), .B(n3384), .CI(n3383), .CO(n3282), .S(n3776) );
  NOR2_X1 U3377 ( .A1(n4069), .A2(n4068), .ZN(n4899) );
  NOR2_X1 U3378 ( .A1(n4901), .A2(n4899), .ZN(n4928) );
  NAND2_X1 U3379 ( .A1(n4077), .A2(n4928), .ZN(n4079) );
  INV_X1 U3380 ( .A(n2472), .ZN(n4342) );
  XNOR2_X1 U3381 ( .A(n5992), .B(n4342), .ZN(n3392) );
  XNOR2_X1 U3382 ( .A(n19), .B(n4342), .ZN(n3701) );
  OAI22_X1 U3383 ( .A1(n3392), .A2(n10), .B1(n3701), .B2(n2585), .ZN(n3399) );
  XNOR2_X1 U3384 ( .A(n21), .B(n4337), .ZN(n3404) );
  XNOR2_X1 U3385 ( .A(n20), .B(n5985), .ZN(n3389) );
  OAI22_X1 U3386 ( .A1(n3404), .A2(n5635), .B1(n3389), .B2(n3241), .ZN(n3398)
         );
  OR2_X1 U3387 ( .A1(n6116), .A2(n3386), .ZN(n3387) );
  OAI22_X1 U3388 ( .A1(n3387), .A2(n2871), .B1(n5822), .B2(n3386), .ZN(n3705)
         );
  XNOR2_X1 U3389 ( .A(n56), .B(n25), .ZN(n3702) );
  XNOR2_X1 U3390 ( .A(n55), .B(n25), .ZN(n3394) );
  OAI22_X1 U3391 ( .A1(n3702), .A2(n2867), .B1(n3394), .B2(n5809), .ZN(n3828)
         );
  AND2_X1 U3392 ( .A1(n6116), .A2(n3388), .ZN(n3827) );
  INV_X1 U3393 ( .A(n2527), .ZN(n4337) );
  XNOR2_X1 U3394 ( .A(n54), .B(n4337), .ZN(n3830) );
  OAI22_X1 U3395 ( .A1(n3830), .A2(n3241), .B1(n3389), .B2(n5635), .ZN(n3826)
         );
  XNOR2_X1 U3396 ( .A(n6002), .B(n27), .ZN(n3396) );
  OAI22_X1 U3397 ( .A1(n3396), .A2(n5822), .B1(n3390), .B2(n4546), .ZN(n3592)
         );
  OAI22_X1 U3398 ( .A1(n3392), .A2(n2585), .B1(n3391), .B2(n10), .ZN(n3591) );
  XNOR2_X1 U3399 ( .A(n22), .B(n25), .ZN(n3395) );
  OAI22_X1 U3400 ( .A1(n3395), .A2(n2867), .B1(n3393), .B2(n5809), .ZN(n3590)
         );
  XNOR2_X1 U3401 ( .A(n56), .B(n5919), .ZN(n3401) );
  XNOR2_X1 U3402 ( .A(n5848), .B(n5919), .ZN(n3700) );
  OAI22_X1 U3403 ( .A1(n3401), .A2(n5922), .B1(n3700), .B2(n3128), .ZN(n3699)
         );
  OAI22_X1 U3404 ( .A1(n3395), .A2(n6010), .B1(n3394), .B2(n2867), .ZN(n3698)
         );
  XNOR2_X1 U3405 ( .A(n6116), .B(n27), .ZN(n3397) );
  OAI22_X1 U3406 ( .A1(n3397), .A2(n5822), .B1(n3396), .B2(n4546), .ZN(n3697)
         );
  HA_X1 U3407 ( .A(n3399), .B(n3398), .CO(n3585), .S(n3706) );
  OAI22_X1 U3408 ( .A1(n3401), .A2(n3128), .B1(n3400), .B2(n5922), .ZN(n3595)
         );
  AND2_X1 U3409 ( .A1(n6116), .A2(n3402), .ZN(n3594) );
  OAI22_X1 U3410 ( .A1(n3404), .A2(n3241), .B1(n3403), .B2(n5635), .ZN(n3593)
         );
  XNOR2_X1 U3411 ( .A(dot_op_b_i[17]), .B(dot_op_a_i[23]), .ZN(n3477) );
  XNOR2_X1 U3412 ( .A(n3405), .B(dot_op_b_i[17]), .ZN(n3446) );
  OAI22_X1 U3413 ( .A1(n3479), .A2(n3477), .B1(n3446), .B2(n1662), .ZN(n3419)
         );
  XNOR2_X1 U3414 ( .A(dot_op_b_i[19]), .B(dot_op_a_i[21]), .ZN(n3462) );
  OAI22_X1 U3415 ( .A1(n3465), .A2(n3462), .B1(n60), .B2(n3406), .ZN(n3418) );
  XNOR2_X1 U3416 ( .A(dot_op_b_i[25]), .B(dot_op_a_i[31]), .ZN(n3480) );
  XNOR2_X1 U3417 ( .A(n3407), .B(dot_op_b_i[25]), .ZN(n3444) );
  OAI22_X1 U3418 ( .A1(n3482), .A2(n3480), .B1(n3444), .B2(n1312), .ZN(n3417)
         );
  XNOR2_X1 U3419 ( .A(dot_op_b_i[21]), .B(dot_op_a_i[19]), .ZN(n3413) );
  OAI22_X1 U3420 ( .A1(n3721), .A2(n3413), .B1(n59), .B2(n3408), .ZN(n3423) );
  XNOR2_X1 U3421 ( .A(dot_op_b_i[23]), .B(dot_op_a_i[17]), .ZN(n3466) );
  OAI22_X1 U3422 ( .A1(n3469), .A2(n3466), .B1(n61), .B2(n3409), .ZN(n3422) );
  XNOR2_X1 U3423 ( .A(dot_op_b_i[27]), .B(dot_op_a_i[29]), .ZN(n3476) );
  OAI22_X1 U3424 ( .A1(n3713), .A2(n3476), .B1(n3711), .B2(n3410), .ZN(n3421)
         );
  INV_X1 U3425 ( .A(n3467), .ZN(n3411) );
  AND2_X1 U3426 ( .A1(dot_op_a_i[16]), .A2(n3411), .ZN(n3843) );
  INV_X1 U3427 ( .A(n62), .ZN(n3412) );
  AND2_X1 U3428 ( .A1(dot_op_a_i[24]), .A2(n3412), .ZN(n3842) );
  XNOR2_X1 U3429 ( .A(dot_op_b_i[21]), .B(dot_op_a_i[18]), .ZN(n3718) );
  OAI22_X1 U3430 ( .A1(n3721), .A2(n3718), .B1(n59), .B2(n3413), .ZN(n3851) );
  XNOR2_X1 U3431 ( .A(dot_op_b_i[17]), .B(dot_op_a_i[22]), .ZN(n3478) );
  OAI22_X1 U3432 ( .A1(n3479), .A2(n3414), .B1(n3478), .B2(n1662), .ZN(n3919)
         );
  XNOR2_X1 U3433 ( .A(dot_op_b_i[25]), .B(dot_op_a_i[30]), .ZN(n3481) );
  OAI22_X1 U3434 ( .A1(n3482), .A2(n3415), .B1(n3481), .B2(n1312), .ZN(n3918)
         );
  XNOR2_X1 U3435 ( .A(dot_op_b_i[19]), .B(dot_op_a_i[20]), .ZN(n3464) );
  OAI22_X1 U3436 ( .A1(n3465), .A2(n3416), .B1(n60), .B2(n3464), .ZN(n3917) );
  FA_X1 U3437 ( .A(n3419), .B(n3418), .CI(n3417), .CO(n3437), .S(n3838) );
  INV_X1 U3438 ( .A(dot_op_a_i[25]), .ZN(n3420) );
  NOR2_X1 U3439 ( .A1(n3420), .A2(n3430), .ZN(n3436) );
  FA_X1 U3440 ( .A(n3423), .B(n3422), .CI(n3421), .CO(n3435), .S(n3837) );
  FA_X1 U3441 ( .A(n3426), .B(n3425), .CI(n3424), .CO(n3443), .S(n3455) );
  FA_X1 U3442 ( .A(n3429), .B(n3428), .CI(n3427), .CO(n3441), .S(n3454) );
  INV_X1 U3443 ( .A(n3430), .ZN(n3431) );
  AND2_X1 U3444 ( .A1(dot_op_a_i[24]), .A2(n3431), .ZN(n3727) );
  INV_X1 U3445 ( .A(n3448), .ZN(n3432) );
  AND2_X1 U3446 ( .A1(dot_op_a_i[16]), .A2(n3432), .ZN(n3726) );
  XNOR2_X1 U3447 ( .A(dot_op_b_i[29]), .B(dot_op_a_i[27]), .ZN(n3475) );
  OAI22_X1 U3448 ( .A1(n3717), .A2(n3475), .B1(n3715), .B2(n3433), .ZN(n3457)
         );
  XNOR2_X1 U3449 ( .A(dot_op_b_i[31]), .B(dot_op_a_i[25]), .ZN(n3471) );
  OAI22_X1 U3450 ( .A1(n3474), .A2(n3471), .B1(n62), .B2(n3434), .ZN(n3456) );
  FA_X1 U3451 ( .A(n3437), .B(n3436), .CI(n3435), .CO(n3611), .S(n3735) );
  FA_X1 U3452 ( .A(n3440), .B(n3439), .CI(n3438), .CO(n3604), .S(n3610) );
  FA_X1 U3453 ( .A(n3443), .B(n3442), .CI(n3441), .CO(n3601), .S(n3609) );
  AOI21_X1 U3454 ( .B1(n3482), .B2(n1312), .A(n3444), .ZN(n3445) );
  INV_X1 U3455 ( .A(n3445), .ZN(n3460) );
  AOI21_X1 U3456 ( .B1(n3479), .B2(n1662), .A(n3446), .ZN(n3447) );
  INV_X1 U3457 ( .A(n3447), .ZN(n3459) );
  INV_X1 U3458 ( .A(dot_op_a_i[17]), .ZN(n3449) );
  NOR2_X1 U3459 ( .A1(n3449), .A2(n3448), .ZN(n3458) );
  FA_X1 U3460 ( .A(n3452), .B(n3451), .CI(n3450), .CO(n3605), .S(n3607) );
  FA_X1 U3461 ( .A(n3455), .B(n3454), .CI(n3453), .CO(n3600), .S(n3734) );
  HA_X1 U3462 ( .A(n3457), .B(n3456), .CO(n3733), .S(n3725) );
  FA_X1 U3463 ( .A(n3460), .B(n3459), .CI(n3458), .CO(n3608), .S(n3732) );
  OR2_X1 U3464 ( .A1(dot_op_a_i[16]), .A2(n2929), .ZN(n3461) );
  OAI22_X1 U3465 ( .A1(n3469), .A2(n2929), .B1(n3461), .B2(n61), .ZN(n3709) );
  OAI22_X1 U3466 ( .A1(n3465), .A2(n3464), .B1(n60), .B2(n3462), .ZN(n3708) );
  XNOR2_X1 U3467 ( .A(dot_op_b_i[23]), .B(dot_op_a_i[16]), .ZN(n3468) );
  OAI22_X1 U3468 ( .A1(n3469), .A2(n3468), .B1(n61), .B2(n3466), .ZN(n3707) );
  OR2_X1 U3469 ( .A1(dot_op_a_i[24]), .A2(n2925), .ZN(n3470) );
  OAI22_X1 U3470 ( .A1(n3474), .A2(n2925), .B1(n3470), .B2(n62), .ZN(n3849) );
  XNOR2_X1 U3471 ( .A(dot_op_b_i[31]), .B(dot_op_a_i[24]), .ZN(n3473) );
  OAI22_X1 U3472 ( .A1(n3474), .A2(n3473), .B1(n62), .B2(n3471), .ZN(n3848) );
  XNOR2_X1 U3473 ( .A(dot_op_b_i[29]), .B(dot_op_a_i[26]), .ZN(n3714) );
  OAI22_X1 U3474 ( .A1(n3717), .A2(n3714), .B1(n3715), .B2(n3475), .ZN(n3847)
         );
  XNOR2_X1 U3475 ( .A(dot_op_b_i[27]), .B(dot_op_a_i[28]), .ZN(n3710) );
  OAI22_X1 U3476 ( .A1(n3713), .A2(n3710), .B1(n3711), .B2(n3476), .ZN(n3724)
         );
  OAI22_X1 U3477 ( .A1(n3479), .A2(n3478), .B1(n3477), .B2(n1662), .ZN(n3723)
         );
  OAI22_X1 U3478 ( .A1(n3482), .A2(n3481), .B1(n3480), .B2(n1312), .ZN(n3722)
         );
  MUX2_X1 U3479 ( .A(n3484), .B(n3483), .S(n6145), .Z(n3747) );
  OR2_X1 U3480 ( .A1(dot_op_a_i[0]), .A2(n2836), .ZN(n3485) );
  OAI22_X1 U3481 ( .A1(n3489), .A2(n2836), .B1(n3485), .B2(n63), .ZN(n3506) );
  XNOR2_X1 U3482 ( .A(dot_op_b_i[3]), .B(dot_op_a_i[4]), .ZN(n3548) );
  OAI22_X1 U3483 ( .A1(n3551), .A2(n3548), .B1(n3486), .B2(n3549), .ZN(n3505)
         );
  XNOR2_X1 U3484 ( .A(dot_op_b_i[7]), .B(dot_op_a_i[0]), .ZN(n3488) );
  OAI22_X1 U3485 ( .A1(n3489), .A2(n3488), .B1(n3487), .B2(n63), .ZN(n3504) );
  XNOR2_X1 U3486 ( .A(dot_op_b_i[11]), .B(dot_op_a_i[12]), .ZN(n3495) );
  OAI22_X1 U3487 ( .A1(n3496), .A2(n3490), .B1(n3493), .B2(n3495), .ZN(n3807)
         );
  XNOR2_X1 U3488 ( .A(dot_op_b_i[13]), .B(dot_op_a_i[10]), .ZN(n3513) );
  OAI22_X1 U3489 ( .A1(n3514), .A2(n3491), .B1(n3511), .B2(n3513), .ZN(n3806)
         );
  XNOR2_X1 U3490 ( .A(dot_op_b_i[5]), .B(dot_op_a_i[2]), .ZN(n3538) );
  OAI22_X1 U3491 ( .A1(n3539), .A2(n3492), .B1(n3536), .B2(n3538), .ZN(n3805)
         );
  OAI22_X1 U3492 ( .A1(n3496), .A2(n3495), .B1(n3494), .B2(n3493), .ZN(n3517)
         );
  XNOR2_X1 U3493 ( .A(dot_op_b_i[1]), .B(dot_op_a_i[6]), .ZN(n3541) );
  OAI22_X1 U3494 ( .A1(n3543), .A2(n3541), .B1(n3497), .B2(n3540), .ZN(n3516)
         );
  XNOR2_X1 U3495 ( .A(dot_op_b_i[9]), .B(dot_op_a_i[14]), .ZN(n3545) );
  XNOR2_X1 U3496 ( .A(dot_op_a_i[15]), .B(dot_op_b_i[9]), .ZN(n3498) );
  OAI22_X1 U3497 ( .A1(n3547), .A2(n3545), .B1(n3498), .B2(n3544), .ZN(n3515)
         );
  OAI22_X1 U3498 ( .A1(n3499), .A2(n3544), .B1(n3547), .B2(n3498), .ZN(n3563)
         );
  INV_X1 U3499 ( .A(n3500), .ZN(n3501) );
  AND2_X1 U3500 ( .A1(dot_op_a_i[8]), .A2(n3501), .ZN(n3562) );
  HA_X1 U3501 ( .A(n3503), .B(n3502), .CO(n3519), .S(n3561) );
  FA_X1 U3502 ( .A(n3506), .B(n3505), .CI(n3504), .CO(n3525), .S(n3804) );
  OR2_X1 U3503 ( .A1(dot_op_a_i[8]), .A2(n2833), .ZN(n3507) );
  OAI22_X1 U3504 ( .A1(n3510), .A2(n2833), .B1(n3507), .B2(n3534), .ZN(n3682)
         );
  XNOR2_X1 U3505 ( .A(dot_op_b_i[15]), .B(dot_op_a_i[8]), .ZN(n3509) );
  OAI22_X1 U3506 ( .A1(n3510), .A2(n3509), .B1(n3508), .B2(n3534), .ZN(n3681)
         );
  OAI22_X1 U3507 ( .A1(n3514), .A2(n3513), .B1(n3512), .B2(n3511), .ZN(n3680)
         );
  FA_X1 U3508 ( .A(n3517), .B(n3516), .CI(n3515), .CO(n3523), .S(n3802) );
  FA_X1 U3509 ( .A(n3520), .B(n3519), .CI(n3518), .CO(n3582), .S(n3577) );
  AOI21_X1 U3510 ( .B1(n3543), .B2(n3540), .A(n3521), .ZN(n3522) );
  INV_X1 U3511 ( .A(n3522), .ZN(n3576) );
  FA_X1 U3512 ( .A(n3525), .B(n3524), .CI(n3523), .CO(n3575), .S(n3686) );
  FA_X1 U3513 ( .A(n3528), .B(n3527), .CI(n3526), .CO(n3552), .S(n3671) );
  FA_X1 U3514 ( .A(n3531), .B(n3530), .CI(n3529), .CO(n3554), .S(n3670) );
  INV_X1 U3515 ( .A(n3532), .ZN(n3533) );
  AND2_X1 U3516 ( .A1(dot_op_a_i[0]), .A2(n3533), .ZN(n3676) );
  INV_X1 U3517 ( .A(n3534), .ZN(n3535) );
  AND2_X1 U3518 ( .A1(dot_op_a_i[8]), .A2(n3535), .ZN(n3675) );
  OAI22_X1 U3519 ( .A1(n3539), .A2(n3538), .B1(n3537), .B2(n3536), .ZN(n3684)
         );
  OAI22_X1 U3520 ( .A1(n3543), .A2(n3542), .B1(n3541), .B2(n3540), .ZN(n3813)
         );
  OAI22_X1 U3521 ( .A1(n3547), .A2(n3546), .B1(n3545), .B2(n3544), .ZN(n3812)
         );
  OAI22_X1 U3522 ( .A1(n3551), .A2(n3550), .B1(n3549), .B2(n3548), .ZN(n3811)
         );
  FA_X1 U3523 ( .A(n3554), .B(n3553), .CI(n3552), .CO(n3574), .S(n3570) );
  FA_X1 U3524 ( .A(n3557), .B(n3556), .CI(n3555), .CO(n3323), .S(n3580) );
  FA_X1 U3525 ( .A(n3560), .B(n3559), .CI(n3558), .CO(n3321), .S(n3579) );
  FA_X1 U3526 ( .A(n3563), .B(n3562), .CI(n3561), .CO(n3578), .S(n3687) );
  INV_X1 U3527 ( .A(op_b_i[10]), .ZN(n3564) );
  NOR2_X1 U3528 ( .A1(n6118), .A2(n3564), .ZN(n3565) );
  MUX2_X1 U3529 ( .A(n3566), .B(n3565), .S(n29), .Z(n3741) );
  INV_X1 U3530 ( .A(op_c_i[10]), .ZN(n3567) );
  OAI22_X1 U3531 ( .A1(n6146), .A2(n3568), .B1(n2525), .B2(n3567), .ZN(n3740)
         );
  FA_X1 U3532 ( .A(n3571), .B(n3570), .CI(n3569), .CO(n3635), .S(n3693) );
  FA_X1 U3533 ( .A(n3574), .B(n3573), .CI(n3572), .CO(n3646), .S(n3634) );
  FA_X1 U3534 ( .A(n3577), .B(n3576), .CI(n3575), .CO(n3642), .S(n3694) );
  FA_X1 U3535 ( .A(n3580), .B(n3579), .CI(n3578), .CO(n3641), .S(n3569) );
  AND2_X1 U3536 ( .A1(n3583), .A2(n6144), .ZN(n3739) );
  FA_X1 U3537 ( .A(n3586), .B(n3585), .CI(n3584), .CO(n3651), .S(n3866) );
  FA_X1 U3538 ( .A(n3589), .B(n3588), .CI(n3587), .CO(n3620), .S(n3650) );
  FA_X1 U3539 ( .A(n3592), .B(n3591), .CI(n3590), .CO(n3619), .S(n3867) );
  FA_X1 U3540 ( .A(n3595), .B(n3594), .CI(n3593), .CO(n3618), .S(n3584) );
  FA_X1 U3541 ( .A(n3598), .B(n3597), .CI(n3596), .CO(n3614), .S(n3617) );
  FA_X1 U3542 ( .A(n104), .B(n3600), .CI(n3599), .CO(n3654), .S(n3869) );
  FA_X1 U3543 ( .A(n3603), .B(n3602), .CI(n3601), .CO(n3628), .S(n3653) );
  FA_X1 U3544 ( .A(n3606), .B(n3605), .CI(n3604), .CO(n3629), .S(n3624) );
  FA_X1 U3545 ( .A(n3611), .B(n3610), .CI(n3609), .CO(n3623), .S(n3870) );
  MUX2_X1 U3546 ( .A(n3613), .B(n3612), .S(n6117), .Z(n3745) );
  FA_X1 U3547 ( .A(n3616), .B(n3615), .CI(n3614), .CO(n3346), .S(n3767) );
  FA_X1 U3548 ( .A(n3619), .B(n3618), .CI(n3617), .CO(n3766), .S(n3649) );
  FA_X1 U3549 ( .A(n3622), .B(n3621), .CI(n3620), .CO(n3753), .S(n3765) );
  FA_X1 U3550 ( .A(n3624), .B(n103), .CI(n3623), .CO(n3770), .S(n3652) );
  FA_X1 U3551 ( .A(n3627), .B(n3626), .CI(n3625), .CO(n3378), .S(n3769) );
  FA_X1 U3552 ( .A(n3630), .B(n3629), .CI(n3628), .CO(n3756), .S(n3768) );
  MUX2_X1 U3553 ( .A(n3632), .B(n3631), .S(n6144), .Z(n3774) );
  FA_X1 U3554 ( .A(n3635), .B(n3634), .CI(n3633), .CO(n3638), .S(n3583) );
  INV_X1 U3555 ( .A(op_b_i[11]), .ZN(n3636) );
  NOR2_X1 U3556 ( .A1(n6119), .A2(n3636), .ZN(n3637) );
  MUX2_X1 U3557 ( .A(n3638), .B(n3637), .S(n29), .Z(n3744) );
  INV_X1 U3558 ( .A(op_c_i[11]), .ZN(n3639) );
  OAI22_X1 U3559 ( .A1(n6146), .A2(n3640), .B1(n2525), .B2(n3639), .ZN(n3743)
         );
  FA_X1 U3560 ( .A(n3642), .B(n3641), .CI(n100), .CO(n3665), .S(n3633) );
  FA_X1 U3561 ( .A(n3645), .B(n3644), .CI(n3643), .CO(n3327), .S(n3664) );
  FA_X1 U3562 ( .A(n3647), .B(n99), .CI(n3646), .CO(n3659), .S(n3663) );
  AND2_X1 U3563 ( .A1(n3648), .A2(n6145), .ZN(n3742) );
  FA_X1 U3564 ( .A(n3651), .B(n3650), .CI(n3649), .CO(n3656), .S(n3613) );
  FA_X1 U3565 ( .A(n3654), .B(n3653), .CI(n3652), .CO(n3655), .S(n3612) );
  MUX2_X1 U3566 ( .A(n3656), .B(n3655), .S(n6144), .Z(n3749) );
  FA_X1 U3567 ( .A(n3659), .B(n3658), .CI(n3657), .CO(n3332), .S(n3660) );
  AND2_X1 U3568 ( .A1(n3660), .A2(n6144), .ZN(n3764) );
  INV_X1 U3569 ( .A(op_c_i[12]), .ZN(n3661) );
  OAI22_X1 U3570 ( .A1(n6112), .A2(n3662), .B1(n2525), .B2(n3661), .ZN(n3763)
         );
  FA_X1 U3571 ( .A(n3665), .B(n3664), .CI(n3663), .CO(n3668), .S(n3648) );
  INV_X1 U3572 ( .A(op_b_i[12]), .ZN(n3666) );
  NOR2_X1 U3573 ( .A1(n6118), .A2(n3666), .ZN(n3667) );
  MUX2_X1 U3574 ( .A(n3668), .B(n3667), .S(n29), .Z(n3762) );
  FA_X1 U3575 ( .A(n3671), .B(n3670), .CI(n3669), .CO(n3571), .S(n3824) );
  FA_X1 U3576 ( .A(n3674), .B(n3673), .CI(n3672), .CO(n3885), .S(n3880) );
  HA_X1 U3577 ( .A(n3676), .B(n3675), .CO(n3685), .S(n3884) );
  FA_X1 U3578 ( .A(n3679), .B(n3678), .CI(n3677), .CO(n3883), .S(n3882) );
  FA_X1 U3579 ( .A(n3682), .B(n3681), .CI(n3680), .CO(n3524), .S(n3815) );
  FA_X1 U3580 ( .A(n3685), .B(n3684), .CI(n3683), .CO(n3669), .S(n3814) );
  FA_X1 U3581 ( .A(n3688), .B(n3687), .CI(n3686), .CO(n3695), .S(n3822) );
  NOR2_X1 U3582 ( .A1(n6118), .A2(n3386), .ZN(n3689) );
  MUX2_X1 U3583 ( .A(n3690), .B(n3689), .S(n29), .Z(n3935) );
  INV_X1 U3584 ( .A(op_c_i[9]), .ZN(n3691) );
  OAI22_X1 U3585 ( .A1(n6146), .A2(n3692), .B1(n2525), .B2(n3691), .ZN(n3934)
         );
  FA_X1 U3586 ( .A(n3695), .B(n3694), .CI(n3693), .CO(n3566), .S(n3696) );
  AND2_X1 U3587 ( .A1(n3696), .A2(n6143), .ZN(n3933) );
  FA_X1 U3588 ( .A(n3699), .B(n3698), .CI(n3697), .CO(n3586), .S(n3860) );
  XNOR2_X1 U3589 ( .A(n6002), .B(n5919), .ZN(n3831) );
  OAI22_X1 U3590 ( .A1(n3831), .A2(n3128), .B1(n3700), .B2(n5922), .ZN(n3835)
         );
  XNOR2_X1 U3591 ( .A(n22), .B(n4342), .ZN(n3703) );
  OAI22_X1 U3592 ( .A1(n3703), .A2(n2585), .B1(n3701), .B2(n10), .ZN(n3834) );
  XNOR2_X1 U3593 ( .A(n5848), .B(n25), .ZN(n3941) );
  OAI22_X1 U3594 ( .A1(n3702), .A2(n5809), .B1(n3941), .B2(n2867), .ZN(n3904)
         );
  XNOR2_X1 U3595 ( .A(n55), .B(n4342), .ZN(n3901) );
  OAI22_X1 U3596 ( .A1(n3703), .A2(n10), .B1(n3901), .B2(n2585), .ZN(n3903) );
  FA_X1 U3597 ( .A(n3706), .B(n3705), .CI(n3704), .CO(n3868), .S(n3858) );
  FA_X1 U3598 ( .A(n3709), .B(n3708), .CI(n3707), .CO(n3730), .S(n3910) );
  OAI22_X1 U3599 ( .A1(n3713), .A2(n3712), .B1(n3711), .B2(n3710), .ZN(n3913)
         );
  OAI22_X1 U3600 ( .A1(n3717), .A2(n3716), .B1(n3715), .B2(n3714), .ZN(n3912)
         );
  OAI22_X1 U3601 ( .A1(n3721), .A2(n3720), .B1(n59), .B2(n3718), .ZN(n3911) );
  FA_X1 U3602 ( .A(n3724), .B(n3723), .CI(n3722), .CO(n3728), .S(n3908) );
  FA_X1 U3603 ( .A(n3727), .B(n3726), .CI(n3725), .CO(n3453), .S(n3854) );
  FA_X1 U3604 ( .A(n3730), .B(n3729), .CI(n3728), .CO(n3731), .S(n3853) );
  FA_X1 U3605 ( .A(n3733), .B(n3732), .CI(n3731), .CO(n3599), .S(n3862) );
  FA_X1 U3606 ( .A(n3736), .B(n3735), .CI(n3734), .CO(n3871), .S(n3861) );
  MUX2_X1 U3607 ( .A(n3738), .B(n3737), .S(n6141), .Z(n3875) );
  FA_X1 U3608 ( .A(n3741), .B(n3740), .CI(n3739), .CO(n3746), .S(n3874) );
  FA_X1 U3609 ( .A(n3744), .B(n3743), .CI(n3742), .CO(n3750), .S(n3800) );
  FA_X1 U3610 ( .A(n3747), .B(n3746), .CI(n3745), .CO(n3775), .S(n3799) );
  NOR2_X1 U3611 ( .A1(n4054), .A2(n4053), .ZN(n5492) );
  INV_X1 U3612 ( .A(n5492), .ZN(n5468) );
  FA_X1 U3613 ( .A(n3750), .B(n3749), .CI(n3748), .CO(n3798), .S(n3773) );
  FA_X1 U3614 ( .A(n3753), .B(n3752), .CI(n3751), .CO(n3382), .S(n3758) );
  FA_X1 U3615 ( .A(n3756), .B(n3755), .CI(n3754), .CO(n3381), .S(n3757) );
  MUX2_X1 U3616 ( .A(n3758), .B(n3757), .S(n6145), .Z(n3797) );
  FA_X1 U3617 ( .A(n3761), .B(n3760), .CI(n3759), .CO(n3791), .S(n3781) );
  FA_X1 U3618 ( .A(n3764), .B(n3763), .CI(n3762), .CO(n3780), .S(n3748) );
  FA_X1 U3619 ( .A(n3767), .B(n3766), .CI(n3765), .CO(n3772), .S(n3632) );
  FA_X1 U3620 ( .A(n3770), .B(n3769), .CI(n3768), .CO(n3771), .S(n3631) );
  MUX2_X1 U3621 ( .A(n3772), .B(n3771), .S(n6144), .Z(n3779) );
  FA_X1 U3622 ( .A(n3775), .B(n3774), .CI(n3773), .CO(n4055), .S(n4054) );
  OR2_X1 U3623 ( .A1(n4056), .A2(n4055), .ZN(n5495) );
  NAND2_X1 U3624 ( .A1(n5468), .A2(n5495), .ZN(n5151) );
  FA_X1 U3625 ( .A(n3778), .B(n3777), .CI(n3776), .CO(n4068), .S(n4062) );
  FA_X1 U3626 ( .A(n3781), .B(n3780), .CI(n3779), .CO(n3795), .S(n3796) );
  FA_X1 U3627 ( .A(n3784), .B(n3783), .CI(n3782), .CO(n3277), .S(n3789) );
  FA_X1 U3628 ( .A(n3787), .B(n3786), .CI(n3785), .CO(n3276), .S(n3788) );
  MUX2_X1 U3629 ( .A(n3789), .B(n3788), .S(n6145), .Z(n3794) );
  FA_X1 U3630 ( .A(n3792), .B(n3791), .CI(n3790), .CO(n3777), .S(n3793) );
  OR2_X1 U3631 ( .A1(n4062), .A2(n4061), .ZN(n5154) );
  FA_X1 U3632 ( .A(n3795), .B(n3794), .CI(n3793), .CO(n4061), .S(n4060) );
  FA_X1 U3633 ( .A(n3798), .B(n3797), .CI(n3796), .CO(n4059), .S(n4056) );
  OR2_X1 U3634 ( .A1(n4060), .A2(n4059), .ZN(n5526) );
  NAND2_X1 U3635 ( .A1(n5154), .A2(n5526), .ZN(n4065) );
  NOR2_X1 U3636 ( .A1(n5151), .A2(n4065), .ZN(n4067) );
  FA_X1 U3637 ( .A(n3801), .B(n3800), .CI(n3799), .CO(n4053), .S(n4049) );
  FA_X1 U3638 ( .A(n3804), .B(n3803), .CI(n3802), .CO(n3688), .S(n3896) );
  FA_X1 U3639 ( .A(n3807), .B(n3806), .CI(n3805), .CO(n3803), .S(n3888) );
  FA_X1 U3640 ( .A(n3810), .B(n3809), .CI(n3808), .CO(n3887), .S(n3975) );
  FA_X1 U3641 ( .A(n3813), .B(n3812), .CI(n3811), .CO(n3683), .S(n3886) );
  FA_X1 U3642 ( .A(n3816), .B(n3815), .CI(n3814), .CO(n3823), .S(n3894) );
  INV_X1 U3643 ( .A(op_b_i[8]), .ZN(n3817) );
  NOR2_X1 U3644 ( .A1(n6119), .A2(n3817), .ZN(n3818) );
  MUX2_X1 U3645 ( .A(n3819), .B(n3818), .S(n29), .Z(n4028) );
  INV_X1 U3646 ( .A(op_c_i[8]), .ZN(n3820) );
  OAI22_X1 U3647 ( .A1(n6146), .A2(n3821), .B1(n2525), .B2(n3820), .ZN(n4027)
         );
  FA_X1 U3648 ( .A(n3824), .B(n3823), .CI(n3822), .CO(n3690), .S(n3825) );
  AND2_X1 U3649 ( .A1(n3825), .A2(n6144), .ZN(n4026) );
  FA_X1 U3650 ( .A(n3828), .B(n3827), .CI(n3826), .CO(n3704), .S(n3927) );
  OR2_X1 U3651 ( .A1(n6116), .A2(n3889), .ZN(n3829) );
  OAI22_X1 U3652 ( .A1(n3829), .A2(n5922), .B1(n3128), .B2(n3889), .ZN(n3907)
         );
  XNOR2_X1 U3653 ( .A(n19), .B(n4337), .ZN(n3898) );
  OAI22_X1 U3654 ( .A1(n3830), .A2(n5635), .B1(n3898), .B2(n3241), .ZN(n3906)
         );
  XNOR2_X1 U3655 ( .A(n6116), .B(n5919), .ZN(n3832) );
  OAI22_X1 U3656 ( .A1(n3832), .A2(n3128), .B1(n3831), .B2(n5922), .ZN(n3905)
         );
  FA_X1 U3657 ( .A(n3835), .B(n3834), .CI(n3833), .CO(n3859), .S(n3925) );
  FA_X1 U3658 ( .A(n3838), .B(n3837), .CI(n3836), .CO(n3736), .S(n3930) );
  FA_X1 U3659 ( .A(n3841), .B(n3840), .CI(n3839), .CO(n3951), .S(n3946) );
  HA_X1 U3660 ( .A(n3843), .B(n3842), .CO(n3852), .S(n3950) );
  FA_X1 U3661 ( .A(n3846), .B(n3845), .CI(n3844), .CO(n3949), .S(n3948) );
  FA_X1 U3662 ( .A(n3849), .B(n3848), .CI(n3847), .CO(n3729), .S(n3921) );
  FA_X1 U3663 ( .A(n3852), .B(n3851), .CI(n3850), .CO(n3836), .S(n3920) );
  FA_X1 U3664 ( .A(n3855), .B(n3854), .CI(n3853), .CO(n3863), .S(n3928) );
  MUX2_X1 U3665 ( .A(n3857), .B(n3856), .S(n6145), .Z(n3937) );
  FA_X1 U3666 ( .A(n3860), .B(n3859), .CI(n3858), .CO(n3738), .S(n3865) );
  FA_X1 U3667 ( .A(n3863), .B(n3862), .CI(n3861), .CO(n3737), .S(n3864) );
  MUX2_X1 U3668 ( .A(n3865), .B(n3864), .S(n6144), .Z(n3936) );
  FA_X1 U3669 ( .A(n3868), .B(n3867), .CI(n3866), .CO(n3484), .S(n3873) );
  FA_X1 U3670 ( .A(n3871), .B(n3870), .CI(n3869), .CO(n3483), .S(n3872) );
  MUX2_X1 U3671 ( .A(n3873), .B(n3872), .S(n6144), .Z(n3878) );
  FA_X1 U3672 ( .A(n3876), .B(n3875), .CI(n3874), .CO(n3801), .S(n3877) );
  OR2_X1 U3673 ( .A1(n4049), .A2(n4048), .ZN(n5436) );
  FA_X1 U3674 ( .A(n3879), .B(n3878), .CI(n3877), .CO(n4048), .S(n4047) );
  FA_X1 U3675 ( .A(n3882), .B(n3881), .CI(n3880), .CO(n3984), .S(n3974) );
  FA_X1 U3676 ( .A(n3885), .B(n3884), .CI(n3883), .CO(n3816), .S(n3983) );
  FA_X1 U3677 ( .A(n3888), .B(n3887), .CI(n3886), .CO(n3895), .S(n3982) );
  INV_X1 U3678 ( .A(op_b_i[7]), .ZN(n3889) );
  NOR2_X1 U3679 ( .A1(n6118), .A2(n3889), .ZN(n3890) );
  MUX2_X1 U3680 ( .A(n3891), .B(n3890), .S(n29), .Z(n3997) );
  INV_X1 U3681 ( .A(op_c_i[7]), .ZN(n3892) );
  OAI22_X1 U3682 ( .A1(n6146), .A2(n3893), .B1(n2525), .B2(n3892), .ZN(n3996)
         );
  FA_X1 U3683 ( .A(n3896), .B(n3895), .CI(n3894), .CO(n3819), .S(n3897) );
  AND2_X1 U3684 ( .A1(n3897), .A2(n6145), .ZN(n3995) );
  OAI22_X1 U3685 ( .A1(n3899), .A2(n3241), .B1(n3898), .B2(n5635), .ZN(n3945)
         );
  AND2_X1 U3686 ( .A1(n6116), .A2(n3900), .ZN(n3944) );
  OAI22_X1 U3687 ( .A1(n3902), .A2(n2585), .B1(n3901), .B2(n10), .ZN(n3943) );
  HA_X1 U3688 ( .A(n3904), .B(n3903), .CO(n3833), .S(n4010) );
  FA_X1 U3689 ( .A(n3907), .B(n3906), .CI(n3905), .CO(n3926), .S(n4009) );
  FA_X1 U3690 ( .A(n3910), .B(n3909), .CI(n3908), .CO(n3855), .S(n4014) );
  FA_X1 U3691 ( .A(n3913), .B(n3912), .CI(n3911), .CO(n3909), .S(n3954) );
  FA_X1 U3692 ( .A(n3916), .B(n3915), .CI(n3914), .CO(n3953), .S(n3967) );
  FA_X1 U3693 ( .A(n3919), .B(n3918), .CI(n3917), .CO(n3850), .S(n3952) );
  FA_X1 U3694 ( .A(n3922), .B(n3921), .CI(n3920), .CO(n3929), .S(n4012) );
  MUX2_X1 U3695 ( .A(n3924), .B(n3923), .S(n6145), .Z(n4030) );
  FA_X1 U3696 ( .A(n3927), .B(n3926), .CI(n3925), .CO(n3857), .S(n3932) );
  FA_X1 U3697 ( .A(n3930), .B(n3929), .CI(n3928), .CO(n3856), .S(n3931) );
  MUX2_X1 U3698 ( .A(n3932), .B(n3931), .S(n6145), .Z(n4029) );
  FA_X1 U3699 ( .A(n3935), .B(n3934), .CI(n3933), .CO(n3876), .S(n4038) );
  FA_X1 U3700 ( .A(n3938), .B(n3937), .CI(n3936), .CO(n3879), .S(n4037) );
  OR2_X1 U3701 ( .A1(n4047), .A2(n4046), .ZN(n5433) );
  NAND2_X1 U3702 ( .A1(n5436), .A2(n5433), .ZN(n4052) );
  HA_X1 U3703 ( .A(n3940), .B(n3939), .CO(n4000), .S(n3963) );
  OAI22_X1 U3704 ( .A1(n3942), .A2(n2867), .B1(n3941), .B2(n5809), .ZN(n3999)
         );
  FA_X1 U3705 ( .A(n3945), .B(n3944), .CI(n3943), .CO(n4011), .S(n3998) );
  FA_X1 U3706 ( .A(n3948), .B(n3947), .CI(n3946), .CO(n4003), .S(n3966) );
  FA_X1 U3707 ( .A(n3951), .B(n3950), .CI(n3949), .CO(n3922), .S(n4002) );
  FA_X1 U3708 ( .A(n3954), .B(n3953), .CI(n3952), .CO(n4013), .S(n4001) );
  MUX2_X1 U3709 ( .A(n3956), .B(n3955), .S(n6145), .Z(n4019) );
  FA_X1 U3710 ( .A(n3959), .B(n3958), .CI(n3957), .CO(n4018), .S(n2594) );
  FA_X1 U3711 ( .A(n3962), .B(n3961), .CI(n3960), .CO(n4017), .S(n2595) );
  FA_X1 U3712 ( .A(n3965), .B(n3964), .CI(n3963), .CO(n3970), .S(n2424) );
  FA_X1 U3713 ( .A(n3968), .B(n3967), .CI(n3966), .CO(n3969), .S(n2423) );
  MUX2_X1 U3714 ( .A(n3970), .B(n3969), .S(n6143), .Z(n3994) );
  FA_X1 U3715 ( .A(n3973), .B(n3972), .CI(n3971), .CO(n3993), .S(n3961) );
  FA_X1 U3716 ( .A(n3976), .B(n3975), .CI(n3974), .CO(n3979), .S(n2558) );
  INV_X1 U3717 ( .A(op_b_i[6]), .ZN(n3977) );
  NOR2_X1 U3718 ( .A1(n6119), .A2(n3977), .ZN(n3978) );
  MUX2_X1 U3719 ( .A(n3979), .B(n3978), .S(n29), .Z(n4008) );
  INV_X1 U3720 ( .A(op_c_i[6]), .ZN(n3980) );
  OAI22_X1 U3721 ( .A1(n6112), .A2(n3981), .B1(n2525), .B2(n3980), .ZN(n4007)
         );
  FA_X1 U3722 ( .A(n3984), .B(n3983), .CI(n3982), .CO(n3891), .S(n3985) );
  AND2_X1 U3723 ( .A1(n3985), .A2(n6141), .ZN(n4006) );
  NOR2_X1 U3724 ( .A1(n3991), .A2(n3990), .ZN(n5353) );
  INV_X1 U3725 ( .A(n3986), .ZN(n3987) );
  AOI21_X1 U3726 ( .B1(n3989), .B2(n3988), .A(n3987), .ZN(n5356) );
  NAND2_X1 U3727 ( .A1(n3991), .A2(n3990), .ZN(n5354) );
  OAI21_X1 U3728 ( .B1(n5353), .B2(n5356), .A(n5354), .ZN(n5043) );
  FA_X1 U3729 ( .A(n3994), .B(n3993), .CI(n3992), .CO(n4034), .S(n3990) );
  FA_X1 U3730 ( .A(n3997), .B(n3996), .CI(n3995), .CO(n4031), .S(n4033) );
  FA_X1 U3731 ( .A(n4000), .B(n3999), .CI(n3998), .CO(n4005), .S(n3956) );
  FA_X1 U3732 ( .A(n4003), .B(n4002), .CI(n4001), .CO(n4004), .S(n3955) );
  MUX2_X1 U3733 ( .A(n4005), .B(n4004), .S(n6144), .Z(n4025) );
  FA_X1 U3734 ( .A(n4008), .B(n4007), .CI(n4006), .CO(n4024), .S(n3992) );
  FA_X1 U3735 ( .A(n4011), .B(n4010), .CI(n4009), .CO(n3924), .S(n4016) );
  FA_X1 U3736 ( .A(n4014), .B(n4013), .CI(n4012), .CO(n3923), .S(n4015) );
  MUX2_X1 U3737 ( .A(n4016), .B(n4015), .S(n6144), .Z(n4023) );
  FA_X1 U3738 ( .A(n4019), .B(n4018), .CI(n4017), .CO(n4020), .S(n3991) );
  OR2_X1 U3739 ( .A1(n4021), .A2(n4020), .ZN(n5042) );
  NAND2_X1 U3740 ( .A1(n4021), .A2(n4020), .ZN(n5041) );
  INV_X1 U3741 ( .A(n5041), .ZN(n4022) );
  AOI21_X1 U3742 ( .B1(n5043), .B2(n5042), .A(n4022), .ZN(n5390) );
  FA_X1 U3743 ( .A(n4025), .B(n4024), .CI(n4023), .CO(n4042), .S(n4032) );
  FA_X1 U3744 ( .A(n4028), .B(n4027), .CI(n4026), .CO(n3938), .S(n4041) );
  FA_X1 U3745 ( .A(n4031), .B(n4030), .CI(n4029), .CO(n4039), .S(n4040) );
  FA_X1 U3746 ( .A(n4034), .B(n4033), .CI(n4032), .CO(n4035), .S(n4021) );
  NOR2_X1 U3747 ( .A1(n4036), .A2(n4035), .ZN(n5387) );
  NAND2_X1 U3748 ( .A1(n4036), .A2(n4035), .ZN(n5388) );
  OAI21_X1 U3749 ( .B1(n5390), .B2(n5387), .A(n5388), .ZN(n5408) );
  FA_X1 U3750 ( .A(n4039), .B(n4038), .CI(n4037), .CO(n4046), .S(n4044) );
  FA_X1 U3751 ( .A(n4042), .B(n4041), .CI(n4040), .CO(n4043), .S(n4036) );
  OR2_X1 U3752 ( .A1(n4044), .A2(n4043), .ZN(n5407) );
  NAND2_X1 U3753 ( .A1(n4044), .A2(n4043), .ZN(n5406) );
  INV_X1 U3754 ( .A(n5406), .ZN(n4045) );
  AOI21_X1 U3755 ( .B1(n5408), .B2(n5407), .A(n4045), .ZN(n4983) );
  NAND2_X1 U3756 ( .A1(n4047), .A2(n4046), .ZN(n4982) );
  INV_X1 U3757 ( .A(n4982), .ZN(n5432) );
  NAND2_X1 U3758 ( .A1(n4049), .A2(n4048), .ZN(n5435) );
  INV_X1 U3759 ( .A(n5435), .ZN(n4050) );
  AOI21_X1 U3760 ( .B1(n5436), .B2(n5432), .A(n4050), .ZN(n4051) );
  OAI21_X1 U3761 ( .B1(n4052), .B2(n4983), .A(n4051), .ZN(n5149) );
  NAND2_X1 U3762 ( .A1(n4054), .A2(n4053), .ZN(n5491) );
  INV_X1 U3763 ( .A(n5491), .ZN(n4058) );
  NAND2_X1 U3764 ( .A1(n4056), .A2(n4055), .ZN(n5494) );
  INV_X1 U3765 ( .A(n5494), .ZN(n4057) );
  AOI21_X1 U3766 ( .B1(n5495), .B2(n4058), .A(n4057), .ZN(n5150) );
  NAND2_X1 U3767 ( .A1(n4060), .A2(n4059), .ZN(n5525) );
  INV_X1 U3768 ( .A(n5525), .ZN(n5152) );
  NAND2_X1 U3769 ( .A1(n4062), .A2(n4061), .ZN(n5153) );
  INV_X1 U3770 ( .A(n5153), .ZN(n4063) );
  AOI21_X1 U3771 ( .B1(n5154), .B2(n5152), .A(n4063), .ZN(n4064) );
  OAI21_X1 U3772 ( .B1(n4065), .B2(n5150), .A(n4064), .ZN(n4066) );
  AOI21_X1 U3773 ( .B1(n4067), .B2(n5149), .A(n4066), .ZN(n4898) );
  NAND2_X1 U3774 ( .A1(n4069), .A2(n4068), .ZN(n5559) );
  NAND2_X1 U3775 ( .A1(n4071), .A2(n4070), .ZN(n4902) );
  OAI21_X1 U3776 ( .B1(n4901), .B2(n5559), .A(n4902), .ZN(n4927) );
  NAND2_X1 U3777 ( .A1(n4073), .A2(n4072), .ZN(n5178) );
  NAND2_X1 U3778 ( .A1(n4075), .A2(n4074), .ZN(n4930) );
  OAI21_X1 U3779 ( .B1(n4929), .B2(n5178), .A(n4930), .ZN(n4076) );
  AOI21_X1 U3780 ( .B1(n4077), .B2(n4927), .A(n4076), .ZN(n4078) );
  OAI21_X1 U3781 ( .B1(n4079), .B2(n4898), .A(n4078), .ZN(n4885) );
  INV_X1 U3782 ( .A(op_b_i[22]), .ZN(n4080) );
  NOR2_X1 U3783 ( .A1(n6119), .A2(n4080), .ZN(n4081) );
  OR2_X1 U3784 ( .A1(n4081), .A2(n6145), .ZN(n4228) );
  INV_X1 U3785 ( .A(op_c_i[22]), .ZN(n4082) );
  OAI22_X1 U3786 ( .A1(n6146), .A2(n4083), .B1(n2525), .B2(n4082), .ZN(n4227)
         );
  INV_X1 U3787 ( .A(op_b_i[21]), .ZN(n4084) );
  NOR2_X1 U3788 ( .A1(n6119), .A2(n4084), .ZN(n4085) );
  OR2_X1 U3789 ( .A1(n4085), .A2(n6145), .ZN(n4240) );
  INV_X1 U3790 ( .A(op_c_i[21]), .ZN(n4086) );
  OAI22_X1 U3791 ( .A1(n6146), .A2(n4087), .B1(n2525), .B2(n4086), .ZN(n4239)
         );
  XNOR2_X1 U3792 ( .A(n55), .B(op_b_i[17]), .ZN(n4109) );
  OAI22_X1 U3793 ( .A1(n4088), .A2(n5915), .B1(n4109), .B2(n5917), .ZN(n4134)
         );
  XNOR2_X1 U3794 ( .A(n52), .B(n5941), .ZN(n4108) );
  OAI22_X1 U3795 ( .A1(n4089), .A2(n5943), .B1(n4108), .B2(n26), .ZN(n4133) );
  XNOR2_X1 U3796 ( .A(n19), .B(n4123), .ZN(n4124) );
  OAI22_X1 U3797 ( .A1(n4090), .A2(n5925), .B1(n4124), .B2(n5927), .ZN(n4132)
         );
  XNOR2_X1 U3798 ( .A(n5848), .B(op_b_i[19]), .ZN(n4119) );
  OAI22_X1 U3799 ( .A1(n4091), .A2(n6032), .B1(n4119), .B2(n6034), .ZN(n4112)
         );
  XNOR2_X1 U3800 ( .A(op_b_i[20]), .B(op_b_i[19]), .ZN(n5999) );
  AND2_X1 U3801 ( .A1(n6116), .A2(n67), .ZN(n4111) );
  XNOR2_X1 U3802 ( .A(n5853), .B(n27), .ZN(n4125) );
  OAI22_X1 U3803 ( .A1(n4092), .A2(n5822), .B1(n4125), .B2(n4546), .ZN(n4110)
         );
  XNOR2_X1 U3804 ( .A(n20), .B(op_b_i[13]), .ZN(n4120) );
  OAI22_X1 U3805 ( .A1(n4093), .A2(n5934), .B1(n4120), .B2(n72), .ZN(n4131) );
  XNOR2_X1 U3806 ( .A(n5844), .B(n4383), .ZN(n4127) );
  OAI22_X1 U3807 ( .A1(n4094), .A2(n3128), .B1(n4127), .B2(n5922), .ZN(n4130)
         );
  XNOR2_X1 U3808 ( .A(n6119), .B(op_a_i[20]), .ZN(n5867) );
  XNOR2_X1 U3809 ( .A(n5867), .B(n4337), .ZN(n4128) );
  OAI22_X1 U3810 ( .A1(n4095), .A2(n3241), .B1(n4128), .B2(n5635), .ZN(n4129)
         );
  FA_X1 U3811 ( .A(n4098), .B(n4097), .CI(n4096), .CO(n4115), .S(n4150) );
  FA_X1 U3812 ( .A(n4101), .B(n4100), .CI(n4099), .CO(n4114), .S(n4148) );
  FA_X1 U3813 ( .A(n4104), .B(n4103), .CI(n4102), .CO(n4113), .S(n4106) );
  FA_X1 U3814 ( .A(n4107), .B(n4106), .CI(n4105), .CO(n4250), .S(n4269) );
  XNOR2_X1 U3815 ( .A(n51), .B(n5941), .ZN(n4168) );
  OAI22_X1 U3816 ( .A1(n4168), .A2(n26), .B1(n4108), .B2(n5943), .ZN(n4192) );
  XNOR2_X1 U3817 ( .A(n22), .B(op_b_i[17]), .ZN(n4155) );
  OAI22_X1 U3818 ( .A1(n4155), .A2(n5917), .B1(n4109), .B2(n5915), .ZN(n4191)
         );
  XNOR2_X1 U3819 ( .A(n5933), .B(n6015), .ZN(n4153) );
  XNOR2_X1 U3820 ( .A(n5824), .B(n6015), .ZN(n4138) );
  OAI22_X1 U3821 ( .A1(n4153), .A2(n10), .B1(n4138), .B2(n2585), .ZN(n4159) );
  FA_X1 U3822 ( .A(n4112), .B(n4111), .CI(n4110), .CO(n4158), .S(n4117) );
  FA_X1 U3823 ( .A(n4115), .B(n4114), .CI(n4113), .CO(n4171), .S(n4251) );
  FA_X1 U3824 ( .A(n4118), .B(n4117), .CI(n4116), .CO(n4170), .S(n4252) );
  XNOR2_X1 U3825 ( .A(n5976), .B(op_b_i[19]), .ZN(n4167) );
  OAI22_X1 U3826 ( .A1(n4167), .A2(n6034), .B1(n4119), .B2(n6032), .ZN(n4190)
         );
  XNOR2_X1 U3827 ( .A(n21), .B(op_b_i[13]), .ZN(n4156) );
  OAI22_X1 U3828 ( .A1(n4156), .A2(n5936), .B1(n4120), .B2(n5934), .ZN(n4189)
         );
  XNOR2_X1 U3829 ( .A(n6116), .B(op_b_i[21]), .ZN(n4122) );
  XOR2_X1 U3830 ( .A(op_b_i[20]), .B(op_b_i[21]), .Z(n4121) );
  NAND2_X1 U3831 ( .A1(n4121), .A2(n5999), .ZN(n5997) );
  XNOR2_X1 U3832 ( .A(n6002), .B(op_b_i[21]), .ZN(n4161) );
  OAI22_X1 U3833 ( .A1(n4122), .A2(n5997), .B1(n4161), .B2(n68), .ZN(n4188) );
  XNOR2_X1 U3834 ( .A(n54), .B(n4123), .ZN(n4169) );
  OAI22_X1 U3835 ( .A1(n4169), .A2(n5927), .B1(n4124), .B2(n5925), .ZN(n4195)
         );
  XNOR2_X1 U3836 ( .A(n6031), .B(n27), .ZN(n4163) );
  OAI22_X1 U3837 ( .A1(n4163), .A2(n4546), .B1(n4125), .B2(n5822), .ZN(n4194)
         );
  OR2_X1 U3838 ( .A1(n6116), .A2(n4084), .ZN(n4126) );
  OAI22_X1 U3839 ( .A1(n4126), .A2(n68), .B1(n5997), .B2(n4084), .ZN(n4193) );
  XNOR2_X1 U3840 ( .A(n5914), .B(n4383), .ZN(n4152) );
  OAI22_X1 U3841 ( .A1(n4152), .A2(n5922), .B1(n4127), .B2(n3128), .ZN(n4166)
         );
  XNOR2_X1 U3842 ( .A(n6119), .B(op_a_i[21]), .ZN(n5942) );
  XNOR2_X1 U3843 ( .A(n5942), .B(n4337), .ZN(n4157) );
  OAI22_X1 U3844 ( .A1(n4157), .A2(n5635), .B1(n4128), .B2(n3241), .ZN(n4165)
         );
  XNOR2_X1 U3845 ( .A(n5924), .B(n25), .ZN(n4154) );
  XNOR2_X1 U3846 ( .A(n5819), .B(n25), .ZN(n4135) );
  OAI22_X1 U3847 ( .A1(n4154), .A2(n5809), .B1(n4135), .B2(n2867), .ZN(n4164)
         );
  FA_X1 U3848 ( .A(n4131), .B(n4130), .CI(n4129), .CO(n4218), .S(n4116) );
  FA_X1 U3849 ( .A(n4134), .B(n4133), .CI(n4132), .CO(n4217), .S(n4118) );
  OAI22_X1 U3850 ( .A1(n4136), .A2(n2867), .B1(n4135), .B2(n5809), .ZN(n4147)
         );
  OAI22_X1 U3851 ( .A1(n4139), .A2(n2585), .B1(n4138), .B2(n10), .ZN(n4146) );
  HA_X1 U3852 ( .A(n4141), .B(n4140), .CO(n4145), .S(n4143) );
  FA_X1 U3853 ( .A(n4144), .B(n4143), .CI(n4142), .CO(n4249), .S(n4245) );
  FA_X1 U3854 ( .A(n4147), .B(n4146), .CI(n4145), .CO(n4216), .S(n4248) );
  FA_X1 U3855 ( .A(n4150), .B(n4149), .CI(n4148), .CO(n4247), .S(n4244) );
  OR2_X1 U3856 ( .A1(n4151), .A2(n6145), .ZN(n4258) );
  XNOR2_X1 U3857 ( .A(n5819), .B(n4383), .ZN(n4198) );
  OAI22_X1 U3858 ( .A1(n4152), .A2(n3128), .B1(n4198), .B2(n5922), .ZN(n4209)
         );
  XNOR2_X1 U3859 ( .A(n5867), .B(n4342), .ZN(n4200) );
  OAI22_X1 U3860 ( .A1(n4153), .A2(n2585), .B1(n4200), .B2(n10), .ZN(n4208) );
  XNOR2_X1 U3861 ( .A(n5824), .B(n25), .ZN(n4199) );
  OAI22_X1 U3862 ( .A1(n4154), .A2(n2867), .B1(n4199), .B2(n5809), .ZN(n4207)
         );
  XNOR2_X1 U3863 ( .A(n19), .B(op_b_i[17]), .ZN(n4210) );
  OAI22_X1 U3864 ( .A1(n4155), .A2(n5915), .B1(n4210), .B2(n5917), .ZN(n4181)
         );
  XNOR2_X1 U3865 ( .A(n52), .B(op_b_i[13]), .ZN(n4204) );
  OAI22_X1 U3866 ( .A1(n4156), .A2(n5934), .B1(n4204), .B2(n5936), .ZN(n4180)
         );
  XNOR2_X1 U3867 ( .A(n6119), .B(op_a_i[22]), .ZN(n5821) );
  XNOR2_X1 U3868 ( .A(n5821), .B(n4337), .ZN(n4197) );
  OAI22_X1 U3869 ( .A1(n4157), .A2(n3241), .B1(n4197), .B2(n5635), .ZN(n4179)
         );
  FA_X1 U3870 ( .A(n4160), .B(n4159), .CI(n4158), .CO(n4185), .S(n4172) );
  XNOR2_X1 U3871 ( .A(n5848), .B(op_b_i[21]), .ZN(n4203) );
  OAI22_X1 U3872 ( .A1(n4161), .A2(n5997), .B1(n4203), .B2(n68), .ZN(n4178) );
  INV_X1 U3873 ( .A(n5983), .ZN(n4162) );
  AND2_X1 U3874 ( .A1(n6116), .A2(n4162), .ZN(n4177) );
  XNOR2_X1 U3875 ( .A(n5844), .B(n27), .ZN(n4196) );
  OAI22_X1 U3876 ( .A1(n4163), .A2(n5822), .B1(n4196), .B2(n4546), .ZN(n4176)
         );
  FA_X1 U3877 ( .A(n4166), .B(n4165), .CI(n4164), .CO(n4183), .S(n4219) );
  XNOR2_X1 U3878 ( .A(n55), .B(op_b_i[19]), .ZN(n4202) );
  OAI22_X1 U3879 ( .A1(n4167), .A2(n6032), .B1(n4202), .B2(n6034), .ZN(n4175)
         );
  XNOR2_X1 U3880 ( .A(n5853), .B(n5941), .ZN(n4201) );
  OAI22_X1 U3881 ( .A1(n4168), .A2(n5943), .B1(n4201), .B2(n26), .ZN(n4174) );
  XNOR2_X1 U3882 ( .A(n20), .B(n4123), .ZN(n4211) );
  OAI22_X1 U3883 ( .A1(n4169), .A2(n5925), .B1(n4211), .B2(n5927), .ZN(n4173)
         );
  FA_X1 U3884 ( .A(n4172), .B(n4171), .CI(n4170), .CO(n4235), .S(n4273) );
  FA_X1 U3885 ( .A(n4175), .B(n4174), .CI(n4173), .CO(n4335), .S(n4182) );
  FA_X1 U3886 ( .A(n4178), .B(n4177), .CI(n4176), .CO(n4334), .S(n4184) );
  FA_X1 U3887 ( .A(n4181), .B(n4180), .CI(n4179), .CO(n4333), .S(n4186) );
  FA_X1 U3888 ( .A(n4184), .B(n4183), .CI(n4182), .CO(n4322), .S(n4236) );
  FA_X1 U3889 ( .A(n4187), .B(n4186), .CI(n4185), .CO(n4321), .S(n4237) );
  FA_X1 U3890 ( .A(n4190), .B(n4189), .CI(n4188), .CO(n4215), .S(n4221) );
  HA_X1 U3891 ( .A(n4192), .B(n4191), .CO(n4214), .S(n4160) );
  FA_X1 U3892 ( .A(n4195), .B(n4194), .CI(n4193), .CO(n4213), .S(n4220) );
  XNOR2_X1 U3893 ( .A(n5914), .B(n27), .ZN(n4336) );
  OAI22_X1 U3894 ( .A1(n4336), .A2(n4546), .B1(n4196), .B2(n5822), .ZN(n4364)
         );
  XNOR2_X1 U3895 ( .A(n6119), .B(op_a_i[23]), .ZN(n5938) );
  XNOR2_X1 U3896 ( .A(n5938), .B(n4337), .ZN(n4338) );
  OAI22_X1 U3897 ( .A1(n4338), .A2(n5635), .B1(n4197), .B2(n3241), .ZN(n4363)
         );
  XNOR2_X1 U3898 ( .A(n5924), .B(n4383), .ZN(n4339) );
  OAI22_X1 U3899 ( .A1(n4339), .A2(n5922), .B1(n4198), .B2(n3128), .ZN(n4362)
         );
  XNOR2_X1 U3900 ( .A(n5933), .B(n25), .ZN(n4332) );
  OAI22_X1 U3901 ( .A1(n4332), .A2(n5809), .B1(n4199), .B2(n2867), .ZN(n4326)
         );
  XNOR2_X1 U3902 ( .A(n5942), .B(n4342), .ZN(n4343) );
  OAI22_X1 U3903 ( .A1(n4343), .A2(n10), .B1(n4200), .B2(n2585), .ZN(n4325) );
  XNOR2_X1 U3904 ( .A(n66), .B(n5941), .ZN(n4371) );
  OAI22_X1 U3905 ( .A1(n4371), .A2(n26), .B1(n4201), .B2(n5943), .ZN(n4341) );
  XNOR2_X1 U3906 ( .A(n22), .B(op_b_i[19]), .ZN(n4327) );
  OAI22_X1 U3907 ( .A1(n4327), .A2(n6034), .B1(n4202), .B2(n6032), .ZN(n4340)
         );
  XNOR2_X1 U3908 ( .A(n56), .B(op_b_i[21]), .ZN(n4329) );
  OAI22_X1 U3909 ( .A1(n4329), .A2(n68), .B1(n4203), .B2(n5997), .ZN(n4346) );
  XNOR2_X1 U3910 ( .A(n51), .B(op_b_i[13]), .ZN(n4328) );
  OAI22_X1 U3911 ( .A1(n4328), .A2(n5936), .B1(n4204), .B2(n5934), .ZN(n4345)
         );
  XNOR2_X1 U3912 ( .A(n6116), .B(op_b_i[23]), .ZN(n4206) );
  XOR2_X1 U3913 ( .A(op_b_i[22]), .B(op_b_i[23]), .Z(n4205) );
  NAND2_X1 U3914 ( .A1(n4205), .A2(n5983), .ZN(n5981) );
  XNOR2_X1 U3915 ( .A(n6002), .B(op_b_i[23]), .ZN(n4369) );
  OAI22_X1 U3916 ( .A1(n4206), .A2(n5981), .B1(n4369), .B2(n5983), .ZN(n4344)
         );
  FA_X1 U3917 ( .A(n4209), .B(n4208), .CI(n4207), .CO(n4398), .S(n4187) );
  XNOR2_X1 U3918 ( .A(n5992), .B(op_b_i[17]), .ZN(n4330) );
  OAI22_X1 U3919 ( .A1(n4330), .A2(n5917), .B1(n4210), .B2(n5915), .ZN(n4367)
         );
  XNOR2_X1 U3920 ( .A(n21), .B(n4123), .ZN(n4331) );
  OAI22_X1 U3921 ( .A1(n4331), .A2(n5927), .B1(n4211), .B2(n5925), .ZN(n4366)
         );
  OR2_X1 U3922 ( .A1(n6116), .A2(n4223), .ZN(n4212) );
  OAI22_X1 U3923 ( .A1(n4212), .A2(n5983), .B1(n5981), .B2(n4223), .ZN(n4365)
         );
  FA_X1 U3924 ( .A(n4215), .B(n4214), .CI(n4213), .CO(n4402), .S(n4234) );
  FA_X1 U3925 ( .A(n4218), .B(n4217), .CI(n4216), .CO(n4233), .S(n4230) );
  FA_X1 U3926 ( .A(n4221), .B(n4220), .CI(n4219), .CO(n4232), .S(n4231) );
  AND2_X1 U3927 ( .A1(n4222), .A2(n29), .ZN(n4432) );
  INV_X1 U3928 ( .A(op_b_i[23]), .ZN(n4223) );
  NOR2_X1 U3929 ( .A1(n6119), .A2(n4223), .ZN(n4224) );
  OR2_X1 U3930 ( .A1(n4224), .A2(n6143), .ZN(n4316) );
  INV_X1 U3931 ( .A(op_c_i[23]), .ZN(n4225) );
  OAI22_X1 U3932 ( .A1(n6146), .A2(n4226), .B1(n2525), .B2(n4225), .ZN(n4315)
         );
  HA_X1 U3933 ( .A(n4228), .B(n4227), .CO(n4419), .S(n4260) );
  FA_X1 U3934 ( .A(n4231), .B(n4230), .CI(n4229), .CO(n4256), .S(n4272) );
  FA_X1 U3935 ( .A(n4234), .B(n4233), .CI(n4232), .CO(n4408), .S(n4255) );
  FA_X1 U3936 ( .A(n4237), .B(n4236), .CI(n4235), .CO(n4319), .S(n4254) );
  OR2_X1 U3937 ( .A1(n4238), .A2(n6145), .ZN(n4418) );
  HA_X1 U3938 ( .A(n4240), .B(n4239), .CO(n4259), .S(n4278) );
  INV_X1 U3939 ( .A(op_b_i[20]), .ZN(n4241) );
  NOR2_X1 U3940 ( .A1(n6118), .A2(n4241), .ZN(n4242) );
  OR2_X1 U3941 ( .A1(n4242), .A2(n6144), .ZN(n4265) );
  OAI22_X1 U3942 ( .A1(n6146), .A2(n4243), .B1(n2525), .B2(n699), .ZN(n4264)
         );
  FA_X1 U3943 ( .A(n4246), .B(n4245), .CI(n4244), .CO(n4287), .S(n4268) );
  FA_X1 U3944 ( .A(n4249), .B(n4248), .CI(n4247), .CO(n4229), .S(n4286) );
  FA_X1 U3945 ( .A(n4252), .B(n4251), .CI(n4250), .CO(n4274), .S(n4285) );
  OR2_X1 U3946 ( .A1(n4253), .A2(n6144), .ZN(n4276) );
  FA_X1 U3947 ( .A(n4256), .B(n4255), .CI(n4254), .CO(n4238), .S(n4257) );
  AND2_X1 U3948 ( .A1(n4257), .A2(n29), .ZN(n4262) );
  FA_X1 U3949 ( .A(n4260), .B(n4259), .CI(n4258), .CO(n4433), .S(n4261) );
  OR2_X1 U3950 ( .A1(n4307), .A2(n4306), .ZN(n5598) );
  FA_X1 U3951 ( .A(n4263), .B(n4262), .CI(n4261), .CO(n4306), .S(n4305) );
  HA_X1 U3952 ( .A(n4265), .B(n4264), .CO(n4277), .S(n4291) );
  HA_X1 U3953 ( .A(n4267), .B(n4266), .CO(n4290), .S(n4283) );
  FA_X1 U3954 ( .A(n4270), .B(n4269), .CI(n4268), .CO(n4271), .S(n2990) );
  OR2_X1 U3955 ( .A1(n4271), .A2(n6144), .ZN(n4289) );
  FA_X1 U3956 ( .A(n4274), .B(n4273), .CI(n4272), .CO(n4151), .S(n4275) );
  AND2_X1 U3957 ( .A1(n4275), .A2(n29), .ZN(n4280) );
  FA_X1 U3958 ( .A(n4278), .B(n4277), .CI(n4276), .CO(n4263), .S(n4279) );
  OR2_X1 U3959 ( .A1(n4305), .A2(n4304), .ZN(n5595) );
  NAND2_X1 U3960 ( .A1(n5598), .A2(n5595), .ZN(n4310) );
  FA_X1 U3961 ( .A(n4281), .B(n4280), .CI(n4279), .CO(n4304), .S(n4301) );
  FA_X1 U3962 ( .A(n4284), .B(n4283), .CI(n4282), .CO(n4294), .S(n4295) );
  FA_X1 U3963 ( .A(n4287), .B(n4286), .CI(n4285), .CO(n4253), .S(n4288) );
  AND2_X1 U3964 ( .A1(n4288), .A2(n29), .ZN(n4293) );
  FA_X1 U3965 ( .A(n4291), .B(n4290), .CI(n4289), .CO(n4281), .S(n4292) );
  OR2_X1 U3966 ( .A1(n4301), .A2(n4300), .ZN(n5570) );
  FA_X1 U3967 ( .A(n4294), .B(n4293), .CI(n4292), .CO(n4300), .S(n4299) );
  FA_X1 U3968 ( .A(n4297), .B(n4296), .CI(n4295), .CO(n4298), .S(n4075) );
  NOR2_X1 U3969 ( .A1(n4299), .A2(n4298), .ZN(n5568) );
  INV_X1 U3970 ( .A(n5568), .ZN(n4886) );
  NAND2_X1 U3971 ( .A1(n5570), .A2(n4886), .ZN(n5582) );
  NOR2_X1 U3972 ( .A1(n4310), .A2(n5582), .ZN(n4312) );
  NAND2_X1 U3973 ( .A1(n4299), .A2(n4298), .ZN(n5567) );
  INV_X1 U3974 ( .A(n5567), .ZN(n4303) );
  NAND2_X1 U3975 ( .A1(n4301), .A2(n4300), .ZN(n5569) );
  INV_X1 U3976 ( .A(n5569), .ZN(n4302) );
  AOI21_X1 U3977 ( .B1(n5570), .B2(n4303), .A(n4302), .ZN(n5581) );
  NAND2_X1 U3978 ( .A1(n4305), .A2(n4304), .ZN(n5584) );
  INV_X1 U3979 ( .A(n5584), .ZN(n5594) );
  NAND2_X1 U3980 ( .A1(n4307), .A2(n4306), .ZN(n5597) );
  INV_X1 U3981 ( .A(n5597), .ZN(n4308) );
  AOI21_X1 U3982 ( .B1(n5598), .B2(n5594), .A(n4308), .ZN(n4309) );
  OAI21_X1 U3983 ( .B1(n5581), .B2(n4310), .A(n4309), .ZN(n4311) );
  AOI21_X1 U3984 ( .B1(n4885), .B2(n4312), .A(n4311), .ZN(n5718) );
  INV_X1 U3985 ( .A(n5718), .ZN(n5614) );
  INV_X1 U3986 ( .A(op_b_i[24]), .ZN(n4313) );
  NOR2_X1 U3987 ( .A1(n6118), .A2(n4313), .ZN(n4314) );
  OR2_X1 U3988 ( .A1(n4314), .A2(n6144), .ZN(n4407) );
  INV_X1 U3989 ( .A(dot_op_c_i[24]), .ZN(n5617) );
  OAI22_X1 U3990 ( .A1(n6146), .A2(n5617), .B1(n2525), .B2(n825), .ZN(n4406)
         );
  HA_X1 U3991 ( .A(n4316), .B(n4315), .CO(n4426), .S(n4420) );
  FA_X1 U3992 ( .A(n4319), .B(n4318), .CI(n4317), .CO(n4320), .S(n4222) );
  OR2_X1 U3993 ( .A1(n4320), .A2(n6145), .ZN(n4425) );
  FA_X1 U3994 ( .A(n4323), .B(n4322), .CI(n4321), .CO(n4416), .S(n4318) );
  FA_X1 U3995 ( .A(n4326), .B(n4325), .CI(n4324), .CO(n4358), .S(n4400) );
  XNOR2_X1 U3996 ( .A(n19), .B(op_b_i[19]), .ZN(n4388) );
  OAI22_X1 U3997 ( .A1(n4327), .A2(n6032), .B1(n4388), .B2(n6034), .ZN(n4382)
         );
  XNOR2_X1 U3998 ( .A(n6120), .B(op_b_i[13]), .ZN(n4387) );
  OAI22_X1 U3999 ( .A1(n4328), .A2(n5934), .B1(n4387), .B2(n72), .ZN(n4381) );
  XNOR2_X1 U4000 ( .A(n55), .B(op_b_i[21]), .ZN(n4379) );
  OAI22_X1 U4001 ( .A1(n4329), .A2(n5997), .B1(n4379), .B2(n68), .ZN(n4380) );
  XNOR2_X1 U4002 ( .A(n20), .B(op_b_i[17]), .ZN(n4353) );
  OAI22_X1 U4003 ( .A1(n4330), .A2(n5915), .B1(n4353), .B2(n5917), .ZN(n4352)
         );
  XNOR2_X1 U4004 ( .A(n52), .B(n4123), .ZN(n4378) );
  OAI22_X1 U4005 ( .A1(n4331), .A2(n5925), .B1(n4378), .B2(n5927), .ZN(n4351)
         );
  XNOR2_X1 U4006 ( .A(n5867), .B(n25), .ZN(n4386) );
  OAI22_X1 U4007 ( .A1(n4332), .A2(n2867), .B1(n4386), .B2(n5809), .ZN(n4350)
         );
  FA_X1 U4008 ( .A(n4335), .B(n4334), .CI(n4333), .CO(n4361), .S(n4323) );
  XNOR2_X1 U4009 ( .A(n5819), .B(n27), .ZN(n4393) );
  OAI22_X1 U4010 ( .A1(n4336), .A2(n5822), .B1(n4393), .B2(n4546), .ZN(n4349)
         );
  XNOR2_X1 U4011 ( .A(n6119), .B(op_a_i[24]), .ZN(n5814) );
  XNOR2_X1 U4012 ( .A(n5814), .B(n4337), .ZN(n4392) );
  OAI22_X1 U4013 ( .A1(n4338), .A2(n3241), .B1(n4392), .B2(n5635), .ZN(n4348)
         );
  XNOR2_X1 U4014 ( .A(n5824), .B(n4383), .ZN(n4384) );
  OAI22_X1 U4015 ( .A1(n4339), .A2(n3128), .B1(n4384), .B2(n5922), .ZN(n4347)
         );
  HA_X1 U4016 ( .A(n4341), .B(n4340), .CO(n4374), .S(n4324) );
  XNOR2_X1 U4017 ( .A(n5821), .B(n4342), .ZN(n4385) );
  OAI22_X1 U4018 ( .A1(n4343), .A2(n2585), .B1(n4385), .B2(n10), .ZN(n4373) );
  FA_X1 U4019 ( .A(n4346), .B(n4345), .CI(n4344), .CO(n4372), .S(n4399) );
  FA_X1 U4020 ( .A(n4349), .B(n4348), .CI(n4347), .CO(n4464), .S(n4360) );
  FA_X1 U4021 ( .A(n4352), .B(n4351), .CI(n4350), .CO(n4463), .S(n4356) );
  XNOR2_X1 U4022 ( .A(n56), .B(op_b_i[23]), .ZN(n4447) );
  XNOR2_X1 U4023 ( .A(n5848), .B(op_b_i[23]), .ZN(n4368) );
  OAI22_X1 U4024 ( .A1(n4447), .A2(n5983), .B1(n4368), .B2(n5981), .ZN(n4473)
         );
  XNOR2_X1 U4025 ( .A(n21), .B(op_b_i[17]), .ZN(n4446) );
  OAI22_X1 U4026 ( .A1(n4446), .A2(n5917), .B1(n4353), .B2(n5915), .ZN(n4472)
         );
  XNOR2_X1 U4027 ( .A(n6116), .B(op_b_i[25]), .ZN(n4355) );
  XOR2_X1 U4028 ( .A(op_b_i[24]), .B(op_b_i[25]), .Z(n4354) );
  XNOR2_X1 U4029 ( .A(op_b_i[24]), .B(op_b_i[23]), .ZN(n5995) );
  NAND2_X1 U4030 ( .A1(n4354), .A2(n5995), .ZN(n5993) );
  XNOR2_X1 U4031 ( .A(n6002), .B(op_b_i[25]), .ZN(n4440) );
  OAI22_X1 U4032 ( .A1(n4355), .A2(n5993), .B1(n4440), .B2(n5995), .ZN(n4471)
         );
  FA_X1 U4033 ( .A(n4358), .B(n4357), .CI(n4356), .CO(n4481), .S(n4415) );
  FA_X1 U4034 ( .A(n4361), .B(n4360), .CI(n4359), .CO(n4480), .S(n4414) );
  FA_X1 U4035 ( .A(n4364), .B(n4363), .CI(n4362), .CO(n4396), .S(n4401) );
  FA_X1 U4036 ( .A(n4367), .B(n4366), .CI(n4365), .CO(n4395), .S(n4397) );
  OAI22_X1 U4037 ( .A1(n4369), .A2(n5981), .B1(n4368), .B2(n5983), .ZN(n4377)
         );
  INV_X1 U4038 ( .A(n5995), .ZN(n4370) );
  AND2_X1 U4039 ( .A1(n6116), .A2(n4370), .ZN(n4376) );
  XNOR2_X1 U4040 ( .A(n5844), .B(n5941), .ZN(n4391) );
  OAI22_X1 U4041 ( .A1(n4371), .A2(n5943), .B1(n4391), .B2(n26), .ZN(n4375) );
  FA_X1 U4042 ( .A(n4374), .B(n4373), .CI(n4372), .CO(n4478), .S(n4359) );
  FA_X1 U4043 ( .A(n4377), .B(n4376), .CI(n4375), .CO(n4467), .S(n4394) );
  XNOR2_X1 U4044 ( .A(n51), .B(n4123), .ZN(n4448) );
  OAI22_X1 U4045 ( .A1(n4448), .A2(n5927), .B1(n4378), .B2(n5925), .ZN(n4461)
         );
  XNOR2_X1 U4046 ( .A(n22), .B(op_b_i[21]), .ZN(n4442) );
  OAI22_X1 U4047 ( .A1(n4442), .A2(n68), .B1(n4379), .B2(n5997), .ZN(n4460) );
  FA_X1 U4048 ( .A(n4382), .B(n4381), .CI(n4380), .CO(n4465), .S(n4357) );
  XNOR2_X1 U4049 ( .A(n5933), .B(n4383), .ZN(n4458) );
  OAI22_X1 U4050 ( .A1(n4458), .A2(n5922), .B1(n4384), .B2(n3128), .ZN(n4445)
         );
  XNOR2_X1 U4051 ( .A(n5938), .B(n5811), .ZN(n4453) );
  OAI22_X1 U4052 ( .A1(n4453), .A2(n10), .B1(n4385), .B2(n2585), .ZN(n4444) );
  XNOR2_X1 U4053 ( .A(n5942), .B(n5807), .ZN(n4459) );
  OAI22_X1 U4054 ( .A1(n4459), .A2(n6010), .B1(n4386), .B2(n2867), .ZN(n4443)
         );
  XNOR2_X1 U4055 ( .A(n65), .B(op_b_i[13]), .ZN(n4455) );
  OAI22_X1 U4056 ( .A1(n4455), .A2(n72), .B1(n4387), .B2(n5934), .ZN(n4470) );
  XNOR2_X1 U4057 ( .A(n54), .B(op_b_i[19]), .ZN(n4456) );
  OAI22_X1 U4058 ( .A1(n4456), .A2(n6034), .B1(n4388), .B2(n6032), .ZN(n4469)
         );
  INV_X1 U4059 ( .A(op_b_i[25]), .ZN(n4389) );
  OR2_X1 U4060 ( .A1(n6116), .A2(n4389), .ZN(n4390) );
  OAI22_X1 U4061 ( .A1(n4390), .A2(n5995), .B1(n5993), .B2(n4389), .ZN(n4468)
         );
  XNOR2_X1 U4062 ( .A(n5914), .B(n5941), .ZN(n4452) );
  OAI22_X1 U4063 ( .A1(n4452), .A2(n26), .B1(n4391), .B2(n5943), .ZN(n4476) );
  XNOR2_X1 U4064 ( .A(n6118), .B(op_a_i[25]), .ZN(n5920) );
  XNOR2_X1 U4065 ( .A(n5920), .B(n5856), .ZN(n4457) );
  OAI22_X1 U4066 ( .A1(n4457), .A2(n5635), .B1(n4392), .B2(n3241), .ZN(n4475)
         );
  XNOR2_X1 U4067 ( .A(n5924), .B(n27), .ZN(n4454) );
  OAI22_X1 U4068 ( .A1(n4454), .A2(n4546), .B1(n4393), .B2(n5822), .ZN(n4474)
         );
  FA_X1 U4069 ( .A(n4396), .B(n4395), .CI(n4394), .CO(n4479), .S(n4413) );
  FA_X1 U4070 ( .A(n4399), .B(n4398), .CI(n4397), .CO(n4412), .S(n4409) );
  FA_X1 U4071 ( .A(n4402), .B(n4401), .CI(n4400), .CO(n4411), .S(n4410) );
  AND2_X1 U4072 ( .A1(n4403), .A2(n29), .ZN(n4493) );
  NOR2_X1 U4073 ( .A1(n6118), .A2(n4389), .ZN(n4404) );
  OR2_X1 U4074 ( .A1(n4404), .A2(n6145), .ZN(n4487) );
  INV_X1 U4075 ( .A(dot_op_c_i[25]), .ZN(n5204) );
  INV_X1 U4076 ( .A(op_c_i[25]), .ZN(n4405) );
  OAI22_X1 U4077 ( .A1(n6146), .A2(n5204), .B1(n2525), .B2(n4405), .ZN(n4486)
         );
  HA_X1 U4078 ( .A(n4407), .B(n4406), .CO(n4435), .S(n4427) );
  FA_X1 U4079 ( .A(n4410), .B(n4409), .CI(n4408), .CO(n4423), .S(n4317) );
  FA_X1 U4080 ( .A(n4413), .B(n4412), .CI(n4411), .CO(n4437), .S(n4422) );
  FA_X1 U4081 ( .A(n4416), .B(n4415), .CI(n4414), .CO(n4490), .S(n4421) );
  OR2_X1 U4082 ( .A1(n4417), .A2(n6144), .ZN(n4434) );
  FA_X1 U4083 ( .A(n4420), .B(n4419), .CI(n4418), .CO(n4430), .S(n4431) );
  FA_X1 U4084 ( .A(n4423), .B(n4422), .CI(n4421), .CO(n4417), .S(n4424) );
  AND2_X1 U4085 ( .A1(n4424), .A2(n29), .ZN(n4429) );
  FA_X1 U4086 ( .A(n4427), .B(n4426), .CI(n4425), .CO(n4494), .S(n4428) );
  OR2_X1 U4087 ( .A1(n4498), .A2(n4497), .ZN(n5198) );
  FA_X1 U4088 ( .A(n4430), .B(n4429), .CI(n4428), .CO(n4497), .S(n4496) );
  FA_X1 U4089 ( .A(n4433), .B(n4432), .CI(n4431), .CO(n4495), .S(n4307) );
  OR2_X1 U4090 ( .A1(n4496), .A2(n4495), .ZN(n5612) );
  NAND2_X1 U4091 ( .A1(n5198), .A2(n5612), .ZN(n4941) );
  FA_X1 U4092 ( .A(n4436), .B(n4435), .CI(n4434), .CO(n4567), .S(n4492) );
  FA_X1 U4093 ( .A(n4439), .B(n4438), .CI(n4437), .CO(n4563), .S(n4488) );
  XNOR2_X1 U4094 ( .A(n5848), .B(op_b_i[25]), .ZN(n4516) );
  OAI22_X1 U4095 ( .A1(n4440), .A2(n5993), .B1(n4516), .B2(n5995), .ZN(n4533)
         );
  XNOR2_X1 U4096 ( .A(op_b_i[26]), .B(op_b_i[25]), .ZN(n6038) );
  INV_X1 U4097 ( .A(n6038), .ZN(n4441) );
  AND2_X1 U4098 ( .A1(n6116), .A2(n4441), .ZN(n4532) );
  XNOR2_X1 U4099 ( .A(n19), .B(op_b_i[21]), .ZN(n4529) );
  OAI22_X1 U4100 ( .A1(n4442), .A2(n5997), .B1(n4529), .B2(n68), .ZN(n4531) );
  FA_X1 U4101 ( .A(n4445), .B(n4444), .CI(n4443), .CO(n4526), .S(n4451) );
  XNOR2_X1 U4102 ( .A(n52), .B(op_b_i[17]), .ZN(n4528) );
  OAI22_X1 U4103 ( .A1(n4446), .A2(n5915), .B1(n4528), .B2(n5917), .ZN(n4539)
         );
  XNOR2_X1 U4104 ( .A(n55), .B(op_b_i[23]), .ZN(n4508) );
  OAI22_X1 U4105 ( .A1(n4447), .A2(n5981), .B1(n4508), .B2(n5983), .ZN(n4538)
         );
  XNOR2_X1 U4106 ( .A(n6120), .B(n4123), .ZN(n4509) );
  OAI22_X1 U4107 ( .A1(n4448), .A2(n5925), .B1(n4509), .B2(n5927), .ZN(n4537)
         );
  FA_X1 U4108 ( .A(n4451), .B(n4450), .CI(n4449), .CO(n4554), .S(n4438) );
  XNOR2_X1 U4109 ( .A(n5819), .B(n5941), .ZN(n4543) );
  OAI22_X1 U4110 ( .A1(n4452), .A2(n5943), .B1(n4543), .B2(n26), .ZN(n4542) );
  XNOR2_X1 U4111 ( .A(n5814), .B(n5811), .ZN(n4549) );
  OAI22_X1 U4112 ( .A1(n4453), .A2(n2585), .B1(n4549), .B2(n10), .ZN(n4541) );
  XNOR2_X1 U4113 ( .A(n5824), .B(n27), .ZN(n4545) );
  OAI22_X1 U4114 ( .A1(n4454), .A2(n5822), .B1(n4545), .B2(n4546), .ZN(n4540)
         );
  XNOR2_X1 U4115 ( .A(n5844), .B(op_b_i[13]), .ZN(n4547) );
  OAI22_X1 U4116 ( .A1(n4455), .A2(n5934), .B1(n4547), .B2(n72), .ZN(n4536) );
  XNOR2_X1 U4117 ( .A(n20), .B(op_b_i[19]), .ZN(n4517) );
  OAI22_X1 U4118 ( .A1(n4456), .A2(n6032), .B1(n4517), .B2(n6034), .ZN(n4535)
         );
  XNOR2_X1 U4119 ( .A(n6118), .B(op_a_i[26]), .ZN(n5808) );
  XNOR2_X1 U4120 ( .A(n5808), .B(n5856), .ZN(n4548) );
  OAI22_X1 U4121 ( .A1(n4457), .A2(n3241), .B1(n4548), .B2(n5635), .ZN(n4534)
         );
  XNOR2_X1 U4122 ( .A(n5867), .B(n5919), .ZN(n4530) );
  OAI22_X1 U4123 ( .A1(n4458), .A2(n3128), .B1(n4530), .B2(n5922), .ZN(n4515)
         );
  XNOR2_X1 U4124 ( .A(n5821), .B(n5807), .ZN(n4544) );
  OAI22_X1 U4125 ( .A1(n4459), .A2(n2867), .B1(n4544), .B2(n5809), .ZN(n4514)
         );
  HA_X1 U4126 ( .A(n4461), .B(n4460), .CO(n4513), .S(n4466) );
  FA_X1 U4127 ( .A(n4464), .B(n4463), .CI(n4462), .CO(n4524), .S(n4482) );
  FA_X1 U4128 ( .A(n4467), .B(n4466), .CI(n4465), .CO(n4523), .S(n4477) );
  FA_X1 U4129 ( .A(n4470), .B(n4469), .CI(n4468), .CO(n4552), .S(n4450) );
  FA_X1 U4130 ( .A(n4473), .B(n4472), .CI(n4471), .CO(n4551), .S(n4462) );
  FA_X1 U4131 ( .A(n4476), .B(n4475), .CI(n4474), .CO(n4550), .S(n4449) );
  FA_X1 U4132 ( .A(n4479), .B(n4478), .CI(n4477), .CO(n4506), .S(n4439) );
  FA_X1 U4133 ( .A(n4482), .B(n4481), .CI(n4480), .CO(n4505), .S(n4489) );
  AND2_X1 U4134 ( .A1(n4483), .A2(n29), .ZN(n4566) );
  INV_X1 U4135 ( .A(op_b_i[26]), .ZN(n4484) );
  NOR2_X1 U4136 ( .A1(n6119), .A2(n4484), .ZN(n4485) );
  OR2_X1 U4137 ( .A1(n4485), .A2(n6144), .ZN(n4560) );
  INV_X1 U4138 ( .A(dot_op_c_i[26]), .ZN(n4667) );
  OAI22_X1 U4139 ( .A1(n6146), .A2(n4667), .B1(n2525), .B2(n877), .ZN(n4559)
         );
  HA_X1 U4140 ( .A(n4487), .B(n4486), .CO(n4503), .S(n4436) );
  FA_X1 U4141 ( .A(n4490), .B(n4489), .CI(n4488), .CO(n4491), .S(n4403) );
  OR2_X1 U4142 ( .A1(n4491), .A2(n6145), .ZN(n4502) );
  FA_X1 U4143 ( .A(n4494), .B(n4493), .CI(n4492), .CO(n4500), .S(n4498) );
  NOR2_X1 U4144 ( .A1(n4501), .A2(n4500), .ZN(n4945) );
  NOR2_X1 U4145 ( .A1(n4941), .A2(n4945), .ZN(n5710) );
  NAND2_X1 U4146 ( .A1(n4496), .A2(n4495), .ZN(n5611) );
  INV_X1 U4147 ( .A(n5611), .ZN(n5196) );
  NAND2_X1 U4148 ( .A1(n4498), .A2(n4497), .ZN(n5197) );
  INV_X1 U4149 ( .A(n5197), .ZN(n4499) );
  AOI21_X1 U4150 ( .B1(n5198), .B2(n5196), .A(n4499), .ZN(n4942) );
  NAND2_X1 U4151 ( .A1(n4501), .A2(n4500), .ZN(n4946) );
  OAI21_X1 U4152 ( .B1(n4942), .B2(n4945), .A(n4946), .ZN(n5715) );
  AOI21_X1 U4153 ( .B1(n5614), .B2(n5710), .A(n5715), .ZN(n5626) );
  FA_X1 U4154 ( .A(n4504), .B(n4503), .CI(n4502), .CO(n5692), .S(n4565) );
  FA_X1 U4155 ( .A(n4507), .B(n4506), .CI(n4505), .CO(n5688), .S(n4561) );
  XNOR2_X1 U4156 ( .A(n22), .B(op_b_i[23]), .ZN(n5638) );
  OAI22_X1 U4157 ( .A1(n5638), .A2(n5983), .B1(n4508), .B2(n5981), .ZN(n5659)
         );
  XNOR2_X1 U4158 ( .A(n65), .B(n4123), .ZN(n5634) );
  OAI22_X1 U4159 ( .A1(n5634), .A2(n5927), .B1(n4509), .B2(n5925), .ZN(n5658)
         );
  INV_X1 U4160 ( .A(op_b_i[27]), .ZN(n4511) );
  OR2_X1 U4161 ( .A1(n6116), .A2(n4511), .ZN(n4512) );
  XOR2_X1 U4162 ( .A(op_b_i[26]), .B(op_b_i[27]), .Z(n4510) );
  NAND2_X1 U4163 ( .A1(n4510), .A2(n6038), .ZN(n6036) );
  OAI22_X1 U4164 ( .A1(n4512), .A2(n6038), .B1(n6036), .B2(n4511), .ZN(n5657)
         );
  FA_X1 U4165 ( .A(n4515), .B(n4514), .CI(n4513), .CO(n5650), .S(n4519) );
  XNOR2_X1 U4166 ( .A(n56), .B(op_b_i[25]), .ZN(n5639) );
  OAI22_X1 U4167 ( .A1(n5639), .A2(n5995), .B1(n4516), .B2(n5993), .ZN(n5654)
         );
  XNOR2_X1 U4168 ( .A(n21), .B(op_b_i[19]), .ZN(n5637) );
  OAI22_X1 U4169 ( .A1(n5637), .A2(n6034), .B1(n4517), .B2(n6032), .ZN(n5653)
         );
  XNOR2_X1 U4170 ( .A(n6116), .B(op_b_i[27]), .ZN(n4518) );
  XNOR2_X1 U4171 ( .A(n6002), .B(op_b_i[27]), .ZN(n5666) );
  OAI22_X1 U4172 ( .A1(n4518), .A2(n6036), .B1(n5666), .B2(n6038), .ZN(n5652)
         );
  FA_X1 U4173 ( .A(n4521), .B(n4520), .CI(n4519), .CO(n5679), .S(n4553) );
  FA_X1 U4174 ( .A(n4524), .B(n4523), .CI(n4522), .CO(n5678), .S(n4507) );
  FA_X1 U4175 ( .A(n4527), .B(n4526), .CI(n4525), .CO(n5648), .S(n4555) );
  XNOR2_X1 U4176 ( .A(n51), .B(op_b_i[17]), .ZN(n5633) );
  OAI22_X1 U4177 ( .A1(n5633), .A2(n5917), .B1(n4528), .B2(n5915), .ZN(n5656)
         );
  XNOR2_X1 U4178 ( .A(n54), .B(op_b_i[21]), .ZN(n5668) );
  OAI22_X1 U4179 ( .A1(n5668), .A2(n68), .B1(n4529), .B2(n5997), .ZN(n5655) );
  XNOR2_X1 U4180 ( .A(n5942), .B(n5919), .ZN(n5642) );
  OAI22_X1 U4181 ( .A1(n5642), .A2(n5922), .B1(n4530), .B2(n3128), .ZN(n5670)
         );
  FA_X1 U4182 ( .A(n4533), .B(n4532), .CI(n4531), .CO(n5669), .S(n4527) );
  FA_X1 U4183 ( .A(n4536), .B(n4535), .CI(n4534), .CO(n5677), .S(n4520) );
  FA_X1 U4184 ( .A(n4539), .B(n4538), .CI(n4537), .CO(n5676), .S(n4525) );
  FA_X1 U4185 ( .A(n4542), .B(n4541), .CI(n4540), .CO(n5675), .S(n4521) );
  XNOR2_X1 U4186 ( .A(n5924), .B(n5941), .ZN(n5674) );
  OAI22_X1 U4187 ( .A1(n5674), .A2(n26), .B1(n4543), .B2(n5943), .ZN(n5662) );
  XNOR2_X1 U4188 ( .A(n5938), .B(n5807), .ZN(n5641) );
  OAI22_X1 U4189 ( .A1(n5641), .A2(n6010), .B1(n4544), .B2(n2867), .ZN(n5661)
         );
  XNOR2_X1 U4190 ( .A(n5933), .B(n27), .ZN(n5640) );
  OAI22_X1 U4191 ( .A1(n5640), .A2(n4546), .B1(n4545), .B2(n5822), .ZN(n5660)
         );
  XNOR2_X1 U4192 ( .A(n5914), .B(op_b_i[13]), .ZN(n5672) );
  OAI22_X1 U4193 ( .A1(n5672), .A2(n72), .B1(n4547), .B2(n5934), .ZN(n5665) );
  XNOR2_X1 U4194 ( .A(n6118), .B(op_a_i[27]), .ZN(n6008) );
  XNOR2_X1 U4195 ( .A(n6008), .B(n5856), .ZN(n5636) );
  OAI22_X1 U4196 ( .A1(n5636), .A2(n5635), .B1(n4548), .B2(n3241), .ZN(n5664)
         );
  XNOR2_X1 U4197 ( .A(n5920), .B(n5811), .ZN(n5673) );
  OAI22_X1 U4198 ( .A1(n5673), .A2(n10), .B1(n4549), .B2(n2585), .ZN(n5663) );
  FA_X1 U4199 ( .A(n4552), .B(n4551), .CI(n4550), .CO(n5643), .S(n4522) );
  FA_X1 U4200 ( .A(n4555), .B(n4554), .CI(n4553), .CO(n5630), .S(n4562) );
  AND2_X1 U4201 ( .A1(n4556), .A2(n29), .ZN(n5691) );
  NOR2_X1 U4202 ( .A1(n6119), .A2(n4511), .ZN(n4557) );
  OR2_X1 U4203 ( .A1(n4557), .A2(n6144), .ZN(n5685) );
  INV_X1 U4204 ( .A(dot_op_c_i[27]), .ZN(n4881) );
  INV_X1 U4205 ( .A(op_c_i[27]), .ZN(n4558) );
  OAI22_X1 U4206 ( .A1(n6146), .A2(n4881), .B1(n2525), .B2(n4558), .ZN(n5684)
         );
  HA_X1 U4207 ( .A(n4560), .B(n4559), .CO(n5628), .S(n4504) );
  FA_X1 U4208 ( .A(n4563), .B(n4562), .CI(n4561), .CO(n4564), .S(n4483) );
  OR2_X1 U4209 ( .A1(n4564), .A2(n6142), .ZN(n5627) );
  FA_X1 U4210 ( .A(n4567), .B(n4566), .CI(n4565), .CO(n4568), .S(n4501) );
  NOR2_X1 U4211 ( .A1(n4569), .A2(n4568), .ZN(n5709) );
  INV_X1 U4212 ( .A(n5709), .ZN(n4570) );
  NAND2_X1 U4213 ( .A1(n4569), .A2(n4568), .ZN(n5712) );
  NAND2_X1 U4214 ( .A1(n4570), .A2(n5712), .ZN(n4571) );
  XOR2_X1 U4215 ( .A(n5626), .B(n4571), .Z(n4572) );
  NAND2_X1 U4216 ( .A1(n4572), .A2(n5615), .ZN(n4884) );
  FA_X1 U4217 ( .A(n4575), .B(n4574), .CI(n4573), .CO(n4762), .S(n4619) );
  FA_X1 U4218 ( .A(n4578), .B(n4577), .CI(n4576), .CO(n4647), .S(n4616) );
  XNOR2_X1 U4219 ( .A(n5076), .B(n4679), .ZN(n4662) );
  OAI22_X1 U4220 ( .A1(n4579), .A2(n4746), .B1(n4662), .B2(n4745), .ZN(n4635)
         );
  OAI21_X1 U4221 ( .B1(n1661), .B2(n5617), .A(n5114), .ZN(n4634) );
  XNOR2_X1 U4222 ( .A(n4673), .B(n1803), .ZN(n4654) );
  OAI22_X1 U4223 ( .A1(n4580), .A2(n5124), .B1(n4654), .B2(n5123), .ZN(n4633)
         );
  FA_X1 U4224 ( .A(n4583), .B(n4582), .CI(n4581), .CO(n4640), .S(n4577) );
  XNOR2_X1 U4225 ( .A(n4681), .B(n17), .ZN(n4648) );
  OAI22_X1 U4226 ( .A1(n5113), .A2(n4584), .B1(n4648), .B2(n6114), .ZN(n4690)
         );
  XNOR2_X1 U4227 ( .A(n4795), .B(n30), .ZN(n4649) );
  OAI22_X1 U4228 ( .A1(n4585), .A2(n4830), .B1(n4649), .B2(n4829), .ZN(n4689)
         );
  XNOR2_X1 U4229 ( .A(n4780), .B(n6111), .ZN(n4650) );
  OAI22_X1 U4230 ( .A1(n6125), .A2(n4586), .B1(n6123), .B2(n4650), .ZN(n4688)
         );
  XNOR2_X1 U4231 ( .A(n5083), .B(n4587), .ZN(n4659) );
  OAI22_X1 U4232 ( .A1(n4661), .A2(n4588), .B1(n4659), .B2(n4660), .ZN(n4653)
         );
  XNOR2_X1 U4233 ( .A(n4683), .B(n5078), .ZN(n4632) );
  OAI22_X1 U4234 ( .A1(n4732), .A2(n4589), .B1(n4632), .B2(n4731), .ZN(n4652)
         );
  INV_X1 U4235 ( .A(n4602), .ZN(n4651) );
  XNOR2_X1 U4236 ( .A(n4590), .B(n15), .ZN(n4591) );
  NOR2_X1 U4237 ( .A1(n4591), .A2(n5109), .ZN(n4687) );
  INV_X1 U4238 ( .A(n4592), .ZN(n4593) );
  NOR2_X1 U4239 ( .A1(n4593), .A2(n5116), .ZN(n4686) );
  XNOR2_X1 U4240 ( .A(n5085), .B(n1307), .ZN(n4628) );
  OAI22_X1 U4241 ( .A1(n4628), .A2(n4629), .B1(n4594), .B2(n4630), .ZN(n4685)
         );
  FA_X1 U4242 ( .A(n4597), .B(n4596), .CI(n4595), .CO(n4697), .S(n4614) );
  FA_X1 U4243 ( .A(n4600), .B(n4599), .CI(n4598), .CO(n4638), .S(n4611) );
  FA_X1 U4244 ( .A(n4603), .B(n4602), .CI(n4601), .CO(n4637), .S(n4609) );
  FA_X1 U4245 ( .A(n4606), .B(n4605), .CI(n4604), .CO(n4636), .S(n4612) );
  FA_X1 U4246 ( .A(n4609), .B(n4608), .CI(n4607), .CO(n4643), .S(n4615) );
  FA_X1 U4247 ( .A(n4612), .B(n4611), .CI(n4610), .CO(n4642), .S(n4617) );
  FA_X1 U4248 ( .A(n4615), .B(n4614), .CI(n4613), .CO(n4707), .S(n4575) );
  FA_X1 U4249 ( .A(n4618), .B(n4617), .CI(n4616), .CO(n4706), .S(n4620) );
  FA_X1 U4250 ( .A(n4621), .B(n4620), .CI(n4619), .CO(n4622), .S(n2265) );
  NOR2_X1 U4251 ( .A1(n4623), .A2(n4622), .ZN(n5033) );
  NOR2_X1 U4252 ( .A1(n5028), .A2(n5033), .ZN(n4625) );
  NAND2_X1 U4253 ( .A1(n5024), .A2(n4625), .ZN(n4863) );
  INV_X1 U4254 ( .A(n4863), .ZN(n4627) );
  NAND2_X1 U4255 ( .A1(n4623), .A2(n4622), .ZN(n5034) );
  OAI21_X1 U4256 ( .B1(n5033), .B2(n5027), .A(n5034), .ZN(n4624) );
  AOI21_X1 U4257 ( .B1(n5026), .B2(n4625), .A(n4624), .ZN(n4870) );
  INV_X1 U4258 ( .A(n4870), .ZN(n4626) );
  AOI21_X1 U4259 ( .B1(n5032), .B2(n4627), .A(n4626), .ZN(n4953) );
  AOI21_X1 U4260 ( .B1(n4630), .B2(n4629), .A(n4628), .ZN(n4631) );
  INV_X1 U4261 ( .A(n4631), .ZN(n4678) );
  XNOR2_X1 U4262 ( .A(n4683), .B(n5107), .ZN(n4684) );
  OAI22_X1 U4263 ( .A1(n4732), .A2(n4632), .B1(n4684), .B2(n4731), .ZN(n4677)
         );
  FA_X1 U4264 ( .A(n4635), .B(n4634), .CI(n4633), .CO(n4676), .S(n4641) );
  FA_X1 U4265 ( .A(n4638), .B(n4637), .CI(n4636), .CO(n4695), .S(n4644) );
  FA_X1 U4266 ( .A(n4641), .B(n4640), .CI(n4639), .CO(n4694), .S(n4646) );
  FA_X1 U4267 ( .A(n4644), .B(n4643), .CI(n4642), .CO(n4713), .S(n4708) );
  FA_X1 U4268 ( .A(n4647), .B(n4646), .CI(n4645), .CO(n4712), .S(n4761) );
  XNOR2_X1 U4269 ( .A(n4740), .B(n17), .ZN(n4672) );
  OAI22_X1 U4270 ( .A1(n5113), .A2(n4648), .B1(n4672), .B2(n6114), .ZN(n4665)
         );
  XNOR2_X1 U4271 ( .A(n4839), .B(n30), .ZN(n4666) );
  OAI22_X1 U4272 ( .A1(n4649), .A2(n4830), .B1(n4666), .B2(n4829), .ZN(n4664)
         );
  XNOR2_X1 U4273 ( .A(n4841), .B(n6111), .ZN(n4675) );
  OAI22_X1 U4274 ( .A1(n6125), .A2(n4650), .B1(n6123), .B2(n4675), .ZN(n4663)
         );
  FA_X1 U4275 ( .A(n4653), .B(n4652), .CI(n4651), .CO(n4704), .S(n4699) );
  XNOR2_X1 U4276 ( .A(n4742), .B(n1803), .ZN(n4668) );
  OAI22_X1 U4277 ( .A1(n4654), .A2(n5124), .B1(n4668), .B2(n5123), .ZN(n4671)
         );
  INV_X1 U4278 ( .A(n4655), .ZN(n4656) );
  NOR2_X1 U4279 ( .A1(n4656), .A2(n5116), .ZN(n4670) );
  XNOR2_X1 U4280 ( .A(n4657), .B(n15), .ZN(n4658) );
  NOR2_X1 U4281 ( .A1(n4658), .A2(n5109), .ZN(n4669) );
  OAI21_X1 U4282 ( .B1(n1661), .B2(n5204), .A(n5114), .ZN(n4693) );
  AOI21_X1 U4283 ( .B1(n4661), .B2(n4660), .A(n4659), .ZN(n4692) );
  XNOR2_X1 U4284 ( .A(n5115), .B(n4679), .ZN(n4680) );
  OAI22_X1 U4285 ( .A1(n4662), .A2(n4746), .B1(n4680), .B2(n4745), .ZN(n4691)
         );
  INV_X1 U4286 ( .A(n4692), .ZN(n4722) );
  FA_X1 U4287 ( .A(n4665), .B(n4664), .CI(n4663), .CO(n4721), .S(n4705) );
  XNOR2_X1 U4288 ( .A(n5076), .B(n30), .ZN(n4733) );
  OAI22_X1 U4289 ( .A1(n4666), .A2(n4830), .B1(n4733), .B2(n4829), .ZN(n4729)
         );
  OAI21_X1 U4290 ( .B1(n1661), .B2(n4667), .A(n5114), .ZN(n4728) );
  XNOR2_X1 U4291 ( .A(n4795), .B(n1803), .ZN(n4735) );
  OAI22_X1 U4292 ( .A1(n4668), .A2(n5124), .B1(n4735), .B2(n5123), .ZN(n4727)
         );
  FA_X1 U4293 ( .A(n4671), .B(n4670), .CI(n4669), .CO(n4719), .S(n4703) );
  XNOR2_X1 U4294 ( .A(n4780), .B(n17), .ZN(n4734) );
  OAI22_X1 U4295 ( .A1(n5113), .A2(n4672), .B1(n4734), .B2(n6114), .ZN(n4726)
         );
  INV_X1 U4296 ( .A(n4673), .ZN(n4674) );
  NOR2_X1 U4297 ( .A1(n4674), .A2(n5116), .ZN(n4725) );
  XNOR2_X1 U4298 ( .A(n5078), .B(n6111), .ZN(n4736) );
  OAI22_X1 U4299 ( .A1(n6125), .A2(n4675), .B1(n6123), .B2(n4736), .ZN(n4724)
         );
  FA_X1 U4300 ( .A(n4678), .B(n4677), .CI(n4676), .CO(n4750), .S(n4696) );
  XNOR2_X1 U4301 ( .A(n5085), .B(n4679), .ZN(n4744) );
  OAI22_X1 U4302 ( .A1(n4744), .A2(n4745), .B1(n4680), .B2(n4746), .ZN(n4739)
         );
  XNOR2_X1 U4303 ( .A(n4681), .B(n15), .ZN(n4682) );
  NOR2_X1 U4304 ( .A1(n4682), .A2(n5109), .ZN(n4738) );
  XNOR2_X1 U4305 ( .A(n5083), .B(n4683), .ZN(n4730) );
  OAI22_X1 U4306 ( .A1(n4732), .A2(n4684), .B1(n4730), .B2(n4731), .ZN(n4737)
         );
  FA_X1 U4307 ( .A(n4687), .B(n4686), .CI(n4685), .CO(n4702), .S(n4698) );
  FA_X1 U4308 ( .A(n4690), .B(n4689), .CI(n4688), .CO(n4701), .S(n4639) );
  FA_X1 U4309 ( .A(n4693), .B(n4692), .CI(n4691), .CO(n4723), .S(n4700) );
  FA_X1 U4310 ( .A(n4696), .B(n4695), .CI(n4694), .CO(n4716), .S(n4714) );
  FA_X1 U4311 ( .A(n4699), .B(n4698), .CI(n4697), .CO(n4711), .S(n4645) );
  FA_X1 U4312 ( .A(n4702), .B(n4701), .CI(n4700), .CO(n4748), .S(n4710) );
  FA_X1 U4313 ( .A(n4705), .B(n4704), .CI(n4703), .CO(n4753), .S(n4709) );
  FA_X1 U4314 ( .A(n4708), .B(n4707), .CI(n4706), .CO(n4759), .S(n4760) );
  FA_X1 U4315 ( .A(n4711), .B(n4710), .CI(n4709), .CO(n4715), .S(n4758) );
  FA_X1 U4316 ( .A(n4714), .B(n4713), .CI(n4712), .CO(n4756), .S(n4757) );
  NOR2_X1 U4317 ( .A1(n4766), .A2(n4765), .ZN(n4859) );
  FA_X1 U4318 ( .A(n4717), .B(n4716), .CI(n4715), .CO(n4805), .S(n4754) );
  FA_X1 U4319 ( .A(n4720), .B(n4719), .CI(n4718), .CO(n4802), .S(n4751) );
  FA_X1 U4320 ( .A(n4723), .B(n4722), .CI(n4721), .CO(n4801), .S(n4752) );
  FA_X1 U4321 ( .A(n4726), .B(n4725), .CI(n4724), .CO(n4779), .S(n4718) );
  FA_X1 U4322 ( .A(n4729), .B(n4728), .CI(n4727), .CO(n4778), .S(n4720) );
  OAI21_X1 U4323 ( .B1(n1661), .B2(n4881), .A(n5114), .ZN(n4787) );
  AOI21_X1 U4324 ( .B1(n4732), .B2(n4731), .A(n4730), .ZN(n4786) );
  XNOR2_X1 U4325 ( .A(n5115), .B(n30), .ZN(n4783) );
  OAI22_X1 U4326 ( .A1(n4733), .A2(n4830), .B1(n4783), .B2(n4829), .ZN(n4785)
         );
  XNOR2_X1 U4327 ( .A(n4841), .B(n17), .ZN(n4782) );
  OAI22_X1 U4328 ( .A1(n5113), .A2(n4734), .B1(n4782), .B2(n6114), .ZN(n4793)
         );
  XNOR2_X1 U4329 ( .A(n4839), .B(n1803), .ZN(n4794) );
  OAI22_X1 U4330 ( .A1(n4735), .A2(n5124), .B1(n4794), .B2(n5123), .ZN(n4792)
         );
  XNOR2_X1 U4331 ( .A(n5107), .B(n6111), .ZN(n4784) );
  OAI22_X1 U4332 ( .A1(n6125), .A2(n4736), .B1(n6123), .B2(n4784), .ZN(n4791)
         );
  FA_X1 U4333 ( .A(n4739), .B(n4738), .CI(n4737), .CO(n4798), .S(n4749) );
  XNOR2_X1 U4334 ( .A(n4740), .B(n15), .ZN(n4741) );
  NOR2_X1 U4335 ( .A1(n4741), .A2(n5109), .ZN(n4790) );
  INV_X1 U4336 ( .A(n4742), .ZN(n4743) );
  NOR2_X1 U4337 ( .A1(n4743), .A2(n5116), .ZN(n4789) );
  AOI21_X1 U4338 ( .B1(n4746), .B2(n4745), .A(n4744), .ZN(n4747) );
  INV_X1 U4339 ( .A(n4747), .ZN(n4788) );
  FA_X1 U4340 ( .A(n4750), .B(n4749), .CI(n4748), .CO(n4775), .S(n4717) );
  FA_X1 U4341 ( .A(n4753), .B(n4752), .CI(n4751), .CO(n4774), .S(n4755) );
  FA_X1 U4342 ( .A(n4756), .B(n4755), .CI(n4754), .CO(n4767), .S(n4766) );
  NOR2_X1 U4343 ( .A1(n4768), .A2(n4767), .ZN(n4873) );
  OR2_X1 U4344 ( .A1(n4859), .A2(n4873), .ZN(n4771) );
  FA_X1 U4345 ( .A(n4759), .B(n4758), .CI(n4757), .CO(n4765), .S(n4764) );
  FA_X1 U4346 ( .A(n4762), .B(n4761), .CI(n4760), .CO(n4763), .S(n4623) );
  NOR2_X1 U4347 ( .A1(n4764), .A2(n4763), .ZN(n4862) );
  NOR2_X1 U4348 ( .A1(n4771), .A2(n4862), .ZN(n4810) );
  INV_X1 U4349 ( .A(n4810), .ZN(n4773) );
  NAND2_X1 U4350 ( .A1(n4764), .A2(n4763), .ZN(n4950) );
  NAND2_X1 U4351 ( .A1(n4766), .A2(n4765), .ZN(n4864) );
  NAND2_X1 U4352 ( .A1(n4768), .A2(n4767), .ZN(n4874) );
  OAI21_X1 U4353 ( .B1(n4873), .B2(n4864), .A(n4874), .ZN(n4769) );
  INV_X1 U4354 ( .A(n4769), .ZN(n4770) );
  OAI21_X1 U4355 ( .B1(n4771), .B2(n4950), .A(n4770), .ZN(n4814) );
  INV_X1 U4356 ( .A(n4814), .ZN(n4772) );
  OAI21_X1 U4357 ( .B1(n4953), .B2(n4773), .A(n4772), .ZN(n4809) );
  FA_X1 U4358 ( .A(n4776), .B(n4775), .CI(n4774), .CO(n4852), .S(n4803) );
  FA_X1 U4359 ( .A(n4779), .B(n4778), .CI(n4777), .CO(n4824), .S(n4800) );
  XNOR2_X1 U4360 ( .A(n4780), .B(n15), .ZN(n4781) );
  NOR2_X1 U4361 ( .A1(n4781), .A2(n5109), .ZN(n4834) );
  XNOR2_X1 U4362 ( .A(n5078), .B(n17), .ZN(n4838) );
  OAI22_X1 U4363 ( .A1(n5113), .A2(n4782), .B1(n4838), .B2(n6114), .ZN(n4833)
         );
  XNOR2_X1 U4364 ( .A(n5085), .B(n30), .ZN(n4828) );
  OAI22_X1 U4365 ( .A1(n4828), .A2(n4829), .B1(n4783), .B2(n4830), .ZN(n4832)
         );
  INV_X1 U4366 ( .A(n4786), .ZN(n4849) );
  XNOR2_X1 U4367 ( .A(n5083), .B(n6111), .ZN(n4843) );
  OAI22_X1 U4368 ( .A1(n4843), .A2(n6123), .B1(n6125), .B2(n4784), .ZN(n4848)
         );
  FA_X1 U4369 ( .A(n4787), .B(n4786), .CI(n4785), .CO(n4847), .S(n4777) );
  FA_X1 U4370 ( .A(n4790), .B(n4789), .CI(n4788), .CO(n4837), .S(n4797) );
  FA_X1 U4371 ( .A(n4793), .B(n4792), .CI(n4791), .CO(n4836), .S(n4799) );
  XNOR2_X1 U4372 ( .A(n5076), .B(n1803), .ZN(n4846) );
  OAI22_X1 U4373 ( .A1(n4794), .A2(n5124), .B1(n4846), .B2(n5123), .ZN(n4827)
         );
  INV_X1 U4374 ( .A(dot_op_c_i[28]), .ZN(n5699) );
  OAI21_X1 U4375 ( .B1(n1661), .B2(n5699), .A(n5114), .ZN(n4826) );
  INV_X1 U4376 ( .A(n4795), .ZN(n4796) );
  NOR2_X1 U4377 ( .A1(n4796), .A2(n5116), .ZN(n4825) );
  FA_X1 U4378 ( .A(n4799), .B(n4798), .CI(n4797), .CO(n4820), .S(n4776) );
  FA_X1 U4379 ( .A(n4802), .B(n4801), .CI(n4800), .CO(n4819), .S(n4804) );
  FA_X1 U4380 ( .A(n4805), .B(n4804), .CI(n4803), .CO(n4806), .S(n4768) );
  OR2_X1 U4381 ( .A1(n4807), .A2(n4806), .ZN(n4813) );
  NAND2_X1 U4382 ( .A1(n4807), .A2(n4806), .ZN(n4811) );
  NAND2_X1 U4383 ( .A1(n4813), .A2(n4811), .ZN(n4808) );
  XNOR2_X1 U4384 ( .A(n4809), .B(n4808), .ZN(n5705) );
  NAND2_X1 U4385 ( .A1(n4810), .A2(n4813), .ZN(n4816) );
  NOR2_X1 U4386 ( .A1(n4863), .A2(n4816), .ZN(n4818) );
  INV_X1 U4387 ( .A(n4811), .ZN(n4812) );
  AOI21_X1 U4388 ( .B1(n4814), .B2(n4813), .A(n4812), .ZN(n4815) );
  OAI21_X1 U4389 ( .B1(n4870), .B2(n4816), .A(n4815), .ZN(n4817) );
  AOI21_X1 U4390 ( .B1(n5032), .B2(n4818), .A(n4817), .ZN(n5064) );
  FA_X1 U4391 ( .A(n4821), .B(n4820), .CI(n4819), .CO(n5067), .S(n4850) );
  FA_X1 U4392 ( .A(n4824), .B(n4823), .CI(n4822), .CO(n5066), .S(n4851) );
  FA_X1 U4393 ( .A(n4827), .B(n4826), .CI(n4825), .CO(n5082), .S(n4835) );
  AOI21_X1 U4394 ( .B1(n4830), .B2(n4829), .A(n4828), .ZN(n4831) );
  INV_X1 U4395 ( .A(n4831), .ZN(n5081) );
  FA_X1 U4396 ( .A(n4834), .B(n4833), .CI(n4832), .CO(n5080), .S(n4823) );
  FA_X1 U4397 ( .A(n4837), .B(n4836), .CI(n4835), .CO(n5069), .S(n4821) );
  XNOR2_X1 U4398 ( .A(n5107), .B(n17), .ZN(n5084) );
  OAI22_X1 U4399 ( .A1(n5113), .A2(n4838), .B1(n5084), .B2(n6114), .ZN(n5073)
         );
  INV_X1 U4400 ( .A(n4839), .ZN(n4840) );
  NOR2_X1 U4401 ( .A1(n4840), .A2(n5116), .ZN(n5072) );
  XNOR2_X1 U4402 ( .A(n4841), .B(n15), .ZN(n4842) );
  NOR2_X1 U4403 ( .A1(n4842), .A2(n5109), .ZN(n5071) );
  INV_X1 U4404 ( .A(dot_op_c_i[29]), .ZN(n5793) );
  OAI21_X1 U4405 ( .B1(n1661), .B2(n5793), .A(n5114), .ZN(n5075) );
  AOI21_X1 U4406 ( .B1(n6125), .B2(n6123), .A(n4843), .ZN(n5087) );
  XNOR2_X1 U4407 ( .A(n5115), .B(dot_op_a_i[15]), .ZN(n5086) );
  OAI22_X1 U4408 ( .A1(n4846), .A2(n5124), .B1(n5086), .B2(n5123), .ZN(n5074)
         );
  FA_X1 U4409 ( .A(n4849), .B(n4848), .CI(n4847), .CO(n5088), .S(n4822) );
  FA_X1 U4410 ( .A(n4852), .B(n4851), .CI(n4850), .CO(n4853), .S(n4807) );
  NOR2_X1 U4411 ( .A1(n4854), .A2(n4853), .ZN(n5063) );
  INV_X1 U4412 ( .A(n5063), .ZN(n4855) );
  NAND2_X1 U4413 ( .A1(n4854), .A2(n4853), .ZN(n5062) );
  NAND2_X1 U4414 ( .A1(n4855), .A2(n5062), .ZN(n4856) );
  XOR2_X1 U4415 ( .A(n5064), .B(n4856), .Z(n5797) );
  AOI22_X1 U4416 ( .A1(n6147), .A2(n5463), .B1(n5797), .B2(n5490), .ZN(n4879)
         );
  NOR2_X1 U4417 ( .A1(n4863), .A2(n4862), .ZN(n4858) );
  OAI21_X1 U4418 ( .B1(n4870), .B2(n4862), .A(n4950), .ZN(n4857) );
  AOI21_X1 U4419 ( .B1(n6127), .B2(n4858), .A(n4857), .ZN(n4861) );
  INV_X1 U4420 ( .A(n4859), .ZN(n4866) );
  NAND2_X1 U4421 ( .A1(n4866), .A2(n4864), .ZN(n4860) );
  XOR2_X1 U4422 ( .A(n4861), .B(n4860), .Z(n5381) );
  INV_X1 U4423 ( .A(n4862), .ZN(n4951) );
  NAND2_X1 U4424 ( .A1(n4951), .A2(n4866), .ZN(n4869) );
  NOR2_X1 U4425 ( .A1(n4863), .A2(n4869), .ZN(n4872) );
  INV_X1 U4426 ( .A(n4950), .ZN(n4867) );
  INV_X1 U4427 ( .A(n4864), .ZN(n4865) );
  AOI21_X1 U4428 ( .B1(n4867), .B2(n4866), .A(n4865), .ZN(n4868) );
  OAI21_X1 U4429 ( .B1(n4870), .B2(n4869), .A(n4868), .ZN(n4871) );
  AOI21_X1 U4430 ( .B1(n6127), .B2(n4872), .A(n4871), .ZN(n4877) );
  INV_X1 U4431 ( .A(n4873), .ZN(n4875) );
  NAND2_X1 U4432 ( .A1(n4875), .A2(n4874), .ZN(n4876) );
  XOR2_X1 U4433 ( .A(n4877), .B(n4876), .Z(n5462) );
  AOI22_X1 U4434 ( .A1(n5521), .A2(n5381), .B1(n5462), .B2(n5519), .ZN(n4878)
         );
  NAND2_X1 U4435 ( .A1(n4879), .A2(n4878), .ZN(n5459) );
  NAND2_X1 U4436 ( .A1(n4880), .A2(n5427), .ZN(n5701) );
  INV_X1 U4437 ( .A(n5701), .ZN(n5620) );
  INV_X1 U4438 ( .A(n5462), .ZN(n5193) );
  OAI22_X1 U4439 ( .A1(n5193), .A2(n6101), .B1(n5894), .B2(n4881), .ZN(n4882)
         );
  AOI211_X1 U4440 ( .C1(n5459), .C2(n5605), .A(n5620), .B(n4882), .ZN(n4883)
         );
  OAI211_X1 U4441 ( .C1(n5461), .C2(n5703), .A(n4884), .B(n4883), .ZN(
        result_o[27]) );
  INV_X1 U4442 ( .A(n4885), .ZN(n5583) );
  NAND2_X1 U4443 ( .A1(n4886), .A2(n5567), .ZN(n4887) );
  XOR2_X1 U4444 ( .A(n5583), .B(n4887), .Z(n4891) );
  AOI22_X1 U4445 ( .A1(n5183), .A2(n5796), .B1(n38), .B2(dot_op_c_i[20]), .ZN(
        n4888) );
  OAI211_X1 U4446 ( .C1(n4889), .C2(n6106), .A(n4888), .B(n5701), .ZN(n4890)
         );
  AOI21_X1 U4447 ( .B1(n4891), .B2(n5615), .A(n4890), .ZN(n4892) );
  OAI21_X1 U4448 ( .B1(n5703), .B2(n4893), .A(n4892), .ZN(result_o[20]) );
  INV_X1 U4449 ( .A(n5261), .ZN(n4895) );
  AOI22_X1 U4450 ( .A1(n5264), .A2(n4894), .B1(n5794), .B2(n4895), .ZN(n4897)
         );
  INV_X1 U4451 ( .A(n5512), .ZN(n5425) );
  NAND2_X1 U4452 ( .A1(n5425), .A2(n5257), .ZN(n4896) );
  OAI211_X1 U4453 ( .C1(n5507), .C2(n5344), .A(n4897), .B(n4896), .ZN(n5300)
         );
  INV_X1 U4454 ( .A(n4898), .ZN(n5562) );
  INV_X1 U4455 ( .A(n4899), .ZN(n5560) );
  INV_X1 U4456 ( .A(n5559), .ZN(n4900) );
  AOI21_X1 U4457 ( .B1(n5562), .B2(n5560), .A(n4900), .ZN(n4905) );
  INV_X1 U4458 ( .A(n4901), .ZN(n4903) );
  NAND2_X1 U4459 ( .A1(n4903), .A2(n4902), .ZN(n4904) );
  XOR2_X1 U4460 ( .A(n4905), .B(n4904), .Z(n4906) );
  NAND2_X1 U4461 ( .A1(n4906), .A2(n5615), .ZN(n4926) );
  NAND2_X1 U4462 ( .A1(n4907), .A2(n5463), .ZN(n4921) );
  NAND2_X1 U4463 ( .A1(n4909), .A2(n4908), .ZN(n4910) );
  XNOR2_X1 U4464 ( .A(n4911), .B(n4910), .ZN(n5184) );
  INV_X1 U4465 ( .A(n4912), .ZN(n5534) );
  OAI21_X1 U4466 ( .B1(n5534), .B2(n4914), .A(n4913), .ZN(n4919) );
  INV_X1 U4467 ( .A(n4915), .ZN(n4917) );
  NAND2_X1 U4468 ( .A1(n4917), .A2(n4916), .ZN(n4918) );
  XNOR2_X1 U4469 ( .A(n4919), .B(n4918), .ZN(n5549) );
  AOI22_X1 U4470 ( .A1(n5184), .A2(n5519), .B1(n5521), .B2(n5549), .ZN(n4920)
         );
  OAI211_X1 U4471 ( .C1(n4922), .C2(n5192), .A(n4921), .B(n4920), .ZN(n5298)
         );
  INV_X1 U4472 ( .A(n5184), .ZN(n5234) );
  OAI22_X1 U4473 ( .A1(n5234), .A2(n6101), .B1(n5894), .B2(n4923), .ZN(n4924)
         );
  AOI211_X1 U4474 ( .C1(n5605), .C2(n5298), .A(n4924), .B(n5620), .ZN(n4925)
         );
  OAI211_X1 U4475 ( .C1(n5703), .C2(n5300), .A(n4926), .B(n4925), .ZN(
        result_o[17]) );
  AOI21_X1 U4476 ( .B1(n5562), .B2(n4928), .A(n4927), .ZN(n5181) );
  OAI21_X1 U4477 ( .B1(n5181), .B2(n5177), .A(n5178), .ZN(n4933) );
  INV_X1 U4478 ( .A(n4929), .ZN(n4931) );
  NAND2_X1 U4479 ( .A1(n4931), .A2(n4930), .ZN(n4932) );
  XNOR2_X1 U4480 ( .A(n4933), .B(n4932), .ZN(n4938) );
  AOI22_X1 U4481 ( .A1(n4934), .A2(n5796), .B1(n38), .B2(dot_op_c_i[19]), .ZN(
        n4935) );
  OAI211_X1 U4482 ( .C1(n4936), .C2(n6106), .A(n4935), .B(n5701), .ZN(n4937)
         );
  AOI21_X1 U4483 ( .B1(n4938), .B2(n5615), .A(n4937), .ZN(n4939) );
  OAI21_X1 U4484 ( .B1(n5703), .B2(n4940), .A(n4939), .ZN(result_o[19]) );
  INV_X1 U4485 ( .A(n4941), .ZN(n4944) );
  INV_X1 U4486 ( .A(n4942), .ZN(n4943) );
  AOI21_X1 U4487 ( .B1(n5614), .B2(n4944), .A(n4943), .ZN(n4949) );
  INV_X1 U4488 ( .A(n4945), .ZN(n4947) );
  NAND2_X1 U4489 ( .A1(n4947), .A2(n4946), .ZN(n4948) );
  XOR2_X1 U4490 ( .A(n4949), .B(n4948), .Z(n4971) );
  NAND2_X1 U4491 ( .A1(n4951), .A2(n4950), .ZN(n4952) );
  XOR2_X1 U4492 ( .A(n4953), .B(n4952), .Z(n5038) );
  INV_X1 U4493 ( .A(n5038), .ZN(n5378) );
  AOI22_X1 U4494 ( .A1(n5519), .A2(n5381), .B1(n5462), .B2(n5463), .ZN(n4955)
         );
  NAND2_X1 U4495 ( .A1(n5705), .A2(n5490), .ZN(n4954) );
  OAI211_X1 U4496 ( .C1(n5378), .C2(n5376), .A(n4955), .B(n4954), .ZN(n5020)
         );
  NAND2_X1 U4497 ( .A1(n5020), .A2(n5605), .ZN(n4969) );
  AOI22_X1 U4498 ( .A1(n5381), .A2(n5796), .B1(n38), .B2(dot_op_c_i[26]), .ZN(
        n4968) );
  AOI22_X1 U4499 ( .A1(n5302), .A2(n4957), .B1(n4956), .B2(n5331), .ZN(n4961)
         );
  AOI22_X1 U4500 ( .A1(n5304), .A2(n4959), .B1(n4958), .B2(n5008), .ZN(n4960)
         );
  NAND2_X1 U4501 ( .A1(n4961), .A2(n4960), .ZN(n5345) );
  INV_X1 U4502 ( .A(n5382), .ZN(n5202) );
  AOI22_X1 U4503 ( .A1(n5302), .A2(n4963), .B1(n4962), .B2(n5304), .ZN(n4964)
         );
  NAND2_X1 U4504 ( .A1(n5897), .A2(n5257), .ZN(n4966) );
  OAI211_X1 U4505 ( .C1(n5544), .C2(n5344), .A(n5202), .B(n4966), .ZN(n4973)
         );
  NAND2_X1 U4506 ( .A1(n4973), .A2(n5622), .ZN(n4967) );
  NAND4_X1 U4507 ( .A1(n4969), .A2(n4968), .A3(n5701), .A4(n4967), .ZN(n4970)
         );
  AOI21_X1 U4508 ( .B1(n4971), .B2(n5615), .A(n4970), .ZN(n4972) );
  INV_X1 U4509 ( .A(n4972), .ZN(result_o[26]) );
  INV_X1 U4510 ( .A(n4973), .ZN(n5022) );
  NAND2_X1 U4511 ( .A1(n4974), .A2(n5008), .ZN(n4981) );
  NAND2_X1 U4512 ( .A1(n4975), .A2(n5304), .ZN(n4980) );
  NAND2_X1 U4513 ( .A1(n4976), .A2(n5331), .ZN(n4979) );
  NAND2_X1 U4514 ( .A1(n4977), .A2(n5302), .ZN(n4978) );
  NAND4_X1 U4515 ( .A1(n4981), .A2(n4980), .A3(n4979), .A4(n4978), .ZN(n5530)
         );
  INV_X1 U4516 ( .A(n5530), .ZN(n5174) );
  INV_X1 U4517 ( .A(n5158), .ZN(n5543) );
  NAND2_X1 U4518 ( .A1(n5433), .A2(n4982), .ZN(n4984) );
  INV_X1 U4519 ( .A(n4983), .ZN(n5434) );
  XNOR2_X1 U4520 ( .A(n4984), .B(n5434), .ZN(n5017) );
  NAND2_X1 U4521 ( .A1(n4985), .A2(n5008), .ZN(n4993) );
  NAND2_X1 U4522 ( .A1(n4986), .A2(n5304), .ZN(n4989) );
  NAND2_X1 U4523 ( .A1(n4987), .A2(n5302), .ZN(n4988) );
  NAND2_X1 U4524 ( .A1(n4989), .A2(n4988), .ZN(n4990) );
  AOI21_X1 U4525 ( .B1(n5331), .B2(n4991), .A(n4990), .ZN(n4992) );
  AND2_X1 U4526 ( .A1(n4993), .A2(n4992), .ZN(n5537) );
  INV_X1 U4527 ( .A(n4994), .ZN(n5442) );
  INV_X1 U4528 ( .A(n5441), .ZN(n4995) );
  NAND2_X1 U4529 ( .A1(n4995), .A2(n5440), .ZN(n4996) );
  XOR2_X1 U4530 ( .A(n5442), .B(n4996), .Z(n4997) );
  AOI22_X1 U4531 ( .A1(n4997), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[10]), 
        .ZN(n5006) );
  INV_X1 U4532 ( .A(n4998), .ZN(n5004) );
  NAND2_X1 U4533 ( .A1(n4999), .A2(n5311), .ZN(n5003) );
  AOI22_X1 U4534 ( .A1(n5001), .A2(n5304), .B1(n5302), .B2(n5000), .ZN(n5002)
         );
  OAI211_X1 U4535 ( .C1(n5004), .C2(n5307), .A(n5003), .B(n5002), .ZN(n5370)
         );
  NAND2_X1 U4536 ( .A1(n5370), .A2(n5898), .ZN(n5005) );
  OAI211_X1 U4537 ( .C1(n5537), .C2(n5477), .A(n5006), .B(n5005), .ZN(n5016)
         );
  INV_X1 U4538 ( .A(n5007), .ZN(n5014) );
  NAND2_X1 U4539 ( .A1(n5009), .A2(n5008), .ZN(n5013) );
  AOI22_X1 U4540 ( .A1(n5304), .A2(n5011), .B1(n5010), .B2(n5302), .ZN(n5012)
         );
  OAI211_X1 U4541 ( .C1(n5014), .C2(n5307), .A(n5013), .B(n5012), .ZN(n5539)
         );
  INV_X1 U4542 ( .A(n5539), .ZN(n5372) );
  NOR2_X1 U4543 ( .A1(n5372), .A2(n5400), .ZN(n5015) );
  AOI211_X1 U4544 ( .C1(n5017), .C2(n5615), .A(n5016), .B(n5015), .ZN(n5018)
         );
  OAI21_X1 U4545 ( .B1(n5174), .B2(n5543), .A(n5018), .ZN(n5019) );
  AOI21_X1 U4546 ( .B1(n38), .B2(n5020), .A(n5019), .ZN(n5021) );
  OAI21_X1 U4547 ( .B1(n5022), .B2(n5553), .A(n5021), .ZN(result_o[10]) );
  OAI22_X1 U4548 ( .A1(n5157), .A2(n5386), .B1(n5431), .B2(n5344), .ZN(n5023)
         );
  INV_X1 U4549 ( .A(n5604), .ZN(n5061) );
  INV_X1 U4550 ( .A(n5024), .ZN(n5025) );
  NOR2_X1 U4551 ( .A1(n5025), .A2(n5028), .ZN(n5031) );
  INV_X1 U4552 ( .A(n5026), .ZN(n5029) );
  OAI21_X1 U4553 ( .B1(n5029), .B2(n5028), .A(n5027), .ZN(n5030) );
  AOI21_X1 U4554 ( .B1(n6127), .B2(n5031), .A(n5030), .ZN(n5037) );
  INV_X1 U4555 ( .A(n5033), .ZN(n5035) );
  NAND2_X1 U4556 ( .A1(n5035), .A2(n5034), .ZN(n5036) );
  XOR2_X1 U4557 ( .A(n5037), .B(n5036), .Z(n5350) );
  AOI22_X1 U4558 ( .A1(n5521), .A2(n5588), .B1(n5350), .B2(n5463), .ZN(n5040)
         );
  AOI22_X1 U4559 ( .A1(n5490), .A2(n5038), .B1(n5602), .B2(n5519), .ZN(n5039)
         );
  NAND2_X1 U4560 ( .A1(n5040), .A2(n5039), .ZN(n5606) );
  NAND2_X1 U4561 ( .A1(n5164), .A2(n5158), .ZN(n5058) );
  NAND2_X1 U4562 ( .A1(n5042), .A2(n5041), .ZN(n5044) );
  XNOR2_X1 U4563 ( .A(n5044), .B(n5043), .ZN(n5054) );
  NAND2_X1 U4564 ( .A1(n5045), .A2(n5898), .ZN(n5052) );
  NAND2_X1 U4565 ( .A1(n5047), .A2(n5046), .ZN(n5049) );
  XNOR2_X1 U4566 ( .A(n5049), .B(n5048), .ZN(n5050) );
  AOI22_X1 U4567 ( .A1(n5050), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[7]), 
        .ZN(n5051) );
  NAND2_X1 U4568 ( .A1(n5052), .A2(n5051), .ZN(n5053) );
  AOI21_X1 U4569 ( .B1(n5054), .B2(n5615), .A(n5053), .ZN(n5057) );
  NAND2_X1 U4570 ( .A1(n5439), .A2(n5529), .ZN(n5056) );
  NAND2_X1 U4571 ( .A1(n5449), .A2(n5540), .ZN(n5055) );
  NAND4_X1 U4572 ( .A1(n5058), .A2(n5057), .A3(n5056), .A4(n5055), .ZN(n5059)
         );
  AOI21_X1 U4573 ( .B1(n5606), .B2(n38), .A(n5059), .ZN(n5060) );
  OAI21_X1 U4574 ( .B1(n5061), .B2(n5553), .A(n5060), .ZN(result_o[7]) );
  OAI21_X1 U4575 ( .B1(n5064), .B2(n5063), .A(n5062), .ZN(n5097) );
  FA_X1 U4576 ( .A(n5067), .B(n5066), .CI(n5065), .CO(n5092), .S(n4854) );
  FA_X1 U4577 ( .A(n5070), .B(n5069), .CI(n5068), .CO(n5100), .S(n5065) );
  FA_X1 U4578 ( .A(n5073), .B(n5072), .CI(n5071), .CO(n5136), .S(n5090) );
  FA_X1 U4579 ( .A(n5075), .B(n5087), .CI(n5074), .CO(n5135), .S(n5089) );
  INV_X1 U4580 ( .A(n5076), .ZN(n5077) );
  NOR2_X1 U4581 ( .A1(n5077), .A2(n5116), .ZN(n5103) );
  INV_X1 U4582 ( .A(dot_op_c_i[30]), .ZN(n5893) );
  OAI21_X1 U4583 ( .B1(n1661), .B2(n5893), .A(n5114), .ZN(n5102) );
  XNOR2_X1 U4584 ( .A(n5078), .B(n15), .ZN(n5079) );
  NOR2_X1 U4585 ( .A1(n5079), .A2(n5109), .ZN(n5101) );
  FA_X1 U4586 ( .A(n5082), .B(n5081), .CI(n5080), .CO(n5139), .S(n5070) );
  XNOR2_X1 U4587 ( .A(n5083), .B(n17), .ZN(n5111) );
  OAI22_X1 U4588 ( .A1(n5111), .A2(n6114), .B1(n5113), .B2(n5084), .ZN(n5106)
         );
  XNOR2_X1 U4589 ( .A(n5085), .B(dot_op_a_i[15]), .ZN(n5122) );
  OAI22_X1 U4590 ( .A1(n5122), .A2(n5123), .B1(n5086), .B2(n5124), .ZN(n5105)
         );
  INV_X1 U4591 ( .A(n5087), .ZN(n5104) );
  FA_X1 U4592 ( .A(n5090), .B(n5089), .CI(n5088), .CO(n5137), .S(n5068) );
  OR2_X1 U4593 ( .A1(n5092), .A2(n5091), .ZN(n5096) );
  NAND2_X1 U4594 ( .A1(n5092), .A2(n5091), .ZN(n5094) );
  NAND2_X1 U4595 ( .A1(n5096), .A2(n5094), .ZN(n5093) );
  XNOR2_X1 U4596 ( .A(n5097), .B(n5093), .ZN(n5520) );
  INV_X1 U4597 ( .A(n5094), .ZN(n5095) );
  FA_X1 U4598 ( .A(n5100), .B(n5099), .CI(n5098), .CO(n5145), .S(n5091) );
  FA_X1 U4599 ( .A(n5103), .B(n5102), .CI(n5101), .CO(n5133), .S(n5134) );
  FA_X1 U4600 ( .A(n5106), .B(n5105), .CI(n5104), .CO(n5131), .S(n5138) );
  XNOR2_X1 U4601 ( .A(n15), .B(n5107), .ZN(n5110) );
  NOR2_X1 U4602 ( .A1(n5110), .A2(n5109), .ZN(n5129) );
  AOI21_X1 U4603 ( .B1(n5113), .B2(n6114), .A(n5111), .ZN(n5121) );
  INV_X1 U4604 ( .A(dot_op_c_i[31]), .ZN(n6076) );
  OAI21_X1 U4605 ( .B1(n1661), .B2(n6076), .A(n5114), .ZN(n5119) );
  INV_X1 U4606 ( .A(n5115), .ZN(n5117) );
  NOR2_X1 U4607 ( .A1(n5117), .A2(n5116), .ZN(n5118) );
  XOR2_X1 U4608 ( .A(n5119), .B(n5118), .Z(n5120) );
  XOR2_X1 U4609 ( .A(n5121), .B(n5120), .Z(n5127) );
  AOI21_X1 U4610 ( .B1(n5124), .B2(n5123), .A(n5122), .ZN(n5125) );
  INV_X1 U4611 ( .A(n5125), .ZN(n5126) );
  XOR2_X1 U4612 ( .A(n5127), .B(n5126), .Z(n5128) );
  XOR2_X1 U4613 ( .A(n5129), .B(n5128), .Z(n5130) );
  XOR2_X1 U4614 ( .A(n5131), .B(n5130), .Z(n5132) );
  XOR2_X1 U4615 ( .A(n5133), .B(n5132), .Z(n5143) );
  FA_X1 U4616 ( .A(n5136), .B(n5135), .CI(n5134), .CO(n5141), .S(n5099) );
  FA_X1 U4617 ( .A(n5139), .B(n5138), .CI(n5137), .CO(n5140), .S(n5098) );
  XOR2_X1 U4618 ( .A(n5141), .B(n5140), .Z(n5142) );
  XOR2_X1 U4619 ( .A(n5143), .B(n5142), .Z(n5144) );
  XOR2_X1 U4620 ( .A(n5145), .B(n5144), .Z(n5146) );
  INV_X1 U4621 ( .A(n5522), .ZN(n6102) );
  NOR2_X1 U4622 ( .A1(n6102), .A2(n5521), .ZN(n5148) );
  AOI21_X1 U4623 ( .B1(n5521), .B2(n5520), .A(n5148), .ZN(n6107) );
  INV_X1 U4624 ( .A(n5149), .ZN(n5493) );
  OAI21_X1 U4625 ( .B1(n5493), .B2(n5151), .A(n5150), .ZN(n5528) );
  AOI21_X1 U4626 ( .B1(n5528), .B2(n5526), .A(n5152), .ZN(n5156) );
  NAND2_X1 U4627 ( .A1(n5154), .A2(n5153), .ZN(n5155) );
  XOR2_X1 U4628 ( .A(n5156), .B(n5155), .Z(n5170) );
  OR2_X1 U4629 ( .A1(n2829), .A2(n5384), .ZN(n5702) );
  NOR2_X1 U4630 ( .A1(n5702), .A2(n5553), .ZN(n5523) );
  AOI22_X1 U4631 ( .A1(n5158), .A2(n5157), .B1(n5431), .B2(n5529), .ZN(n5168)
         );
  OAI21_X1 U4632 ( .B1(n5534), .B2(n5159), .A(n5531), .ZN(n5163) );
  NAND2_X1 U4633 ( .A1(n5161), .A2(n5160), .ZN(n5162) );
  XNOR2_X1 U4634 ( .A(n5163), .B(n5162), .ZN(n5231) );
  AOI22_X1 U4635 ( .A1(n5231), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[15]), 
        .ZN(n5167) );
  NAND2_X1 U4636 ( .A1(n5164), .A2(n5540), .ZN(n5166) );
  NAND2_X1 U4637 ( .A1(n5439), .A2(n5898), .ZN(n5165) );
  NAND4_X1 U4638 ( .A1(n5168), .A2(n5167), .A3(n5166), .A4(n5165), .ZN(n5169)
         );
  AOI211_X1 U4639 ( .C1(n5170), .C2(n5615), .A(n5523), .B(n5169), .ZN(n5173)
         );
  AND2_X1 U4640 ( .A1(n5427), .A2(n5384), .ZN(n5524) );
  NAND2_X1 U4641 ( .A1(n5171), .A2(n5524), .ZN(n5172) );
  OAI211_X1 U4642 ( .C1(n6107), .C2(n5894), .A(n5173), .B(n5172), .ZN(
        result_o[15]) );
  AOI22_X1 U4643 ( .A1(n5544), .A2(n5264), .B1(n5372), .B2(n5384), .ZN(n5176)
         );
  NAND2_X1 U4644 ( .A1(n5174), .A2(n5257), .ZN(n5175) );
  OAI211_X1 U4645 ( .C1(n5261), .C2(n5897), .A(n5176), .B(n5175), .ZN(n5343)
         );
  INV_X1 U4646 ( .A(n5177), .ZN(n5179) );
  NAND2_X1 U4647 ( .A1(n5179), .A2(n5178), .ZN(n5180) );
  XOR2_X1 U4648 ( .A(n5181), .B(n5180), .Z(n5182) );
  NAND2_X1 U4649 ( .A1(n5182), .A2(n5615), .ZN(n5191) );
  AOI22_X1 U4650 ( .A1(n5183), .A2(n5490), .B1(n5519), .B2(n4907), .ZN(n5186)
         );
  AOI22_X1 U4651 ( .A1(n4934), .A2(n5463), .B1(n5521), .B2(n5184), .ZN(n5185)
         );
  NAND2_X1 U4652 ( .A1(n5186), .A2(n5185), .ZN(n5341) );
  OAI22_X1 U4653 ( .A1(n5188), .A2(n6101), .B1(n5894), .B2(n5187), .ZN(n5189)
         );
  AOI211_X1 U4654 ( .C1(n5605), .C2(n5341), .A(n5189), .B(n5620), .ZN(n5190)
         );
  OAI211_X1 U4655 ( .C1(n5703), .C2(n5343), .A(n5191), .B(n5190), .ZN(
        result_o[18]) );
  NOR2_X1 U4656 ( .A1(n5193), .A2(n5192), .ZN(n5195) );
  INV_X1 U4657 ( .A(n5350), .ZN(n5618) );
  OAI22_X1 U4658 ( .A1(n5378), .A2(n5465), .B1(n5618), .B2(n5376), .ZN(n5194)
         );
  AOI211_X1 U4659 ( .C1(n5381), .C2(n5463), .A(n5195), .B(n5194), .ZN(n5430)
         );
  AOI21_X1 U4660 ( .B1(n5614), .B2(n5612), .A(n5196), .ZN(n5200) );
  NAND2_X1 U4661 ( .A1(n5198), .A2(n5197), .ZN(n5199) );
  XOR2_X1 U4662 ( .A(n5200), .B(n5199), .Z(n5201) );
  NAND2_X1 U4663 ( .A1(n5201), .A2(n5615), .ZN(n5207) );
  OAI211_X1 U4664 ( .C1(n4894), .C2(n5344), .A(n5203), .B(n5202), .ZN(n5428)
         );
  OAI22_X1 U4665 ( .A1(n5378), .A2(n6101), .B1(n5894), .B2(n5204), .ZN(n5205)
         );
  AOI211_X1 U4666 ( .C1(n5622), .C2(n5428), .A(n5620), .B(n5205), .ZN(n5206)
         );
  OAI211_X1 U4667 ( .C1(n5430), .C2(n6106), .A(n5207), .B(n5206), .ZN(
        result_o[25]) );
  INV_X1 U4668 ( .A(n109), .ZN(n5208) );
  INV_X1 U4669 ( .A(ex_ready_i), .ZN(n5209) );
  OAI21_X1 U4670 ( .B1(n5209), .B2(n109), .A(mulh_CS[2]), .ZN(n5211) );
  NAND2_X1 U4671 ( .A1(n5211), .A2(n5210), .ZN(n466) );
  NAND3_X1 U4672 ( .A1(n6108), .A2(operator_i[2]), .A3(enable_i), .ZN(n5213)
         );
  NOR3_X1 U4673 ( .A1(n5213), .A2(n5212), .A3(operator_i[0]), .ZN(n5217) );
  INV_X1 U4674 ( .A(n5218), .ZN(n5226) );
  NOR3_X1 U4675 ( .A1(n5217), .A2(mulh_CS[0]), .A3(n5226), .ZN(n5216) );
  NOR2_X1 U4676 ( .A1(n5216), .A2(n5215), .ZN(n467) );
  NOR2_X1 U4677 ( .A1(n5217), .A2(n109), .ZN(ready_o) );
  NAND2_X1 U4678 ( .A1(n5218), .A2(mulh_carry_q), .ZN(n5228) );
  AOI21_X1 U4679 ( .B1(n5221), .B2(n5220), .A(n5219), .ZN(n5225) );
  NAND2_X1 U4680 ( .A1(n5223), .A2(n5222), .ZN(n5224) );
  XOR2_X1 U4681 ( .A(n5225), .B(n5224), .Z(n5552) );
  NAND3_X1 U4682 ( .A1(n5552), .A2(n5226), .A3(n6109), .ZN(n5227) );
  OAI21_X1 U4683 ( .B1(ex_ready_i), .B2(n5228), .A(n5227), .ZN(n464) );
  INV_X1 U4684 ( .A(n5264), .ZN(n5229) );
  INV_X1 U4685 ( .A(n5230), .ZN(n5566) );
  NAND2_X1 U4686 ( .A1(n4907), .A2(n5490), .ZN(n5233) );
  AOI22_X1 U4687 ( .A1(n5521), .A2(n5231), .B1(n5549), .B2(n5519), .ZN(n5232)
         );
  OAI211_X1 U4688 ( .C1(n5234), .C2(n5488), .A(n5233), .B(n5232), .ZN(n5558)
         );
  INV_X1 U4689 ( .A(n5524), .ZN(n5515) );
  FA_X1 U4690 ( .A(n5237), .B(n5236), .CI(n5235), .CO(n5287), .S(n5267) );
  FA_X1 U4691 ( .A(n5240), .B(n5239), .CI(n5238), .CO(n5281), .S(n5241) );
  AOI22_X1 U4692 ( .A1(n5241), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[0]), 
        .ZN(n5242) );
  INV_X1 U4693 ( .A(n5242), .ZN(n5266) );
  INV_X1 U4694 ( .A(n5328), .ZN(n5271) );
  INV_X1 U4695 ( .A(n5243), .ZN(n5245) );
  NAND2_X1 U4696 ( .A1(n5245), .A2(n5244), .ZN(n5246) );
  XOR2_X1 U4697 ( .A(n5247), .B(n5246), .Z(n5326) );
  NOR2_X1 U4698 ( .A1(n5326), .A2(n5307), .ZN(n5256) );
  NAND2_X1 U4699 ( .A1(n5249), .A2(n5248), .ZN(n5251) );
  XNOR2_X1 U4700 ( .A(n5251), .B(n5250), .ZN(n5272) );
  FA_X1 U4701 ( .A(n5253), .B(op_c_i[0]), .CI(n5252), .CO(n5250), .S(n5254) );
  OAI22_X1 U4702 ( .A1(n5272), .A2(n5327), .B1(n5254), .B2(n5325), .ZN(n5255)
         );
  AOI211_X1 U4703 ( .C1(n5271), .C2(n5311), .A(n5256), .B(n5255), .ZN(n5260)
         );
  NAND2_X1 U4704 ( .A1(n5258), .A2(n5257), .ZN(n5259) );
  OAI211_X1 U4705 ( .C1(n5260), .C2(n5344), .A(n5259), .B(n5622), .ZN(n5263)
         );
  NOR2_X1 U4706 ( .A1(n5474), .A2(n5261), .ZN(n5262) );
  AOI211_X1 U4707 ( .C1(n5399), .C2(n5264), .A(n5263), .B(n5262), .ZN(n5265)
         );
  AOI211_X1 U4708 ( .C1(n5267), .C2(n5615), .A(n5266), .B(n5265), .ZN(n5268)
         );
  OAI21_X1 U4709 ( .B1(n5551), .B2(n5515), .A(n5268), .ZN(n5269) );
  AOI21_X1 U4710 ( .B1(n38), .B2(n5558), .A(n5269), .ZN(n5270) );
  OAI21_X1 U4711 ( .B1(n5566), .B2(n5553), .A(n5270), .ZN(result_o[0]) );
  NAND2_X1 U4712 ( .A1(n5271), .A2(n5331), .ZN(n5276) );
  INV_X1 U4713 ( .A(n5326), .ZN(n5274) );
  OAI21_X1 U4714 ( .B1(n5272), .B2(n5325), .A(n5898), .ZN(n5273) );
  AOI21_X1 U4715 ( .B1(n5274), .B2(n5304), .A(n5273), .ZN(n5275) );
  OAI211_X1 U4716 ( .C1(n5277), .C2(n5334), .A(n5276), .B(n5275), .ZN(n5292)
         );
  INV_X1 U4717 ( .A(n5278), .ZN(n5280) );
  NAND2_X1 U4718 ( .A1(n5280), .A2(n5279), .ZN(n5282) );
  XNOR2_X1 U4719 ( .A(n5282), .B(n5281), .ZN(n5283) );
  AOI22_X1 U4720 ( .A1(n5283), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[1]), 
        .ZN(n5291) );
  INV_X1 U4721 ( .A(n5284), .ZN(n5286) );
  NAND2_X1 U4722 ( .A1(n5286), .A2(n5285), .ZN(n5288) );
  XNOR2_X1 U4723 ( .A(n5288), .B(n5287), .ZN(n5289) );
  NAND2_X1 U4724 ( .A1(n5289), .A2(n5615), .ZN(n5290) );
  NAND3_X1 U4725 ( .A1(n5292), .A2(n5291), .A3(n5290), .ZN(n5295) );
  NOR2_X1 U4726 ( .A1(n5293), .A2(n5477), .ZN(n5294) );
  AOI211_X1 U4727 ( .C1(n5418), .C2(n5529), .A(n5295), .B(n5294), .ZN(n5296)
         );
  OAI21_X1 U4728 ( .B1(n5510), .B2(n5543), .A(n5296), .ZN(n5297) );
  AOI21_X1 U4729 ( .B1(n5298), .B2(n38), .A(n5297), .ZN(n5299) );
  OAI21_X1 U4730 ( .B1(n5300), .B2(n5553), .A(n5299), .ZN(result_o[1]) );
  INV_X1 U4731 ( .A(n5301), .ZN(n5308) );
  AOI22_X1 U4732 ( .A1(n5305), .A2(n5304), .B1(n5303), .B2(n5302), .ZN(n5306)
         );
  OAI21_X1 U4733 ( .B1(n5308), .B2(n5307), .A(n5306), .ZN(n5309) );
  AOI21_X1 U4734 ( .B1(n5311), .B2(n5310), .A(n5309), .ZN(n5367) );
  NAND2_X1 U4735 ( .A1(n5313), .A2(n5312), .ZN(n5315) );
  XNOR2_X1 U4736 ( .A(n5315), .B(n5314), .ZN(n5324) );
  INV_X1 U4737 ( .A(n5316), .ZN(n5318) );
  NAND2_X1 U4738 ( .A1(n5318), .A2(n5317), .ZN(n5320) );
  XOR2_X1 U4739 ( .A(n5320), .B(n5319), .Z(n5321) );
  AOI22_X1 U4740 ( .A1(n5321), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[2]), 
        .ZN(n5322) );
  INV_X1 U4741 ( .A(n5322), .ZN(n5323) );
  AOI21_X1 U4742 ( .B1(n5324), .B2(n5615), .A(n5323), .ZN(n5337) );
  OAI21_X1 U4743 ( .B1(n5326), .B2(n5325), .A(n5898), .ZN(n5330) );
  NOR2_X1 U4744 ( .A1(n5328), .A2(n5327), .ZN(n5329) );
  AOI211_X1 U4745 ( .C1(n5332), .C2(n5331), .A(n5330), .B(n5329), .ZN(n5333)
         );
  OAI21_X1 U4746 ( .B1(n5335), .B2(n5334), .A(n5333), .ZN(n5336) );
  OAI211_X1 U4747 ( .C1(n5367), .C2(n5477), .A(n5337), .B(n5336), .ZN(n5338)
         );
  AOI21_X1 U4748 ( .B1(n5529), .B2(n5370), .A(n5338), .ZN(n5339) );
  OAI21_X1 U4749 ( .B1(n5537), .B2(n5543), .A(n5339), .ZN(n5340) );
  AOI21_X1 U4750 ( .B1(n5341), .B2(n38), .A(n5340), .ZN(n5342) );
  OAI21_X1 U4751 ( .B1(n5343), .B2(n5553), .A(n5342), .ZN(result_o[2]) );
  INV_X1 U4752 ( .A(n5897), .ZN(n5349) );
  OAI22_X1 U4753 ( .A1(n5345), .A2(n5386), .B1(n5344), .B2(n5530), .ZN(n5347)
         );
  AOI211_X1 U4754 ( .C1(n5349), .C2(n5348), .A(n5347), .B(n5346), .ZN(n5587)
         );
  INV_X1 U4755 ( .A(n5587), .ZN(n5375) );
  AOI22_X1 U4756 ( .A1(n5519), .A2(n5588), .B1(n5602), .B2(n5463), .ZN(n5352)
         );
  AOI22_X1 U4757 ( .A1(n5350), .A2(n5490), .B1(n5521), .B2(n5573), .ZN(n5351)
         );
  NAND2_X1 U4758 ( .A1(n5352), .A2(n5351), .ZN(n5589) );
  INV_X1 U4759 ( .A(n5353), .ZN(n5355) );
  NAND2_X1 U4760 ( .A1(n5355), .A2(n5354), .ZN(n5357) );
  XOR2_X1 U4761 ( .A(n5357), .B(n5356), .Z(n5358) );
  NAND2_X1 U4762 ( .A1(n5358), .A2(n5615), .ZN(n5366) );
  INV_X1 U4763 ( .A(n5359), .ZN(n5361) );
  NAND2_X1 U4764 ( .A1(n5361), .A2(n5360), .ZN(n5363) );
  XOR2_X1 U4765 ( .A(n5363), .B(n5362), .Z(n5364) );
  AOI22_X1 U4766 ( .A1(n5364), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[6]), 
        .ZN(n5365) );
  OAI211_X1 U4767 ( .C1(n5367), .C2(n6095), .A(n5366), .B(n5365), .ZN(n5369)
         );
  NOR2_X1 U4768 ( .A1(n5537), .A2(n5400), .ZN(n5368) );
  AOI211_X1 U4769 ( .C1(n5540), .C2(n5370), .A(n5369), .B(n5368), .ZN(n5371)
         );
  OAI21_X1 U4770 ( .B1(n5372), .B2(n5543), .A(n5371), .ZN(n5373) );
  AOI21_X1 U4771 ( .B1(n5589), .B2(n38), .A(n5373), .ZN(n5374) );
  OAI21_X1 U4772 ( .B1(n5375), .B2(n5553), .A(n5374), .ZN(result_o[6]) );
  NOR2_X1 U4773 ( .A1(n5377), .A2(n5376), .ZN(n5380) );
  OAI22_X1 U4774 ( .A1(n5378), .A2(n5488), .B1(n5618), .B2(n5465), .ZN(n5379)
         );
  AOI211_X1 U4775 ( .C1(n5381), .C2(n5490), .A(n5380), .B(n5379), .ZN(n5625)
         );
  AOI21_X1 U4776 ( .B1(n5384), .B2(n5383), .A(n5382), .ZN(n5385) );
  OAI21_X1 U4777 ( .B1(n5700), .B2(n5386), .A(n5385), .ZN(n5621) );
  INV_X1 U4778 ( .A(n5387), .ZN(n5389) );
  NAND2_X1 U4779 ( .A1(n5389), .A2(n5388), .ZN(n5391) );
  XOR2_X1 U4780 ( .A(n5391), .B(n5390), .Z(n5392) );
  NAND2_X1 U4781 ( .A1(n5392), .A2(n5615), .ZN(n5398) );
  NAND2_X1 U4782 ( .A1(n5411), .A2(n5393), .ZN(n5395) );
  INV_X1 U4783 ( .A(n5394), .ZN(n5412) );
  XNOR2_X1 U4784 ( .A(n5395), .B(n5412), .ZN(n5396) );
  AOI22_X1 U4785 ( .A1(n5396), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[8]), 
        .ZN(n5397) );
  OAI211_X1 U4786 ( .C1(n5399), .C2(n6095), .A(n5398), .B(n5397), .ZN(n5402)
         );
  NOR2_X1 U4787 ( .A1(n5551), .A2(n5400), .ZN(n5401) );
  AOI211_X1 U4788 ( .C1(n5540), .C2(n5474), .A(n5402), .B(n5401), .ZN(n5403)
         );
  OAI21_X1 U4789 ( .B1(n5481), .B2(n5543), .A(n5403), .ZN(n5404) );
  AOI21_X1 U4790 ( .B1(n5427), .B2(n5621), .A(n5404), .ZN(n5405) );
  OAI21_X1 U4791 ( .B1(n5625), .B2(n5894), .A(n5405), .ZN(result_o[8]) );
  NAND2_X1 U4792 ( .A1(n5407), .A2(n5406), .ZN(n5409) );
  XNOR2_X1 U4793 ( .A(n5409), .B(n5408), .ZN(n5422) );
  AOI21_X1 U4794 ( .B1(n5412), .B2(n5411), .A(n5410), .ZN(n5416) );
  NAND2_X1 U4795 ( .A1(n5414), .A2(n5413), .ZN(n5415) );
  XOR2_X1 U4796 ( .A(n5416), .B(n5415), .Z(n5417) );
  AOI22_X1 U4797 ( .A1(n5417), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[9]), 
        .ZN(n5420) );
  NAND2_X1 U4798 ( .A1(n5418), .A2(n5898), .ZN(n5419) );
  OAI211_X1 U4799 ( .C1(n5510), .C2(n5477), .A(n5420), .B(n5419), .ZN(n5421)
         );
  AOI21_X1 U4800 ( .B1(n5422), .B2(n5615), .A(n5421), .ZN(n5424) );
  NAND2_X1 U4801 ( .A1(n5507), .A2(n5529), .ZN(n5423) );
  OAI211_X1 U4802 ( .C1(n5425), .C2(n5543), .A(n5424), .B(n5423), .ZN(n5426)
         );
  AOI21_X1 U4803 ( .B1(n5428), .B2(n5427), .A(n5426), .ZN(n5429) );
  OAI21_X1 U4804 ( .B1(n5430), .B2(n5894), .A(n5429), .ZN(result_o[9]) );
  INV_X1 U4805 ( .A(n5431), .ZN(n5457) );
  AOI21_X1 U4806 ( .B1(n5434), .B2(n5433), .A(n5432), .ZN(n5438) );
  NAND2_X1 U4807 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  XOR2_X1 U4808 ( .A(n5438), .B(n5437), .Z(n5454) );
  INV_X1 U4809 ( .A(n5439), .ZN(n5452) );
  OAI21_X1 U4810 ( .B1(n5442), .B2(n5441), .A(n5440), .ZN(n5447) );
  INV_X1 U4811 ( .A(n5443), .ZN(n5445) );
  NAND2_X1 U4812 ( .A1(n5445), .A2(n5444), .ZN(n5446) );
  XNOR2_X1 U4813 ( .A(n5447), .B(n5446), .ZN(n5448) );
  AOI22_X1 U4814 ( .A1(n5448), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[11]), 
        .ZN(n5451) );
  NAND2_X1 U4815 ( .A1(n5449), .A2(n5898), .ZN(n5450) );
  OAI211_X1 U4816 ( .C1(n5452), .C2(n5477), .A(n5451), .B(n5450), .ZN(n5453)
         );
  AOI21_X1 U4817 ( .B1(n5454), .B2(n5615), .A(n5453), .ZN(n5456) );
  NAND2_X1 U4818 ( .A1(n5164), .A2(n5529), .ZN(n5455) );
  OAI211_X1 U4819 ( .C1(n5457), .C2(n5543), .A(n5456), .B(n5455), .ZN(n5458)
         );
  AOI21_X1 U4820 ( .B1(n5459), .B2(n38), .A(n5458), .ZN(n5460) );
  OAI21_X1 U4821 ( .B1(n5461), .B2(n5553), .A(n5460), .ZN(result_o[11]) );
  INV_X1 U4822 ( .A(n5705), .ZN(n5466) );
  AOI22_X1 U4823 ( .A1(n5797), .A2(n5463), .B1(n5462), .B2(n5521), .ZN(n5464)
         );
  OAI21_X1 U4824 ( .B1(n5466), .B2(n5465), .A(n5464), .ZN(n5467) );
  AOI21_X1 U4825 ( .B1(n5490), .B2(n5520), .A(n5467), .ZN(n5708) );
  NAND2_X1 U4826 ( .A1(n5468), .A2(n5491), .ZN(n5469) );
  XOR2_X1 U4827 ( .A(n5493), .B(n5469), .Z(n5480) );
  INV_X1 U4828 ( .A(n5470), .ZN(n5501) );
  NAND2_X1 U4829 ( .A1(n5500), .A2(n5471), .ZN(n5472) );
  XNOR2_X1 U4830 ( .A(n5501), .B(n5472), .ZN(n5473) );
  AOI22_X1 U4831 ( .A1(n5473), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[12]), 
        .ZN(n5476) );
  NAND2_X1 U4832 ( .A1(n5474), .A2(n5898), .ZN(n5475) );
  OAI211_X1 U4833 ( .C1(n5551), .C2(n5477), .A(n5476), .B(n5475), .ZN(n5479)
         );
  NOR2_X1 U4834 ( .A1(n5700), .A2(n5515), .ZN(n5478) );
  AOI211_X1 U4835 ( .C1(n5480), .C2(n5615), .A(n5479), .B(n5478), .ZN(n5486)
         );
  INV_X1 U4836 ( .A(n5481), .ZN(n5484) );
  NOR2_X1 U4837 ( .A1(n5482), .A2(n5543), .ZN(n5483) );
  AOI211_X1 U4838 ( .C1(n5529), .C2(n5484), .A(n5523), .B(n5483), .ZN(n5485)
         );
  OAI211_X1 U4839 ( .C1(n5708), .C2(n5894), .A(n5486), .B(n5485), .ZN(
        result_o[12]) );
  INV_X1 U4840 ( .A(n5520), .ZN(n5895) );
  AOI22_X1 U4841 ( .A1(n6147), .A2(n5521), .B1(n5797), .B2(n5519), .ZN(n5487)
         );
  OAI21_X1 U4842 ( .B1(n5895), .B2(n5488), .A(n5487), .ZN(n5489) );
  AOI21_X1 U4843 ( .B1(n5522), .B2(n5490), .A(n5489), .ZN(n5800) );
  OAI21_X1 U4844 ( .B1(n5493), .B2(n5492), .A(n5491), .ZN(n5497) );
  NAND2_X1 U4845 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  XNOR2_X1 U4846 ( .A(n5497), .B(n5496), .ZN(n5498) );
  NAND2_X1 U4847 ( .A1(n5498), .A2(n5615), .ZN(n5514) );
  AOI21_X1 U4848 ( .B1(n5501), .B2(n5500), .A(n5499), .ZN(n5505) );
  NAND2_X1 U4849 ( .A1(n5503), .A2(n5502), .ZN(n5504) );
  XOR2_X1 U4850 ( .A(n5505), .B(n5504), .Z(n5506) );
  AOI22_X1 U4851 ( .A1(n5506), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[13]), 
        .ZN(n5509) );
  NAND2_X1 U4852 ( .A1(n5507), .A2(n5540), .ZN(n5508) );
  OAI211_X1 U4853 ( .C1(n5510), .C2(n6095), .A(n5509), .B(n5508), .ZN(n5511)
         );
  AOI21_X1 U4854 ( .B1(n5512), .B2(n5529), .A(n5511), .ZN(n5513) );
  NAND2_X1 U4855 ( .A1(n5514), .A2(n5513), .ZN(n5517) );
  OAI22_X1 U4856 ( .A1(n4894), .A2(n5543), .B1(n5794), .B2(n5515), .ZN(n5516)
         );
  NOR3_X1 U4857 ( .A1(n5517), .A2(n5516), .A3(n5523), .ZN(n5518) );
  OAI21_X1 U4858 ( .B1(n5800), .B2(n5894), .A(n5518), .ZN(result_o[13]) );
  AOI222_X1 U4859 ( .A1(n5522), .A2(clpx_shift_i[1]), .B1(n5521), .B2(n5797), 
        .C1(n5520), .C2(n5519), .ZN(n5901) );
  AOI21_X1 U4860 ( .B1(n5524), .B2(n5897), .A(n5523), .ZN(n5548) );
  NAND2_X1 U4861 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  XNOR2_X1 U4862 ( .A(n5528), .B(n5527), .ZN(n5546) );
  NAND2_X1 U4863 ( .A1(n5530), .A2(n5529), .ZN(n5542) );
  NAND2_X1 U4864 ( .A1(n5532), .A2(n5531), .ZN(n5533) );
  XOR2_X1 U4865 ( .A(n5534), .B(n5533), .Z(n5535) );
  AOI22_X1 U4866 ( .A1(n5535), .A2(n5796), .B1(n5605), .B2(dot_op_c_i[14]), 
        .ZN(n5536) );
  OAI21_X1 U4867 ( .B1(n5537), .B2(n6095), .A(n5536), .ZN(n5538) );
  AOI21_X1 U4868 ( .B1(n5540), .B2(n5539), .A(n5538), .ZN(n5541) );
  OAI211_X1 U4869 ( .C1(n5544), .C2(n5543), .A(n5542), .B(n5541), .ZN(n5545)
         );
  AOI21_X1 U4870 ( .B1(n5546), .B2(n5615), .A(n5545), .ZN(n5547) );
  OAI211_X1 U4871 ( .C1(n5901), .C2(n5894), .A(n5548), .B(n5547), .ZN(
        result_o[14]) );
  AOI22_X1 U4872 ( .A1(n5549), .A2(n5796), .B1(n38), .B2(dot_op_c_i[16]), .ZN(
        n5550) );
  OAI21_X1 U4873 ( .B1(n5551), .B2(n6095), .A(n5550), .ZN(n5557) );
  INV_X1 U4874 ( .A(n5552), .ZN(n5555) );
  AOI211_X1 U4875 ( .C1(n5555), .C2(n5554), .A(n5553), .B(n2829), .ZN(n5556)
         );
  AOI211_X1 U4876 ( .C1(n5605), .C2(n5558), .A(n5557), .B(n5556), .ZN(n5565)
         );
  NAND2_X1 U4877 ( .A1(n5560), .A2(n5559), .ZN(n5561) );
  XNOR2_X1 U4878 ( .A(n5562), .B(n5561), .ZN(n5563) );
  NAND2_X1 U4879 ( .A1(n5563), .A2(n5615), .ZN(n5564) );
  OAI211_X1 U4880 ( .C1(n5566), .C2(n5703), .A(n5565), .B(n5564), .ZN(
        result_o[16]) );
  OAI21_X1 U4881 ( .B1(n5583), .B2(n5568), .A(n5567), .ZN(n5572) );
  NAND2_X1 U4882 ( .A1(n5570), .A2(n5569), .ZN(n5571) );
  XNOR2_X1 U4883 ( .A(n5572), .B(n5571), .ZN(n5577) );
  AOI22_X1 U4884 ( .A1(n5573), .A2(n5796), .B1(n38), .B2(dot_op_c_i[21]), .ZN(
        n5574) );
  OAI21_X1 U4885 ( .B1(n5575), .B2(n6106), .A(n5574), .ZN(n5576) );
  AOI21_X1 U4886 ( .B1(n5577), .B2(n5615), .A(n5576), .ZN(n5580) );
  NAND2_X1 U4887 ( .A1(n5701), .A2(n5703), .ZN(n5603) );
  OAI21_X1 U4888 ( .B1(n5578), .B2(n5620), .A(n5603), .ZN(n5579) );
  NAND2_X1 U4889 ( .A1(n5580), .A2(n5579), .ZN(result_o[21]) );
  OAI21_X1 U4890 ( .B1(n5583), .B2(n5582), .A(n5581), .ZN(n5596) );
  NAND2_X1 U4891 ( .A1(n5595), .A2(n5584), .ZN(n5585) );
  XNOR2_X1 U4892 ( .A(n5596), .B(n5585), .ZN(n5586) );
  NAND2_X1 U4893 ( .A1(n5586), .A2(n5615), .ZN(n5593) );
  OAI21_X1 U4894 ( .B1(n5587), .B2(n5620), .A(n5603), .ZN(n5592) );
  AOI22_X1 U4895 ( .A1(n5588), .A2(n5796), .B1(n38), .B2(dot_op_c_i[22]), .ZN(
        n5591) );
  NAND2_X1 U4896 ( .A1(n5589), .A2(n5605), .ZN(n5590) );
  NAND4_X1 U4897 ( .A1(n5593), .A2(n5592), .A3(n5591), .A4(n5590), .ZN(
        result_o[22]) );
  AOI21_X1 U4898 ( .B1(n5596), .B2(n5595), .A(n5594), .ZN(n5600) );
  NAND2_X1 U4899 ( .A1(n5598), .A2(n5597), .ZN(n5599) );
  XOR2_X1 U4900 ( .A(n5600), .B(n5599), .Z(n5601) );
  NAND2_X1 U4901 ( .A1(n5601), .A2(n5615), .ZN(n5610) );
  AOI22_X1 U4902 ( .A1(n5602), .A2(n5796), .B1(n38), .B2(dot_op_c_i[23]), .ZN(
        n5609) );
  OAI21_X1 U4903 ( .B1(n5604), .B2(n5620), .A(n5603), .ZN(n5608) );
  NAND2_X1 U4904 ( .A1(n5606), .A2(n5605), .ZN(n5607) );
  NAND4_X1 U4905 ( .A1(n5610), .A2(n5609), .A3(n5608), .A4(n5607), .ZN(
        result_o[23]) );
  NAND2_X1 U4906 ( .A1(n5612), .A2(n5611), .ZN(n5613) );
  XNOR2_X1 U4907 ( .A(n5614), .B(n5613), .ZN(n5616) );
  NAND2_X1 U4908 ( .A1(n5616), .A2(n5615), .ZN(n5624) );
  OAI22_X1 U4909 ( .A1(n5618), .A2(n6101), .B1(n5894), .B2(n5617), .ZN(n5619)
         );
  AOI211_X1 U4910 ( .C1(n5622), .C2(n5621), .A(n5620), .B(n5619), .ZN(n5623)
         );
  OAI211_X1 U4911 ( .C1(n5625), .C2(n6106), .A(n5624), .B(n5623), .ZN(
        result_o[24]) );
  OAI21_X1 U4912 ( .B1(n5626), .B2(n5709), .A(n5712), .ZN(n5697) );
  FA_X1 U4913 ( .A(n5629), .B(n5628), .CI(n5627), .CO(n5788), .S(n5690) );
  FA_X1 U4914 ( .A(n5632), .B(n5631), .CI(n5630), .CO(n5784), .S(n5686) );
  XNOR2_X1 U4915 ( .A(n6121), .B(op_b_i[17]), .ZN(n5730) );
  OAI22_X1 U4916 ( .A1(n5633), .A2(n5915), .B1(n5730), .B2(n5917), .ZN(n5753)
         );
  XNOR2_X1 U4917 ( .A(n5844), .B(n4123), .ZN(n5733) );
  OAI22_X1 U4918 ( .A1(n5634), .A2(n5925), .B1(n5733), .B2(n5927), .ZN(n5752)
         );
  XNOR2_X1 U4919 ( .A(n6118), .B(op_a_i[28]), .ZN(n5812) );
  XNOR2_X1 U4920 ( .A(n5812), .B(n5856), .ZN(n5727) );
  OAI22_X1 U4921 ( .A1(n5636), .A2(n3241), .B1(n5727), .B2(n5635), .ZN(n5751)
         );
  XNOR2_X1 U4922 ( .A(n52), .B(op_b_i[19]), .ZN(n5766) );
  OAI22_X1 U4923 ( .A1(n5637), .A2(n6032), .B1(n5766), .B2(n6034), .ZN(n5747)
         );
  XNOR2_X1 U4924 ( .A(n19), .B(op_b_i[23]), .ZN(n5760) );
  OAI22_X1 U4925 ( .A1(n5638), .A2(n5981), .B1(n5760), .B2(n5983), .ZN(n5746)
         );
  XNOR2_X1 U4926 ( .A(n55), .B(op_b_i[25]), .ZN(n5767) );
  OAI22_X1 U4927 ( .A1(n5639), .A2(n5993), .B1(n5767), .B2(n5995), .ZN(n5745)
         );
  XNOR2_X1 U4928 ( .A(n5867), .B(n27), .ZN(n5765) );
  OAI22_X1 U4929 ( .A1(n5640), .A2(n5822), .B1(n5765), .B2(n4546), .ZN(n5756)
         );
  XNOR2_X1 U4930 ( .A(n5814), .B(n5807), .ZN(n5728) );
  OAI22_X1 U4931 ( .A1(n5641), .A2(n2867), .B1(n5728), .B2(n5809), .ZN(n5755)
         );
  XNOR2_X1 U4932 ( .A(n5821), .B(n5919), .ZN(n5734) );
  OAI22_X1 U4933 ( .A1(n5642), .A2(n3128), .B1(n5734), .B2(n5922), .ZN(n5754)
         );
  FA_X1 U4934 ( .A(n5645), .B(n5644), .CI(n5643), .CO(n5775), .S(n5631) );
  FA_X1 U4935 ( .A(n5648), .B(n5647), .CI(n5646), .CO(n5774), .S(n5632) );
  FA_X1 U4936 ( .A(n5651), .B(n5650), .CI(n5649), .CO(n5741), .S(n5680) );
  FA_X1 U4937 ( .A(n5654), .B(n5653), .CI(n5652), .CO(n5770), .S(n5649) );
  HA_X1 U4938 ( .A(n5656), .B(n5655), .CO(n5769), .S(n5671) );
  FA_X1 U4939 ( .A(n5659), .B(n5658), .CI(n5657), .CO(n5768), .S(n5651) );
  FA_X1 U4940 ( .A(n5662), .B(n5661), .CI(n5660), .CO(n5773), .S(n5645) );
  FA_X1 U4941 ( .A(n5665), .B(n5664), .CI(n5663), .CO(n5772), .S(n5644) );
  XNOR2_X1 U4942 ( .A(n5848), .B(op_b_i[27]), .ZN(n5729) );
  OAI22_X1 U4943 ( .A1(n5666), .A2(n6036), .B1(n5729), .B2(n6038), .ZN(n5750)
         );
  XNOR2_X1 U4944 ( .A(op_b_i[27]), .B(op_b_i[28]), .ZN(n5979) );
  INV_X1 U4945 ( .A(n5979), .ZN(n5667) );
  AND2_X1 U4946 ( .A1(n6116), .A2(n5667), .ZN(n5749) );
  XNOR2_X1 U4947 ( .A(n20), .B(op_b_i[21]), .ZN(n5761) );
  OAI22_X1 U4948 ( .A1(n5668), .A2(n5997), .B1(n5761), .B2(n68), .ZN(n5748) );
  FA_X1 U4949 ( .A(n5671), .B(n5670), .CI(n5669), .CO(n5738), .S(n5647) );
  XNOR2_X1 U4950 ( .A(n5819), .B(op_b_i[13]), .ZN(n5735) );
  OAI22_X1 U4951 ( .A1(n5672), .A2(n5934), .B1(n5735), .B2(n72), .ZN(n5759) );
  XNOR2_X1 U4952 ( .A(n5808), .B(n5811), .ZN(n5726) );
  OAI22_X1 U4953 ( .A1(n5673), .A2(n2585), .B1(n5726), .B2(n10), .ZN(n5758) );
  XNOR2_X1 U4954 ( .A(n5824), .B(n5941), .ZN(n5764) );
  OAI22_X1 U4955 ( .A1(n5674), .A2(n5943), .B1(n5764), .B2(n26), .ZN(n5757) );
  FA_X1 U4956 ( .A(n5677), .B(n5676), .CI(n5675), .CO(n5736), .S(n5646) );
  FA_X1 U4957 ( .A(n5680), .B(n5679), .CI(n5678), .CO(n5723), .S(n5687) );
  AND2_X1 U4958 ( .A1(n5681), .A2(n29), .ZN(n5787) );
  INV_X1 U4959 ( .A(op_b_i[28]), .ZN(n5682) );
  NOR2_X1 U4960 ( .A1(n6118), .A2(n5682), .ZN(n5683) );
  OR2_X1 U4961 ( .A1(n5683), .A2(n6145), .ZN(n5781) );
  OAI22_X1 U4962 ( .A1(n6146), .A2(n5699), .B1(n2525), .B2(n914), .ZN(n5780)
         );
  HA_X1 U4963 ( .A(n5685), .B(n5684), .CO(n5721), .S(n5629) );
  FA_X1 U4964 ( .A(n5688), .B(n5687), .CI(n5686), .CO(n5689), .S(n4556) );
  OR2_X1 U4965 ( .A1(n5689), .A2(n6145), .ZN(n5720) );
  FA_X1 U4966 ( .A(n5692), .B(n5691), .CI(n5690), .CO(n5693), .S(n4569) );
  NOR2_X1 U4967 ( .A1(n5694), .A2(n5693), .ZN(n5713) );
  INV_X1 U4968 ( .A(n5713), .ZN(n5695) );
  NAND2_X1 U4969 ( .A1(n5694), .A2(n5693), .ZN(n5711) );
  NAND2_X1 U4970 ( .A1(n5695), .A2(n5711), .ZN(n5696) );
  XNOR2_X1 U4971 ( .A(n5697), .B(n5696), .ZN(n5698) );
  NAND2_X1 U4972 ( .A1(n5698), .A2(n5615), .ZN(n5707) );
  OAI22_X1 U4973 ( .A1(n5700), .A2(n6095), .B1(n5894), .B2(n5699), .ZN(n5704)
         );
  OAI21_X1 U4974 ( .B1(n5703), .B2(n5702), .A(n5701), .ZN(n6099) );
  AOI211_X1 U4975 ( .C1(n5705), .C2(n5796), .A(n5704), .B(n6099), .ZN(n5706)
         );
  OAI211_X1 U4976 ( .C1(n5708), .C2(n6106), .A(n5707), .B(n5706), .ZN(
        result_o[28]) );
  NOR2_X1 U4977 ( .A1(n5709), .A2(n5713), .ZN(n5716) );
  NAND2_X1 U4978 ( .A1(n5716), .A2(n5710), .ZN(n5719) );
  OAI21_X1 U4979 ( .B1(n5713), .B2(n5712), .A(n5711), .ZN(n5714) );
  AOI21_X1 U4980 ( .B1(n5716), .B2(n5715), .A(n5714), .ZN(n5717) );
  OAI21_X1 U4981 ( .B1(n5719), .B2(n5718), .A(n5717), .ZN(n5890) );
  FA_X1 U4982 ( .A(n5722), .B(n5721), .CI(n5720), .CO(n5886), .S(n5786) );
  FA_X1 U4983 ( .A(n5725), .B(n5724), .CI(n5723), .CO(n5882), .S(n5782) );
  XNOR2_X1 U4984 ( .A(n6008), .B(n5811), .ZN(n5813) );
  OAI22_X1 U4985 ( .A1(n5813), .A2(n10), .B1(n5726), .B2(n2585), .ZN(n5834) );
  XNOR2_X1 U4986 ( .A(n6119), .B(op_a_i[29]), .ZN(n6016) );
  XNOR2_X1 U4987 ( .A(n6016), .B(n5856), .ZN(n5858) );
  OAI22_X1 U4988 ( .A1(n5858), .A2(n5635), .B1(n5727), .B2(n3241), .ZN(n5833)
         );
  XNOR2_X1 U4989 ( .A(n5920), .B(n5807), .ZN(n5810) );
  OAI22_X1 U4990 ( .A1(n5810), .A2(n5809), .B1(n5728), .B2(n2867), .ZN(n5832)
         );
  XNOR2_X1 U4991 ( .A(n56), .B(op_b_i[27]), .ZN(n5846) );
  OAI22_X1 U4992 ( .A1(n5846), .A2(n6038), .B1(n5729), .B2(n6036), .ZN(n5871)
         );
  XNOR2_X1 U4993 ( .A(n66), .B(op_b_i[17]), .ZN(n5845) );
  OAI22_X1 U4994 ( .A1(n5845), .A2(n5917), .B1(n5730), .B2(n5915), .ZN(n5870)
         );
  XNOR2_X1 U4995 ( .A(n6116), .B(op_b_i[29]), .ZN(n5732) );
  XOR2_X1 U4996 ( .A(op_b_i[28]), .B(op_b_i[29]), .Z(n5731) );
  NAND2_X1 U4997 ( .A1(n5731), .A2(n5979), .ZN(n5977) );
  XNOR2_X1 U4998 ( .A(n6002), .B(op_b_i[29]), .ZN(n5849) );
  OAI22_X1 U4999 ( .A1(n5732), .A2(n5977), .B1(n5849), .B2(n5979), .ZN(n5869)
         );
  XNOR2_X1 U5000 ( .A(n5914), .B(n4123), .ZN(n5820) );
  OAI22_X1 U5001 ( .A1(n5820), .A2(n5927), .B1(n5733), .B2(n5925), .ZN(n5840)
         );
  XNOR2_X1 U5002 ( .A(n5938), .B(n5919), .ZN(n5815) );
  OAI22_X1 U5003 ( .A1(n5815), .A2(n5922), .B1(n5734), .B2(n3128), .ZN(n5839)
         );
  XNOR2_X1 U5004 ( .A(n5924), .B(op_b_i[13]), .ZN(n5825) );
  OAI22_X1 U5005 ( .A1(n5825), .A2(n72), .B1(n5735), .B2(n5934), .ZN(n5838) );
  FA_X1 U5006 ( .A(n5738), .B(n5737), .CI(n5736), .CO(n5873), .S(n5724) );
  FA_X1 U5007 ( .A(n5741), .B(n5740), .CI(n5739), .CO(n5872), .S(n5725) );
  FA_X1 U5008 ( .A(n5744), .B(n5743), .CI(n5742), .CO(n5831), .S(n5776) );
  FA_X1 U5009 ( .A(n5747), .B(n5746), .CI(n5745), .CO(n5864), .S(n5743) );
  FA_X1 U5010 ( .A(n5750), .B(n5749), .CI(n5748), .CO(n5863), .S(n5771) );
  FA_X1 U5011 ( .A(n5753), .B(n5752), .CI(n5751), .CO(n5862), .S(n5744) );
  FA_X1 U5012 ( .A(n5756), .B(n5755), .CI(n5754), .CO(n5861), .S(n5742) );
  FA_X1 U5013 ( .A(n5759), .B(n5758), .CI(n5757), .CO(n5860), .S(n5737) );
  XNOR2_X1 U5014 ( .A(n54), .B(op_b_i[23]), .ZN(n5855) );
  OAI22_X1 U5015 ( .A1(n5855), .A2(n5983), .B1(n5760), .B2(n5981), .ZN(n5837)
         );
  XNOR2_X1 U5016 ( .A(n21), .B(op_b_i[21]), .ZN(n5847) );
  OAI22_X1 U5017 ( .A1(n5847), .A2(n68), .B1(n5761), .B2(n5997), .ZN(n5836) );
  INV_X1 U5018 ( .A(op_b_i[29]), .ZN(n5762) );
  OR2_X1 U5019 ( .A1(n6116), .A2(n5762), .ZN(n5763) );
  OAI22_X1 U5020 ( .A1(n5763), .A2(n5979), .B1(n5977), .B2(n5762), .ZN(n5835)
         );
  XNOR2_X1 U5021 ( .A(n5933), .B(n5941), .ZN(n5868) );
  OAI22_X1 U5022 ( .A1(n5868), .A2(n26), .B1(n5764), .B2(n5943), .ZN(n5818) );
  XNOR2_X1 U5023 ( .A(n5942), .B(n27), .ZN(n5823) );
  OAI22_X1 U5024 ( .A1(n5823), .A2(n2871), .B1(n5765), .B2(n5822), .ZN(n5817)
         );
  XNOR2_X1 U5025 ( .A(n51), .B(op_b_i[19]), .ZN(n5854) );
  OAI22_X1 U5026 ( .A1(n5854), .A2(n6034), .B1(n5766), .B2(n6032), .ZN(n5866)
         );
  XNOR2_X1 U5027 ( .A(n22), .B(op_b_i[25]), .ZN(n5852) );
  OAI22_X1 U5028 ( .A1(n5852), .A2(n5995), .B1(n5767), .B2(n5993), .ZN(n5865)
         );
  FA_X1 U5029 ( .A(n5770), .B(n5769), .CI(n5768), .CO(n5827), .S(n5740) );
  FA_X1 U5030 ( .A(n5773), .B(n5772), .CI(n5771), .CO(n5826), .S(n5739) );
  FA_X1 U5031 ( .A(n5776), .B(n5775), .CI(n5774), .CO(n5804), .S(n5783) );
  AND2_X1 U5032 ( .A1(n5777), .A2(n29), .ZN(n5885) );
  NOR2_X1 U5033 ( .A1(n6118), .A2(n5762), .ZN(n5778) );
  OR2_X1 U5034 ( .A1(n5778), .A2(n6145), .ZN(n5879) );
  INV_X1 U5035 ( .A(op_c_i[29]), .ZN(n5779) );
  OAI22_X1 U5036 ( .A1(n6146), .A2(n5793), .B1(n2525), .B2(n5779), .ZN(n5878)
         );
  HA_X1 U5037 ( .A(n5781), .B(n5780), .CO(n5802), .S(n5722) );
  FA_X1 U5038 ( .A(n5784), .B(n5783), .CI(n5782), .CO(n5785), .S(n5681) );
  OR2_X1 U5039 ( .A1(n5785), .A2(n6145), .ZN(n5801) );
  FA_X1 U5040 ( .A(n5788), .B(n5787), .CI(n5786), .CO(n5789), .S(n5694) );
  OR2_X1 U5041 ( .A1(n5790), .A2(n5789), .ZN(n5889) );
  NAND2_X1 U5042 ( .A1(n5790), .A2(n5789), .ZN(n5887) );
  NAND2_X1 U5043 ( .A1(n5889), .A2(n5887), .ZN(n5791) );
  XNOR2_X1 U5044 ( .A(n5890), .B(n5791), .ZN(n5792) );
  NAND2_X1 U5045 ( .A1(n5792), .A2(n5615), .ZN(n5799) );
  OAI22_X1 U5046 ( .A1(n5794), .A2(n6095), .B1(n5894), .B2(n5793), .ZN(n5795)
         );
  AOI211_X1 U5047 ( .C1(n5797), .C2(n5796), .A(n5795), .B(n6099), .ZN(n5798)
         );
  OAI211_X1 U5048 ( .C1(n5800), .C2(n6106), .A(n5799), .B(n5798), .ZN(
        result_o[29]) );
  FA_X1 U5049 ( .A(n5803), .B(n5802), .CI(n5801), .CO(n5907), .S(n5884) );
  FA_X1 U5050 ( .A(n5806), .B(n5805), .CI(n5804), .CO(n6071), .S(n5880) );
  XNOR2_X1 U5051 ( .A(n5808), .B(n5807), .ZN(n6009) );
  OAI22_X1 U5052 ( .A1(n5810), .A2(n2867), .B1(n6009), .B2(n5809), .ZN(n5963)
         );
  XNOR2_X1 U5053 ( .A(n5812), .B(n5811), .ZN(n6017) );
  OAI22_X1 U5054 ( .A1(n5813), .A2(n2585), .B1(n6017), .B2(n10), .ZN(n5962) );
  XNOR2_X1 U5055 ( .A(n5814), .B(n5919), .ZN(n5921) );
  OAI22_X1 U5056 ( .A1(n5815), .A2(n3128), .B1(n5921), .B2(n5922), .ZN(n5961)
         );
  FA_X1 U5057 ( .A(n5818), .B(n5817), .CI(n5816), .CO(n5974), .S(n5828) );
  XNOR2_X1 U5058 ( .A(n5819), .B(op_b_i[15]), .ZN(n5926) );
  OAI22_X1 U5059 ( .A1(n5820), .A2(n5925), .B1(n5926), .B2(n5927), .ZN(n5969)
         );
  XNOR2_X1 U5060 ( .A(n5821), .B(n27), .ZN(n5939) );
  OAI22_X1 U5061 ( .A1(n5823), .A2(n5822), .B1(n5939), .B2(n4546), .ZN(n5968)
         );
  XNOR2_X1 U5062 ( .A(n5824), .B(op_b_i[13]), .ZN(n5935) );
  OAI22_X1 U5063 ( .A1(n5825), .A2(n5934), .B1(n5935), .B2(n72), .ZN(n5967) );
  FA_X1 U5064 ( .A(n5828), .B(n5827), .CI(n5826), .CO(n6058), .S(n5805) );
  FA_X1 U5065 ( .A(n5831), .B(n5830), .CI(n5829), .CO(n6057), .S(n5806) );
  FA_X1 U5066 ( .A(n5834), .B(n5833), .CI(n5832), .CO(n6050), .S(n5843) );
  FA_X1 U5067 ( .A(n5837), .B(n5836), .CI(n5835), .CO(n6049), .S(n5859) );
  FA_X1 U5068 ( .A(n5840), .B(n5839), .CI(n5838), .CO(n6048), .S(n5841) );
  FA_X1 U5069 ( .A(n5843), .B(n5842), .CI(n5841), .CO(n5956), .S(n5874) );
  XNOR2_X1 U5070 ( .A(n5844), .B(op_b_i[17]), .ZN(n5916) );
  OAI22_X1 U5071 ( .A1(n5845), .A2(n5915), .B1(n5916), .B2(n5917), .ZN(n6044)
         );
  XNOR2_X1 U5072 ( .A(n55), .B(op_b_i[27]), .ZN(n6037) );
  OAI22_X1 U5073 ( .A1(n5846), .A2(n6036), .B1(n6037), .B2(n6038), .ZN(n6043)
         );
  XNOR2_X1 U5074 ( .A(n52), .B(op_b_i[21]), .ZN(n5998) );
  OAI22_X1 U5075 ( .A1(n5847), .A2(n5997), .B1(n5998), .B2(n68), .ZN(n6042) );
  XNOR2_X1 U5076 ( .A(n5848), .B(op_b_i[29]), .ZN(n5978) );
  OAI22_X1 U5077 ( .A1(n5849), .A2(n5977), .B1(n5978), .B2(n5979), .ZN(n6030)
         );
  XNOR2_X1 U5078 ( .A(op_b_i[29]), .B(op_b_i[30]), .ZN(n6013) );
  INV_X1 U5079 ( .A(n6013), .ZN(n5850) );
  AND2_X1 U5080 ( .A1(n6116), .A2(n5850), .ZN(n6029) );
  XNOR2_X1 U5081 ( .A(n19), .B(op_b_i[25]), .ZN(n5994) );
  OAI22_X1 U5082 ( .A1(n5852), .A2(n5993), .B1(n5994), .B2(n5995), .ZN(n6028)
         );
  XNOR2_X1 U5083 ( .A(n6120), .B(op_b_i[19]), .ZN(n6033) );
  OAI22_X1 U5084 ( .A1(n5854), .A2(n6032), .B1(n6033), .B2(n6034), .ZN(n5966)
         );
  XNOR2_X1 U5085 ( .A(n20), .B(op_b_i[23]), .ZN(n5982) );
  OAI22_X1 U5086 ( .A1(n5855), .A2(n5981), .B1(n5982), .B2(n5983), .ZN(n5965)
         );
  XNOR2_X1 U5087 ( .A(n6119), .B(op_a_i[30]), .ZN(n5857) );
  XNOR2_X1 U5088 ( .A(n5857), .B(n5856), .ZN(n5987) );
  OAI22_X1 U5089 ( .A1(n5858), .A2(n3241), .B1(n5987), .B2(n5635), .ZN(n5964)
         );
  FA_X1 U5090 ( .A(n5861), .B(n5860), .CI(n5859), .CO(n5913), .S(n5829) );
  FA_X1 U5091 ( .A(n5864), .B(n5863), .CI(n5862), .CO(n5912), .S(n5830) );
  HA_X1 U5092 ( .A(n5866), .B(n5865), .CO(n5951), .S(n5816) );
  XNOR2_X1 U5093 ( .A(n5867), .B(op_b_i[11]), .ZN(n5944) );
  OAI22_X1 U5094 ( .A1(n5868), .A2(n5943), .B1(n5944), .B2(n26), .ZN(n5950) );
  FA_X1 U5095 ( .A(n5871), .B(n5870), .CI(n5869), .CO(n5949), .S(n5842) );
  FA_X1 U5096 ( .A(n5874), .B(n5873), .CI(n5872), .CO(n5908), .S(n5881) );
  AND2_X1 U5097 ( .A1(n5875), .A2(n29), .ZN(n5906) );
  INV_X1 U5098 ( .A(op_b_i[30]), .ZN(n5876) );
  NOR2_X1 U5099 ( .A1(n6118), .A2(n5876), .ZN(n5877) );
  OR2_X1 U5100 ( .A1(n5877), .A2(n6145), .ZN(n6068) );
  OAI22_X1 U5101 ( .A1(n6146), .A2(n5893), .B1(n2525), .B2(n988), .ZN(n6067)
         );
  HA_X1 U5102 ( .A(n5879), .B(n5878), .CO(n6084), .S(n5803) );
  FA_X1 U5103 ( .A(n5882), .B(n5881), .CI(n5880), .CO(n5883), .S(n5777) );
  OR2_X1 U5104 ( .A1(n5883), .A2(n6144), .ZN(n6083) );
  FA_X1 U5105 ( .A(n5886), .B(n5885), .CI(n5884), .CO(n5903), .S(n5790) );
  INV_X1 U5106 ( .A(n5887), .ZN(n5888) );
  AOI21_X1 U5107 ( .B1(n5890), .B2(n5889), .A(n5888), .ZN(n5891) );
  INV_X1 U5108 ( .A(n5891), .ZN(n5902) );
  NAND2_X1 U5109 ( .A1(n5892), .A2(n5615), .ZN(n5900) );
  OAI22_X1 U5110 ( .A1(n5895), .A2(n6101), .B1(n5894), .B2(n5893), .ZN(n5896)
         );
  AOI211_X1 U5111 ( .C1(n5898), .C2(n5897), .A(n6099), .B(n5896), .ZN(n5899)
         );
  OAI211_X1 U5112 ( .C1(n5901), .C2(n6106), .A(n5900), .B(n5899), .ZN(
        result_o[30]) );
  FA_X1 U5113 ( .A(n5904), .B(n5903), .CI(n5902), .CO(n6093), .S(n5892) );
  FA_X1 U5114 ( .A(n5907), .B(n5906), .CI(n5905), .CO(n6091), .S(n5904) );
  FA_X1 U5115 ( .A(n5910), .B(n5909), .CI(n5908), .CO(n6065), .S(n6069) );
  FA_X1 U5116 ( .A(n5913), .B(n5912), .CI(n5911), .CO(n5960), .S(n5909) );
  XNOR2_X1 U5117 ( .A(n5914), .B(op_b_i[17]), .ZN(n5918) );
  OAI22_X1 U5118 ( .A1(n5918), .A2(n5917), .B1(n5916), .B2(n5915), .ZN(n5931)
         );
  XNOR2_X1 U5119 ( .A(n5920), .B(n5919), .ZN(n5923) );
  OAI22_X1 U5120 ( .A1(n5923), .A2(n5922), .B1(n5921), .B2(n3128), .ZN(n5930)
         );
  XNOR2_X1 U5121 ( .A(n5924), .B(op_b_i[15]), .ZN(n5928) );
  OAI22_X1 U5122 ( .A1(n5928), .A2(n5927), .B1(n5926), .B2(n5925), .ZN(n5929)
         );
  FA_X1 U5123 ( .A(n5931), .B(n5930), .CI(n5929), .S(n5954) );
  XNOR2_X1 U5124 ( .A(n5933), .B(op_b_i[13]), .ZN(n5937) );
  OAI22_X1 U5125 ( .A1(n5937), .A2(n72), .B1(n5935), .B2(n5934), .ZN(n5948) );
  XNOR2_X1 U5126 ( .A(n5938), .B(n27), .ZN(n5940) );
  OAI22_X1 U5127 ( .A1(n5940), .A2(n2871), .B1(n5939), .B2(n5822), .ZN(n5947)
         );
  XNOR2_X1 U5128 ( .A(n5942), .B(n5941), .ZN(n5945) );
  OAI22_X1 U5129 ( .A1(n5945), .A2(n26), .B1(n5944), .B2(n5943), .ZN(n5946) );
  FA_X1 U5130 ( .A(n5948), .B(n5947), .CI(n5946), .S(n5953) );
  FA_X1 U5131 ( .A(n5951), .B(n5950), .CI(n5949), .CO(n5952), .S(n5911) );
  FA_X1 U5132 ( .A(n5954), .B(n5953), .CI(n5952), .S(n5959) );
  FA_X1 U5133 ( .A(n5957), .B(n5956), .CI(n5955), .CO(n5958), .S(n5910) );
  FA_X1 U5134 ( .A(n5960), .B(n5959), .CI(n5958), .S(n6064) );
  FA_X1 U5135 ( .A(n5963), .B(n5962), .CI(n5961), .CO(n5972), .S(n5975) );
  FA_X1 U5136 ( .A(n5966), .B(n5965), .CI(n5964), .CO(n5971), .S(n6051) );
  FA_X1 U5137 ( .A(n5969), .B(n5968), .CI(n5967), .CO(n5970), .S(n5973) );
  FA_X1 U5138 ( .A(n5972), .B(n5971), .CI(n5970), .S(n6027) );
  FA_X1 U5139 ( .A(n5975), .B(n5974), .CI(n5973), .CO(n6026), .S(n6059) );
  XNOR2_X1 U5140 ( .A(n56), .B(op_b_i[29]), .ZN(n5980) );
  OAI22_X1 U5141 ( .A1(n5980), .A2(n5979), .B1(n5978), .B2(n5977), .ZN(n5991)
         );
  XNOR2_X1 U5142 ( .A(n21), .B(op_b_i[23]), .ZN(n5984) );
  OAI22_X1 U5143 ( .A1(n5984), .A2(n5983), .B1(n5982), .B2(n5981), .ZN(n5990)
         );
  XNOR2_X1 U5144 ( .A(n6119), .B(op_a_i[31]), .ZN(n5986) );
  XNOR2_X1 U5145 ( .A(n5986), .B(n5985), .ZN(n5988) );
  OAI22_X1 U5146 ( .A1(n5988), .A2(n5635), .B1(n5987), .B2(n3241), .ZN(n5989)
         );
  FA_X1 U5147 ( .A(n5991), .B(n5990), .CI(n5989), .S(n6024) );
  XNOR2_X1 U5148 ( .A(n54), .B(op_b_i[25]), .ZN(n5996) );
  OAI22_X1 U5149 ( .A1(n5996), .A2(n5995), .B1(n5994), .B2(n5993), .ZN(n6007)
         );
  XNOR2_X1 U5150 ( .A(n51), .B(op_b_i[21]), .ZN(n6000) );
  OAI22_X1 U5151 ( .A1(n6000), .A2(n68), .B1(n5998), .B2(n5997), .ZN(n6006) );
  XNOR2_X1 U5152 ( .A(n6116), .B(op_b_i[31]), .ZN(n6004) );
  XOR2_X1 U5153 ( .A(op_b_i[30]), .B(op_b_i[31]), .Z(n6001) );
  NAND2_X1 U5154 ( .A1(n6001), .A2(n6013), .ZN(n6012) );
  XNOR2_X1 U5155 ( .A(n6002), .B(op_b_i[31]), .ZN(n6003) );
  OAI22_X1 U5156 ( .A1(n6004), .A2(n6012), .B1(n6003), .B2(n6013), .ZN(n6005)
         );
  FA_X1 U5157 ( .A(n6007), .B(n6006), .CI(n6005), .S(n6023) );
  XNOR2_X1 U5158 ( .A(n6008), .B(n25), .ZN(n6011) );
  OAI22_X1 U5159 ( .A1(n6011), .A2(n6010), .B1(n6009), .B2(n2867), .ZN(n6021)
         );
  OR2_X1 U5160 ( .A1(n6116), .A2(n6073), .ZN(n6014) );
  OAI22_X1 U5161 ( .A1(n6014), .A2(n6013), .B1(n6012), .B2(n6073), .ZN(n6020)
         );
  XNOR2_X1 U5162 ( .A(n6016), .B(n6015), .ZN(n6018) );
  OAI22_X1 U5163 ( .A1(n6018), .A2(n10), .B1(n6017), .B2(n2585), .ZN(n6019) );
  FA_X1 U5164 ( .A(n6021), .B(n6020), .CI(n6019), .S(n6022) );
  FA_X1 U5165 ( .A(n6024), .B(n6023), .CI(n6022), .S(n6025) );
  FA_X1 U5166 ( .A(n6027), .B(n6026), .CI(n6025), .S(n6062) );
  FA_X1 U5167 ( .A(n6030), .B(n6029), .CI(n6028), .CO(n6047), .S(n6052) );
  XNOR2_X1 U5168 ( .A(n65), .B(op_b_i[19]), .ZN(n6035) );
  OAI22_X1 U5169 ( .A1(n6035), .A2(n6034), .B1(n6033), .B2(n6032), .ZN(n6041)
         );
  XNOR2_X1 U5170 ( .A(n22), .B(op_b_i[27]), .ZN(n6039) );
  OAI22_X1 U5171 ( .A1(n6039), .A2(n6038), .B1(n6037), .B2(n6036), .ZN(n6040)
         );
  HA_X1 U5172 ( .A(n6041), .B(n6040), .S(n6046) );
  FA_X1 U5173 ( .A(n6044), .B(n6043), .CI(n6042), .CO(n6045), .S(n6053) );
  FA_X1 U5174 ( .A(n6047), .B(n6046), .CI(n6045), .S(n6056) );
  FA_X1 U5175 ( .A(n6050), .B(n6049), .CI(n6048), .CO(n6055), .S(n5957) );
  FA_X1 U5176 ( .A(n6053), .B(n6052), .CI(n6051), .CO(n6054), .S(n5955) );
  FA_X1 U5177 ( .A(n6056), .B(n6055), .CI(n6054), .S(n6061) );
  FA_X1 U5178 ( .A(n6059), .B(n6058), .CI(n6057), .CO(n6060), .S(n6070) );
  FA_X1 U5179 ( .A(n6062), .B(n6061), .CI(n6060), .S(n6063) );
  FA_X1 U5180 ( .A(n6065), .B(n6064), .CI(n6063), .S(n6066) );
  AND2_X1 U5181 ( .A1(n6066), .A2(n29), .ZN(n6089) );
  HA_X1 U5182 ( .A(n6068), .B(n6067), .CO(n6082), .S(n6085) );
  FA_X1 U5183 ( .A(n6071), .B(n6070), .CI(n6069), .CO(n6072), .S(n5875) );
  OR2_X1 U5184 ( .A1(n6072), .A2(n6144), .ZN(n6080) );
  NOR2_X1 U5185 ( .A1(n6119), .A2(n6073), .ZN(n6074) );
  OR2_X1 U5186 ( .A1(n6074), .A2(n6143), .ZN(n6078) );
  INV_X1 U5187 ( .A(op_c_i[31]), .ZN(n6075) );
  OAI22_X1 U5188 ( .A1(n6146), .A2(n6076), .B1(n2525), .B2(n6075), .ZN(n6077)
         );
  XOR2_X1 U5189 ( .A(n6078), .B(n6077), .Z(n6079) );
  XOR2_X1 U5190 ( .A(n6080), .B(n6079), .Z(n6081) );
  XOR2_X1 U5191 ( .A(n6082), .B(n6081), .Z(n6087) );
  FA_X1 U5192 ( .A(n6085), .B(n6084), .CI(n6083), .CO(n6086), .S(n5905) );
  XOR2_X1 U5193 ( .A(n6087), .B(n6086), .Z(n6088) );
  XOR2_X1 U5194 ( .A(n6089), .B(n6088), .Z(n6090) );
  XOR2_X1 U5195 ( .A(n6091), .B(n6090), .Z(n6092) );
  XOR2_X1 U5196 ( .A(n6093), .B(n6092), .Z(n6094) );
  NAND2_X1 U5197 ( .A1(n6094), .A2(n5615), .ZN(n6105) );
  OAI211_X1 U5198 ( .C1(n6107), .C2(n6106), .A(n6105), .B(n6104), .ZN(
        result_o[31]) );
  SDFFR_X1 mulh_CS_reg_0_ ( .D(n467), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(mulh_CS[0]), .QN(n6109) );
  SDFFR_X1 mulh_CS_reg_1_ ( .D(n465), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(mulh_CS[1]), .QN(n6110) );
  SDFFR_X1 mulh_CS_reg_2_ ( .D(n466), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(mulh_CS[2]), .QN(n6108) );
  SDFFR_X1 mulh_carry_q_reg ( .D(n464), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(mulh_carry_q) );
  OR2_X1 U111 ( .A1(mulh_CS[0]), .A2(mulh_CS[1]), .ZN(n109) );
  INV_X1 U114 ( .A(dot_op_a_i[0]), .ZN(n1777) );
  INV_X1 U14 ( .A(n3015), .ZN(n1785) );
  INV_X1 U97 ( .A(n1628), .ZN(n1612) );
  INV_X1 U101 ( .A(n3107), .ZN(n4123) );
  CLKBUF_X1 U60 ( .A(n3472), .Z(n62) );
  INV_X1 U15 ( .A(n3078), .ZN(n1808) );
  INV_X1 U10 ( .A(n1313), .ZN(n1307) );
  INV_X1 U12 ( .A(n3084), .ZN(n4679) );
  INV_X1 U9 ( .A(n2848), .ZN(n1803) );
  CLKBUF_X1 U58 ( .A(n3719), .Z(n59) );
  BUF_X1 U92 ( .A(n1089), .Z(n1131) );
  NAND2_X1 U31 ( .A1(n1612), .A2(n1777), .ZN(n1778) );
  INV_X1 U53 ( .A(n23), .ZN(n12) );
  BUF_X1 U11 ( .A(n897), .Z(n6) );
  BUF_X1 U47 ( .A(n5976), .Z(n56) );
  INV_X1 U35 ( .A(n53), .ZN(n15) );
  INV_X1 U67 ( .A(n49), .ZN(n50) );
  BUF_X1 U1071 ( .A(n1002), .Z(n2292) );
  AND2_X2 U61 ( .A1(is_clpx_i), .A2(clpx_img_i), .ZN(n1087) );
  MUX2_X1 U1184 ( .A(dot_op_b_i[0]), .B(dot_op_b_i[16]), .S(n1087), .Z(n1093)
         );
  CLKBUF_X2 U46 ( .A(n5992), .Z(n54) );
  NAND2_X1 U243 ( .A1(n6114), .A2(n1112), .ZN(n5113) );
  OAI21_X1 U2669 ( .B1(n4880), .B2(n5302), .A(n4962), .ZN(n2831) );
  NAND2_X2 U1178 ( .A1(n1086), .A2(n4731), .ZN(n4732) );
  INV_X1 U3 ( .A(n36), .ZN(n6111) );
  INV_X1 U4 ( .A(n6112), .ZN(n6117) );
  OR2_X1 U5 ( .A1(n2840), .A2(n2652), .ZN(n5615) );
  NAND2_X1 U8 ( .A1(n1084), .A2(n1932), .ZN(n1931) );
  BUF_X2 U13 ( .A(n145), .Z(n533) );
  INV_X1 U16 ( .A(n48), .ZN(n6115) );
  BUF_X2 U17 ( .A(n2621), .Z(n6116) );
  BUF_X1 U19 ( .A(n2866), .Z(n2879) );
  INV_X1 U22 ( .A(n3636), .ZN(n5941) );
  INV_X2 U25 ( .A(n2591), .ZN(n6112) );
  OR2_X1 U28 ( .A1(n6133), .A2(n530), .ZN(n6135) );
  INV_X1 U29 ( .A(n530), .ZN(n6132) );
  OR2_X1 U30 ( .A1(n6133), .A2(n530), .ZN(n6134) );
  INV_X1 U32 ( .A(n1611), .ZN(n6122) );
  OR2_X1 U34 ( .A1(n1514), .A2(n6129), .ZN(n6130) );
  OR2_X1 U43 ( .A1(n1164), .A2(n6124), .ZN(n6125) );
  INV_X1 U50 ( .A(n1164), .ZN(n6123) );
  BUF_X1 U54 ( .A(n2233), .Z(n6128) );
  INV_X2 U57 ( .A(n5112), .ZN(n6114) );
  INV_X1 U69 ( .A(n369), .ZN(n6156) );
  OR2_X1 U76 ( .A1(n6149), .A2(n429), .ZN(n6151) );
  OR2_X1 U83 ( .A1(n6137), .A2(n487), .ZN(n6139) );
  INV_X1 U84 ( .A(n487), .ZN(n6136) );
  OR2_X1 U85 ( .A1(n6137), .A2(n487), .ZN(n6138) );
  OR2_X1 U87 ( .A1(n6157), .A2(n369), .ZN(n6159) );
  OR2_X1 U94 ( .A1(n6157), .A2(n369), .ZN(n6158) );
  INV_X1 U95 ( .A(n429), .ZN(n6148) );
  OR2_X1 U96 ( .A1(n6149), .A2(n429), .ZN(n6150) );
  NAND2_X1 U103 ( .A1(n533), .A2(n549), .ZN(n552) );
  OR2_X1 U106 ( .A1(n6153), .A2(n514), .ZN(n6155) );
  INV_X1 U113 ( .A(n514), .ZN(n6152) );
  OR2_X1 U115 ( .A1(n6153), .A2(n514), .ZN(n6154) );
  NAND2_X1 U140 ( .A1(n124), .A2(n34), .ZN(n921) );
  AND3_X1 U151 ( .A1(n985), .A2(short_signed_i[0]), .A3(n144), .ZN(n2673) );
  INV_X1 U153 ( .A(n526), .ZN(n549) );
  INV_X1 U163 ( .A(n37), .ZN(n22) );
  INV_X1 U197 ( .A(n39), .ZN(n55) );
  INV_X1 U200 ( .A(n6143), .ZN(n6146) );
  XOR2_X1 U223 ( .A(n12), .B(dot_op_a_i[29]), .Z(n36) );
  BUF_X2 U248 ( .A(n2866), .Z(n6118) );
  MUX2_X1 U249 ( .A(op_a_i[31]), .B(op_a_i[15]), .S(n149), .Z(n985) );
  BUF_X2 U250 ( .A(n2866), .Z(n6119) );
  NAND2_X1 U279 ( .A1(n110), .A2(n166), .ZN(n6126) );
  MUX2_X1 U282 ( .A(dot_op_b_i[16]), .B(dot_op_b_i[0]), .S(n1087), .Z(n1126)
         );
  OR2_X1 U286 ( .A1(n6110), .A2(mulh_CS[2]), .ZN(n5218) );
  CLKBUF_X2 U289 ( .A(n2840), .Z(n29) );
  XNOR2_X1 U290 ( .A(n2866), .B(op_a_i[12]), .ZN(n6120) );
  XNOR2_X1 U296 ( .A(n2866), .B(op_a_i[12]), .ZN(n6121) );
  XNOR2_X1 U301 ( .A(n2866), .B(op_a_i[12]), .ZN(n5853) );
  AOI21_X1 U303 ( .B1(mulh_CS[1]), .B2(mulh_CS[2]), .A(mulh_CS[0]), .ZN(n166)
         );
  XNOR2_X1 U310 ( .A(n1083), .B(n1095), .ZN(n1932) );
  OR2_X1 U311 ( .A1(n1164), .A2(n6124), .ZN(n4845) );
  XNOR2_X1 U350 ( .A(n1118), .B(n57), .ZN(n6124) );
  XNOR2_X1 U357 ( .A(n1117), .B(n1118), .ZN(n4844) );
  NAND2_X1 U358 ( .A1(n110), .A2(n166), .ZN(n146) );
  OAI21_X1 U384 ( .B1(n2066), .B2(n2273), .A(n2065), .ZN(n6127) );
  OAI21_X1 U385 ( .B1(n2066), .B2(n2273), .A(n2065), .ZN(n5032) );
  OR2_X1 U388 ( .A1(n1514), .A2(n6129), .ZN(n2234) );
  XNOR2_X1 U389 ( .A(n1099), .B(n2147), .ZN(n6129) );
  OR2_X1 U1169 ( .A1(n1514), .A2(n6129), .ZN(n6131) );
  XNOR2_X1 U1232 ( .A(n1130), .B(n1099), .ZN(n2233) );
  OR2_X1 U1233 ( .A1(n6133), .A2(n530), .ZN(n562) );
  XNOR2_X1 U1234 ( .A(n107), .B(n542), .ZN(n6133) );
  XNOR2_X1 U1278 ( .A(n107), .B(n145), .ZN(n560) );
  OR2_X1 U2405 ( .A1(n6137), .A2(n487), .ZN(n737) );
  XNOR2_X1 U5199 ( .A(n111), .B(n730), .ZN(n6137) );
  XNOR2_X1 U5200 ( .A(n111), .B(n113), .ZN(n738) );
  AND2_X1 U5201 ( .A1(n2652), .A2(operator_i[2]), .ZN(n6140) );
  INV_X1 U5202 ( .A(n6112), .ZN(n6141) );
  INV_X1 U5203 ( .A(n6112), .ZN(n6142) );
  INV_X1 U5204 ( .A(n6112), .ZN(n6143) );
  INV_X1 U5205 ( .A(n6112), .ZN(n6144) );
  INV_X1 U5206 ( .A(n6112), .ZN(n6145) );
  AND2_X1 U5207 ( .A1(n2652), .A2(operator_i[2]), .ZN(n2591) );
  XNOR2_X1 U5208 ( .A(n4809), .B(n4808), .ZN(n6147) );
  INV_X1 U5209 ( .A(n36), .ZN(n57) );
  NOR2_X1 U5210 ( .A1(operator_i[1]), .A2(operator_i[0]), .ZN(n2652) );
  OR2_X1 U5211 ( .A1(n6149), .A2(n429), .ZN(n831) );
  XNOR2_X1 U5212 ( .A(n126), .B(n779), .ZN(n6149) );
  XNOR2_X1 U5213 ( .A(n126), .B(n125), .ZN(n832) );
  OR2_X1 U5214 ( .A1(n6153), .A2(n514), .ZN(n686) );
  XNOR2_X1 U5215 ( .A(n115), .B(n653), .ZN(n6153) );
  XNOR2_X1 U5216 ( .A(n115), .B(n114), .ZN(n687) );
  OR2_X1 U5217 ( .A1(n6157), .A2(n369), .ZN(n870) );
  XNOR2_X1 U5218 ( .A(n129), .B(n848), .ZN(n6157) );
  XNOR2_X1 U5219 ( .A(n129), .B(n128), .ZN(n871) );
  INV_X1 U5220 ( .A(n6160), .ZN(n6104) );
  OAI21_X1 U5221 ( .B1(n6101), .B2(n6102), .A(n6100), .ZN(n6160) );
endmodule


module riscv_alu_SHARED_INT_DIV0_FPU0 ( clk, rst_n, operator_i, operand_a_i, 
        operand_b_i, operand_c_i, vector_mode_i, bmask_a_i, bmask_b_i, 
        imm_vec_ext_i, is_clpx_i, is_subrot_i, clpx_shift_i, result_o, 
        comparison_result_o, ready_o, ex_ready_i, enable_i_BAR );
  input [6:0] operator_i;
  input [31:0] operand_a_i;
  input [31:0] operand_b_i;
  input [31:0] operand_c_i;
  input [1:0] vector_mode_i;
  input [4:0] bmask_a_i;
  input [4:0] bmask_b_i;
  input [1:0] imm_vec_ext_i;
  input [1:0] clpx_shift_i;
  output [31:0] result_o;
  input clk, rst_n, is_clpx_i, is_subrot_i, ex_ready_i, enable_i_BAR;
  output comparison_result_o, ready_o;
  wire   div_valid, ff_no_one, int_div_div_op_a_signed, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n33,
         n34, n38, n39, n40, n41, n42, n43, n44, n45, n46, n48, n52, n53, n54,
         n57, n58, n60, n61, n62, n64, n65, n66, n67, n68, n69, n71, n72, n73,
         n74, n75, n76, n77, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n98, n99, n100, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n120, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n222, n223,
         n224, n225, n226, n228, n229, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1324, n1325, n1327, n1328, n1329, n1330,
         n1331, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1403,
         n1404, n1405, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2358, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2408, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3042, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3113, n3114, n3115, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3886,
         n3887, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4083, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4198, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366;
  wire   [5:0] div_shift;
  wire   [5:0] cnt_result;
  wire   [31:0] ff_input;
  wire   [4:0] ff1_result;
  wire   [31:0] result_div;

  AND2_X1 U3 ( .A1(n240), .A2(n41), .ZN(n40) );
  AND2_X1 U4 ( .A1(n3115), .A2(n193), .ZN(n41) );
  NOR2_X1 U7 ( .A1(n1837), .A2(n44), .ZN(n43) );
  INV_X1 U9 ( .A(n71), .ZN(n72) );
  INV_X1 U11 ( .A(n53), .ZN(n54) );
  INV_X1 U14 ( .A(n2605), .ZN(n45) );
  INV_X1 U19 ( .A(n2848), .ZN(n64) );
  AND3_X2 U22 ( .A1(n4159), .A2(n398), .A3(n488), .ZN(div_valid) );
  BUF_X1 U23 ( .A(n1050), .Z(n3133) );
  NAND2_X1 U25 ( .A1(n34), .A2(n33), .ZN(n2886) );
  NAND2_X1 U26 ( .A1(n2412), .A2(n2376), .ZN(n33) );
  NAND2_X1 U27 ( .A1(n2399), .A2(n91), .ZN(n34) );
  NAND2_X1 U29 ( .A1(n38), .A2(n411), .ZN(n3177) );
  NAND2_X1 U30 ( .A1(n4275), .A2(n91), .ZN(n38) );
  NAND2_X1 U31 ( .A1(n397), .A2(n2496), .ZN(n2632) );
  NAND3_X1 U33 ( .A1(n39), .A2(n1711), .A3(n1712), .ZN(n2052) );
  NAND3_X1 U34 ( .A1(n353), .A2(n354), .A3(n1620), .ZN(n39) );
  NOR2_X2 U36 ( .A1(n2170), .A2(n3387), .ZN(n2217) );
  NAND2_X2 U41 ( .A1(n421), .A2(n365), .ZN(n1636) );
  NOR2_X2 U42 ( .A1(n1324), .A2(n1330), .ZN(n1341) );
  NAND3_X1 U43 ( .A1(n1834), .A2(n43), .A3(n1833), .ZN(n2418) );
  NAND2_X1 U44 ( .A1(n1835), .A2(n1832), .ZN(n44) );
  NAND3_X1 U45 ( .A1(n45), .A2(n2637), .A3(n281), .ZN(n2751) );
  NAND2_X1 U48 ( .A1(n46), .A2(n372), .ZN(n369) );
  AOI21_X1 U49 ( .B1(n371), .B2(n2598), .A(n198), .ZN(n46) );
  NAND2_X2 U50 ( .A1(n1364), .A2(n1363), .ZN(n2013) );
  INV_X1 U57 ( .A(operand_a_i[29]), .ZN(n53) );
  INV_X1 U60 ( .A(n1481), .ZN(n57) );
  AOI21_X1 U61 ( .B1(n1535), .B2(n1536), .A(n1031), .ZN(n58) );
  OR2_X1 U66 ( .A1(n2614), .A2(n3387), .ZN(n61) );
  AND3_X1 U67 ( .A1(n2852), .A2(n4037), .A3(n3190), .ZN(n62) );
  NAND2_X1 U69 ( .A1(n655), .A2(n467), .ZN(n65) );
  AND2_X1 U70 ( .A1(n335), .A2(operator_i[4]), .ZN(n66) );
  XNOR2_X1 U72 ( .A(n1286), .B(n68), .ZN(n478) );
  AND2_X1 U73 ( .A1(n1285), .A2(n1284), .ZN(n68) );
  INV_X1 U74 ( .A(n2747), .ZN(n69) );
  OR2_X1 U76 ( .A1(n2616), .A2(n2596), .ZN(n2615) );
  INV_X1 U79 ( .A(operand_a_i[18]), .ZN(n71) );
  NAND2_X1 U80 ( .A1(n2637), .A2(n281), .ZN(n73) );
  NAND2_X1 U82 ( .A1(n2632), .A2(n540), .ZN(n74) );
  OR2_X2 U83 ( .A1(n2023), .A2(n1933), .ZN(n2333) );
  NAND2_X1 U86 ( .A1(n397), .A2(n2496), .ZN(n77) );
  MUX2_X1 U93 ( .A(n2220), .B(n1746), .S(n1884), .Z(n2033) );
  OR2_X1 U96 ( .A1(n492), .A2(n482), .ZN(n80) );
  AND3_X1 U99 ( .A1(n333), .A2(n2290), .A3(n1288), .ZN(n81) );
  OAI21_X1 U102 ( .B1(n783), .B2(n784), .A(n135), .ZN(n1158) );
  CLKBUF_X1 U103 ( .A(n2885), .Z(n125) );
  MUX2_X1 U104 ( .A(n2400), .B(n2411), .S(n2376), .Z(n2885) );
  MUX2_X1 U105 ( .A(n2392), .B(n2419), .S(n91), .Z(n3463) );
  CLKBUF_X1 U107 ( .A(n2967), .Z(n3216) );
  MUX2_X1 U108 ( .A(n2400), .B(n2411), .S(n91), .Z(n3320) );
  OR2_X1 U110 ( .A1(n1782), .A2(n87), .ZN(n129) );
  OAI211_X1 U111 ( .C1(n1770), .C2(n1620), .A(n1561), .B(n1884), .ZN(n156) );
  BUF_X1 U112 ( .A(n1702), .Z(n2206) );
  NAND2_X1 U113 ( .A1(n391), .A2(n2695), .ZN(n2023) );
  INV_X1 U114 ( .A(n1635), .ZN(n86) );
  CLKBUF_X1 U118 ( .A(n1343), .Z(n1356) );
  NOR2_X1 U123 ( .A1(n660), .A2(n2641), .ZN(n635) );
  CLKBUF_X1 U130 ( .A(n2502), .Z(n4160) );
  CLKBUF_X1 U131 ( .A(n2553), .Z(n4071) );
  CLKBUF_X1 U133 ( .A(n2514), .Z(n4072) );
  CLKBUF_X1 U136 ( .A(operand_a_i[10]), .Z(n167) );
  CLKBUF_X1 U138 ( .A(operand_a_i[10]), .Z(n168) );
  NAND4_X1 U142 ( .A1(n115), .A2(n3286), .A3(n3285), .A4(n113), .ZN(
        result_o[21]) );
  OR2_X1 U144 ( .A1(n4286), .A2(n448), .ZN(n2385) );
  OR2_X1 U145 ( .A1(n4118), .A2(n447), .ZN(n3498) );
  OR2_X1 U146 ( .A1(n4118), .A2(n184), .ZN(n3792) );
  AND2_X1 U147 ( .A1(n3349), .A2(n480), .ZN(n103) );
  INV_X1 U148 ( .A(n4118), .ZN(n84) );
  CLKBUF_X1 U149 ( .A(n3010), .Z(n3590) );
  CLKBUF_X1 U151 ( .A(n3280), .Z(n222) );
  MUX2_X1 U152 ( .A(n2392), .B(n2419), .S(n2376), .Z(n3875) );
  CLKBUF_X1 U153 ( .A(n2994), .Z(n3763) );
  CLKBUF_X1 U154 ( .A(n2886), .Z(n3521) );
  OR2_X1 U156 ( .A1(n428), .A2(n1673), .ZN(n2419) );
  AOI21_X1 U158 ( .B1(n2072), .B2(n409), .A(n91), .ZN(n408) );
  NOR2_X1 U159 ( .A1(n1665), .A2(n431), .ZN(n430) );
  AND2_X1 U161 ( .A1(n140), .A2(n139), .ZN(n2072) );
  NOR2_X1 U162 ( .A1(n2071), .A2(n141), .ZN(n140) );
  OR2_X1 U163 ( .A1(n2097), .A2(n142), .ZN(n141) );
  OR2_X1 U164 ( .A1(n130), .A2(n1585), .ZN(n1782) );
  OAI211_X1 U166 ( .C1(n1770), .C2(n4294), .A(n1768), .B(n1769), .ZN(n1977) );
  OAI21_X1 U167 ( .B1(n2174), .B2(n94), .A(n93), .ZN(n2131) );
  OAI211_X1 U168 ( .C1(n1776), .C2(n1984), .A(n1678), .B(n133), .ZN(n132) );
  INV_X1 U174 ( .A(n1795), .ZN(n1260) );
  CLKBUF_X1 U175 ( .A(n1607), .Z(n1647) );
  NOR2_X1 U177 ( .A1(n2069), .A2(n2092), .ZN(n142) );
  INV_X1 U178 ( .A(n2127), .ZN(n94) );
  CLKBUF_X1 U179 ( .A(n2194), .Z(n157) );
  AOI21_X1 U180 ( .B1(n228), .B2(n82), .A(n1334), .ZN(n1895) );
  INV_X1 U187 ( .A(n2169), .ZN(n2230) );
  NAND2_X1 U190 ( .A1(n1788), .A2(n1730), .ZN(n1751) );
  INV_X1 U191 ( .A(n1620), .ZN(n87) );
  AOI21_X1 U192 ( .B1(n1606), .B2(n1605), .A(n1604), .ZN(n2115) );
  CLKBUF_X1 U193 ( .A(n1383), .Z(n1384) );
  NOR2_X1 U194 ( .A1(n1037), .A2(n1467), .ZN(n1492) );
  AND2_X1 U195 ( .A1(n1337), .A2(n1336), .ZN(n1338) );
  INV_X1 U196 ( .A(n1335), .ZN(n88) );
  AND2_X1 U197 ( .A1(n116), .A2(n493), .ZN(div_shift[1]) );
  OR2_X1 U199 ( .A1(n2834), .A2(n1230), .ZN(n1285) );
  XNOR2_X1 U200 ( .A(n484), .B(n105), .ZN(n3464) );
  NOR2_X1 U201 ( .A1(n1377), .A2(n1369), .ZN(n1392) );
  OR2_X1 U202 ( .A1(n3581), .A2(n1032), .ZN(n1472) );
  AND2_X1 U203 ( .A1(n3627), .A2(n1029), .ZN(n1535) );
  AND2_X1 U204 ( .A1(n3242), .A2(n1030), .ZN(n1031) );
  NOR2_X1 U205 ( .A1(n126), .A2(n1045), .ZN(n1382) );
  OR2_X1 U207 ( .A1(n3512), .A2(n1019), .ZN(n1528) );
  INV_X1 U208 ( .A(ff1_result[3]), .ZN(n105) );
  INV_X1 U210 ( .A(n1158), .ZN(n1123) );
  INV_X1 U211 ( .A(ff_no_one), .ZN(n112) );
  INV_X1 U213 ( .A(n1257), .ZN(n108) );
  AND2_X1 U214 ( .A1(n684), .A2(n778), .ZN(n685) );
  INV_X1 U215 ( .A(n1146), .ZN(n89) );
  NOR2_X1 U217 ( .A1(n1089), .A2(n1092), .ZN(n1145) );
  INV_X1 U218 ( .A(n3270), .ZN(n114) );
  NOR2_X1 U220 ( .A1(n643), .A2(n642), .ZN(n907) );
  NOR2_X2 U222 ( .A1(n2788), .A2(n2695), .ZN(n3076) );
  CLKBUF_X1 U223 ( .A(n2597), .Z(n2598) );
  NOR2_X1 U225 ( .A1(n4310), .A2(n3500), .ZN(n447) );
  NOR2_X1 U226 ( .A1(n4310), .A2(n2705), .ZN(n448) );
  NOR2_X1 U227 ( .A1(n4310), .A2(n3799), .ZN(n184) );
  INV_X1 U228 ( .A(n3373), .ZN(n123) );
  OR2_X1 U230 ( .A1(n532), .A2(is_clpx_i), .ZN(n579) );
  NOR2_X1 U232 ( .A1(n2733), .A2(n4130), .ZN(n4117) );
  NOR2_X2 U233 ( .A1(n2726), .A2(n2386), .ZN(n4059) );
  OR3_X1 U234 ( .A1(n2646), .A2(n500), .A3(n499), .ZN(n2726) );
  CLKBUF_X1 U235 ( .A(n2608), .Z(n4163) );
  CLKBUF_X1 U236 ( .A(n3949), .Z(n148) );
  BUF_X1 U238 ( .A(n2463), .Z(n4127) );
  INV_X1 U241 ( .A(n4108), .ZN(n100) );
  AND2_X1 U243 ( .A1(n2641), .A2(vector_mode_i[1]), .ZN(n2784) );
  INV_X1 U245 ( .A(n2561), .ZN(n163) );
  INV_X1 U248 ( .A(operand_a_i[13]), .ZN(n4101) );
  INV_X1 U250 ( .A(operand_b_i[13]), .ZN(n111) );
  INV_X1 U251 ( .A(operand_b_i[26]), .ZN(n3186) );
  CLKBUF_X1 U252 ( .A(operand_b_i[11]), .Z(n150) );
  NAND2_X1 U255 ( .A1(n2174), .A2(n2176), .ZN(n93) );
  OR2_X1 U256 ( .A1(n2058), .A2(n2150), .ZN(n1727) );
  NOR2_X1 U257 ( .A1(n1685), .A2(n1686), .ZN(n2058) );
  NAND2_X1 U258 ( .A1(n96), .A2(n95), .ZN(n654) );
  NAND2_X1 U259 ( .A1(n2949), .A2(n4098), .ZN(n95) );
  NAND2_X1 U260 ( .A1(n704), .A2(n4300), .ZN(n96) );
  NAND2_X1 U261 ( .A1(n99), .A2(n98), .ZN(n606) );
  NAND2_X1 U262 ( .A1(n169), .A2(n4108), .ZN(n98) );
  NAND2_X1 U263 ( .A1(n74), .A2(n100), .ZN(n99) );
  NAND3_X1 U264 ( .A1(n2615), .A2(n61), .A3(n2752), .ZN(n2770) );
  NAND2_X1 U265 ( .A1(n2520), .A2(n2519), .ZN(n2887) );
  NAND2_X1 U267 ( .A1(n104), .A2(n103), .ZN(result_o[10]) );
  NAND2_X1 U269 ( .A1(n492), .A2(n482), .ZN(n484) );
  NAND2_X1 U270 ( .A1(n361), .A2(n287), .ZN(n2089) );
  NAND2_X1 U271 ( .A1(n107), .A2(n106), .ZN(n236) );
  INV_X2 U272 ( .A(n2104), .ZN(n106) );
  NAND2_X1 U273 ( .A1(n2298), .A2(n92), .ZN(n107) );
  NAND3_X1 U274 ( .A1(n283), .A2(n2601), .A3(n3860), .ZN(n276) );
  NAND2_X1 U276 ( .A1(n332), .A2(n81), .ZN(n292) );
  NAND2_X1 U277 ( .A1(n109), .A2(n108), .ZN(n1795) );
  NAND2_X1 U278 ( .A1(n4299), .A2(n82), .ZN(n109) );
  NAND3_X1 U279 ( .A1(n2647), .A2(n4306), .A3(n2502), .ZN(n2608) );
  NAND2_X1 U280 ( .A1(n2565), .A2(n3387), .ZN(n2621) );
  NAND3_X1 U281 ( .A1(n2503), .A2(n2608), .A3(n52), .ZN(n2565) );
  NAND2_X1 U282 ( .A1(operand_a_i[13]), .A2(n111), .ZN(n2581) );
  NAND3_X1 U283 ( .A1(n80), .A2(n484), .A3(n112), .ZN(n490) );
  NAND2_X1 U286 ( .A1(n3258), .A2(n114), .ZN(n113) );
  NAND2_X1 U287 ( .A1(n3257), .A2(n3270), .ZN(n115) );
  NAND3_X1 U288 ( .A1(n3686), .A2(n495), .A3(n112), .ZN(n116) );
  NAND2_X1 U291 ( .A1(n630), .A2(n949), .ZN(n117) );
  NAND2_X1 U292 ( .A1(n120), .A2(n118), .ZN(n2001) );
  NAND2_X1 U293 ( .A1(n2052), .A2(n1884), .ZN(n118) );
  NAND2_X1 U294 ( .A1(n2047), .A2(n1635), .ZN(n120) );
  NOR2_X1 U295 ( .A1(n272), .A2(n273), .ZN(n271) );
  NAND2_X1 U296 ( .A1(n2593), .A2(n197), .ZN(n272) );
  OAI21_X1 U297 ( .B1(n2751), .B2(n123), .A(n122), .ZN(n2756) );
  NAND2_X1 U298 ( .A1(n2751), .A2(n2893), .ZN(n122) );
  OR2_X2 U299 ( .A1(n2636), .A2(n1016), .ZN(n1445) );
  NAND2_X1 U300 ( .A1(n124), .A2(n160), .ZN(n2597) );
  NAND2_X1 U301 ( .A1(n2540), .A2(n2541), .ZN(n124) );
  AND3_X1 U302 ( .A1(n61), .A2(n2752), .A3(n2753), .ZN(n2748) );
  NAND2_X1 U303 ( .A1(n126), .A2(n1045), .ZN(n1396) );
  NAND2_X1 U304 ( .A1(n3923), .A2(n126), .ZN(n3028) );
  XNOR2_X1 U305 ( .A(n686), .B(n685), .ZN(n126) );
  NAND2_X1 U306 ( .A1(n128), .A2(n127), .ZN(n130) );
  NAND3_X1 U307 ( .A1(n1629), .A2(n2171), .A3(n92), .ZN(n127) );
  NAND2_X1 U310 ( .A1(n132), .A2(n87), .ZN(n131) );
  OR2_X1 U311 ( .A1(n1636), .A2(n1985), .ZN(n133) );
  NAND2_X1 U312 ( .A1(n134), .A2(n1156), .ZN(n814) );
  NAND2_X1 U313 ( .A1(n1158), .A2(n89), .ZN(n134) );
  AOI21_X1 U314 ( .B1(n781), .B2(n782), .A(n780), .ZN(n135) );
  NAND2_X1 U315 ( .A1(n770), .A2(n782), .ZN(n784) );
  OAI21_X1 U317 ( .B1(n872), .B2(n867), .A(n873), .ZN(n136) );
  OAI21_X1 U318 ( .B1(n858), .B2(n885), .A(n859), .ZN(n866) );
  NOR2_X1 U319 ( .A1(n872), .A2(n868), .ZN(n672) );
  AOI21_X1 U320 ( .B1(n653), .B2(n137), .A(n652), .ZN(n1143) );
  NAND2_X1 U322 ( .A1(n138), .A2(n1536), .ZN(n1537) );
  INV_X1 U323 ( .A(n1031), .ZN(n138) );
  INV_X1 U324 ( .A(n1841), .ZN(n2070) );
  NAND2_X1 U325 ( .A1(n1841), .A2(n4288), .ZN(n139) );
  NAND2_X1 U327 ( .A1(n143), .A2(n82), .ZN(n1340) );
  XNOR2_X1 U328 ( .A(n144), .B(n1338), .ZN(n143) );
  AOI21_X1 U329 ( .B1(n1322), .B2(n88), .A(n1357), .ZN(n144) );
  XNOR2_X1 U330 ( .A(n832), .B(n145), .ZN(n3274) );
  AND2_X1 U331 ( .A1(n831), .A2(n840), .ZN(n145) );
  XNOR2_X1 U332 ( .A(n1011), .B(n146), .ZN(n3992) );
  AND2_X1 U333 ( .A1(n1010), .A2(n1009), .ZN(n146) );
  XNOR2_X1 U334 ( .A(n1071), .B(n147), .ZN(n4051) );
  AND2_X1 U335 ( .A1(n1070), .A2(n1090), .ZN(n147) );
  AOI21_X1 U336 ( .B1(n1535), .B2(n1536), .A(n1031), .ZN(n1468) );
  XNOR2_X1 U337 ( .A(n1162), .B(n151), .ZN(n3095) );
  AND2_X1 U338 ( .A1(n886), .A2(n885), .ZN(n151) );
  OR2_X1 U344 ( .A1(n3922), .A2(n1046), .ZN(n155) );
  NAND2_X1 U345 ( .A1(n1670), .A2(n156), .ZN(n2330) );
  BUF_X1 U346 ( .A(n2621), .Z(n158) );
  XNOR2_X1 U347 ( .A(n1103), .B(n159), .ZN(n3197) );
  AND2_X1 U348 ( .A1(n1102), .A2(n1149), .ZN(n159) );
  OR2_X1 U349 ( .A1(n2584), .A2(n2542), .ZN(n160) );
  INV_X1 U350 ( .A(n2759), .ZN(n161) );
  INV_X1 U351 ( .A(operand_a_i[12]), .ZN(n162) );
  NAND4_X1 U352 ( .A1(n1745), .A2(n1744), .A3(n1743), .A4(n1742), .ZN(n164) );
  INV_X1 U353 ( .A(n951), .ZN(n165) );
  OR2_X1 U354 ( .A1(n624), .A2(n623), .ZN(n166) );
  BUF_X2 U355 ( .A(n2632), .Z(n2949) );
  AOI21_X1 U356 ( .B1(n3672), .B2(n2372), .A(n2349), .ZN(n263) );
  OR2_X1 U357 ( .A1(n403), .A2(n402), .ZN(n401) );
  OR2_X1 U358 ( .A1(n2391), .A2(n91), .ZN(n2341) );
  NOR2_X1 U360 ( .A1(n2012), .A2(n532), .ZN(n427) );
  OR2_X1 U361 ( .A1(n2745), .A2(n2500), .ZN(n1267) );
  AOI21_X1 U363 ( .B1(n1386), .B2(n186), .A(n305), .ZN(n304) );
  INV_X1 U364 ( .A(operand_b_i[7]), .ZN(n231) );
  OAI21_X1 U365 ( .B1(n635), .B2(n1009), .A(n174), .ZN(n996) );
  CLKBUF_X1 U366 ( .A(n2614), .Z(n2618) );
  AND2_X1 U367 ( .A1(n2351), .A2(n2649), .ZN(n264) );
  AND3_X1 U368 ( .A1(n2852), .A2(n4037), .A3(n3190), .ZN(n284) );
  AND2_X1 U369 ( .A1(n1730), .A2(n425), .ZN(n366) );
  INV_X1 U370 ( .A(n1298), .ZN(n343) );
  OAI21_X1 U371 ( .B1(n1258), .B2(n1257), .A(n422), .ZN(n1566) );
  INV_X1 U372 ( .A(n423), .ZN(n422) );
  OAI21_X1 U373 ( .B1(n1257), .B2(n82), .A(n426), .ZN(n423) );
  NOR2_X1 U374 ( .A1(n1730), .A2(n424), .ZN(n365) );
  AND2_X1 U375 ( .A1(n394), .A2(n176), .ZN(n1581) );
  NOR2_X1 U376 ( .A1(n180), .A2(n1619), .ZN(n327) );
  NOR2_X1 U377 ( .A1(n90), .A2(n298), .ZN(n297) );
  AND2_X1 U378 ( .A1(n522), .A2(n515), .ZN(n298) );
  AND2_X1 U379 ( .A1(n1730), .A2(n416), .ZN(n415) );
  OR2_X1 U380 ( .A1(n3760), .A2(n3767), .ZN(n3761) );
  XNOR2_X1 U381 ( .A(n380), .B(n1362), .ZN(n379) );
  NOR2_X1 U382 ( .A1(n521), .A2(n433), .ZN(n432) );
  NOR2_X1 U383 ( .A1(n90), .A2(n517), .ZN(n433) );
  INV_X1 U384 ( .A(n396), .ZN(n395) );
  OAI21_X1 U385 ( .B1(n90), .B2(n176), .A(n516), .ZN(n396) );
  AND2_X1 U386 ( .A1(n4190), .A2(n319), .ZN(n318) );
  OR2_X1 U387 ( .A1(n4193), .A2(n4192), .ZN(n319) );
  NAND4_X1 U388 ( .A1(n1618), .A2(n1615), .A3(n1616), .A4(n1617), .ZN(n2304)
         );
  NOR2_X1 U390 ( .A1(n817), .A2(n4196), .ZN(n592) );
  INV_X1 U391 ( .A(n2589), .ZN(n212) );
  CLKBUF_X1 U392 ( .A(n2887), .Z(n2888) );
  OR2_X1 U393 ( .A1(n775), .A2(n588), .ZN(n589) );
  AND2_X1 U394 ( .A1(n3095), .A2(n1033), .ZN(n1034) );
  AND2_X1 U396 ( .A1(n2602), .A2(n2599), .ZN(n274) );
  NOR2_X1 U397 ( .A1(n2564), .A2(n214), .ZN(n277) );
  AND2_X1 U398 ( .A1(n264), .A2(n2367), .ZN(n261) );
  AND2_X1 U399 ( .A1(n264), .A2(n2725), .ZN(n260) );
  NAND2_X1 U400 ( .A1(n2421), .A2(n91), .ZN(n405) );
  OR2_X1 U402 ( .A1(n2584), .A2(n2620), .ZN(n2585) );
  AND2_X1 U403 ( .A1(n2604), .A2(n3387), .ZN(n2605) );
  OR2_X1 U404 ( .A1(n2605), .A2(n148), .ZN(n373) );
  OR2_X1 U405 ( .A1(bmask_b_i[4]), .A2(bmask_b_i[3]), .ZN(n1218) );
  INV_X1 U406 ( .A(n2159), .ZN(n341) );
  INV_X1 U407 ( .A(n2155), .ZN(n339) );
  NOR2_X1 U408 ( .A1(n1657), .A2(n532), .ZN(n356) );
  AOI21_X1 U409 ( .B1(n1636), .B2(n1795), .A(n1269), .ZN(n1814) );
  NOR2_X1 U410 ( .A1(n90), .A2(n515), .ZN(n393) );
  INV_X1 U411 ( .A(n2773), .ZN(n224) );
  AND2_X1 U412 ( .A1(n1657), .A2(n343), .ZN(n337) );
  OAI211_X1 U413 ( .C1(n2304), .C2(n321), .A(n1702), .B(n320), .ZN(n1943) );
  NAND2_X1 U414 ( .A1(n2169), .A2(n1566), .ZN(n2104) );
  OAI22_X1 U415 ( .A1(n1944), .A2(n2159), .B1(n342), .B2(n2160), .ZN(n1946) );
  OR2_X1 U416 ( .A1(n1938), .A2(n300), .ZN(n2109) );
  NAND4_X1 U417 ( .A1(n1723), .A2(n1722), .A3(n1720), .A4(n1721), .ZN(n2228)
         );
  INV_X1 U418 ( .A(n2158), .ZN(n2116) );
  INV_X1 U419 ( .A(n352), .ZN(n1713) );
  OAI21_X1 U420 ( .B1(n2194), .B2(n1619), .A(n355), .ZN(n352) );
  AND2_X1 U421 ( .A1(n1702), .A2(n1620), .ZN(n288) );
  OR2_X1 U422 ( .A1(n1775), .A2(n1614), .ZN(n1639) );
  OAI211_X1 U423 ( .C1(n1782), .C2(n1620), .A(n1781), .B(n1780), .ZN(n1978) );
  OR2_X1 U424 ( .A1(n1775), .A2(n4285), .ZN(n1781) );
  NOR2_X1 U425 ( .A1(n2000), .A2(n390), .ZN(n389) );
  INV_X1 U426 ( .A(n2695), .ZN(n390) );
  OAI211_X1 U428 ( .C1(n1316), .C2(n414), .A(n1619), .B(n413), .ZN(n420) );
  OAI21_X1 U429 ( .B1(n1354), .B2(n417), .A(n415), .ZN(n419) );
  NOR2_X1 U431 ( .A1(n487), .A2(n2648), .ZN(n4159) );
  NOR2_X1 U432 ( .A1(n3790), .A2(n3789), .ZN(n3791) );
  AND2_X1 U433 ( .A1(n3788), .A2(n4059), .ZN(n3789) );
  NOR2_X1 U434 ( .A1(n3680), .A2(n3679), .ZN(n3681) );
  INV_X1 U438 ( .A(n3941), .ZN(n246) );
  AOI21_X1 U439 ( .B1(n4011), .B2(n234), .A(n4065), .ZN(n233) );
  INV_X1 U440 ( .A(n4018), .ZN(n234) );
  AND2_X1 U441 ( .A1(n3594), .A2(n3593), .ZN(n229) );
  AND2_X1 U442 ( .A1(n2267), .A2(n2329), .ZN(n347) );
  AOI22_X1 U443 ( .A1(n2322), .A2(n2321), .B1(n2109), .B2(n2323), .ZN(n1950)
         );
  INV_X1 U444 ( .A(n330), .ZN(n329) );
  OAI21_X1 U445 ( .B1(n2209), .B2(n2207), .A(n2148), .ZN(n330) );
  NOR2_X1 U446 ( .A1(n241), .A2(n1910), .ZN(n1912) );
  NOR2_X1 U447 ( .A1(n1664), .A2(n2333), .ZN(n431) );
  INV_X1 U448 ( .A(n587), .ZN(n1180) );
  OR2_X1 U449 ( .A1(n75), .A2(n4097), .ZN(n530) );
  OR2_X1 U451 ( .A1(n1128), .A2(n2566), .ZN(n211) );
  NOR2_X1 U452 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U453 ( .A1(n636), .A2(n210), .ZN(n975) );
  AOI21_X1 U454 ( .B1(n2578), .B2(n2577), .A(n378), .ZN(n377) );
  AND3_X1 U455 ( .A1(n2588), .A2(n3902), .A3(n2589), .ZN(n285) );
  NOR2_X1 U456 ( .A1(n1069), .A2(n1068), .ZN(n1092) );
  NOR2_X1 U457 ( .A1(n708), .A2(n707), .ZN(n779) );
  NOR2_X1 U458 ( .A1(n213), .A2(n212), .ZN(n2977) );
  INV_X1 U459 ( .A(n2588), .ZN(n213) );
  CLKBUF_X1 U460 ( .A(n73), .Z(n2898) );
  INV_X1 U461 ( .A(n2603), .ZN(n2896) );
  NOR2_X1 U462 ( .A1(n667), .A2(n668), .ZN(n858) );
  NOR2_X1 U463 ( .A1(n975), .A2(n979), .ZN(n639) );
  OAI21_X1 U464 ( .B1(n76), .B2(n585), .A(n586), .ZN(n633) );
  NOR2_X1 U465 ( .A1(n270), .A2(n269), .ZN(n3364) );
  INV_X1 U466 ( .A(n273), .ZN(n282) );
  CLKBUF_X1 U467 ( .A(n2637), .Z(n2638) );
  NOR2_X1 U468 ( .A1(n3922), .A2(n1046), .ZN(n1388) );
  NOR2_X1 U469 ( .A1(n646), .A2(n647), .ZN(n897) );
  NOR2_X1 U470 ( .A1(n1311), .A2(n1306), .ZN(n1299) );
  INV_X1 U471 ( .A(n2504), .ZN(n2507) );
  CLKBUF_X1 U472 ( .A(n2503), .Z(n2497) );
  CLKBUF_X1 U473 ( .A(comparison_result_o), .Z(n2832) );
  INV_X1 U474 ( .A(n4127), .ZN(n4198) );
  INV_X1 U475 ( .A(n2292), .ZN(n409) );
  AOI21_X1 U477 ( .B1(n3280), .B2(n259), .A(n258), .ZN(n257) );
  AND2_X1 U478 ( .A1(n264), .A2(n2346), .ZN(n258) );
  AND2_X1 U479 ( .A1(n264), .A2(n2368), .ZN(n259) );
  NOR2_X1 U481 ( .A1(n1050), .A2(n1051), .ZN(n1330) );
  NOR2_X1 U482 ( .A1(n364), .A2(n1026), .ZN(n1493) );
  NOR2_X1 U483 ( .A1(n1467), .A2(n215), .ZN(n1460) );
  INV_X1 U484 ( .A(n1472), .ZN(n215) );
  INV_X1 U485 ( .A(n1034), .ZN(n400) );
  INV_X1 U486 ( .A(operator_i[1]), .ZN(n3834) );
  NOR2_X1 U488 ( .A1(n2335), .A2(bmask_a_i[1]), .ZN(n2725) );
  NOR2_X1 U489 ( .A1(n1795), .A2(n2156), .ZN(n1608) );
  INV_X1 U490 ( .A(n2003), .ZN(n342) );
  NOR2_X1 U491 ( .A1(n1794), .A2(n417), .ZN(n266) );
  OR2_X1 U492 ( .A1(div_valid), .A2(n2464), .ZN(n522) );
  NOR2_X1 U493 ( .A1(n311), .A2(n310), .ZN(n309) );
  INV_X1 U494 ( .A(n1386), .ZN(n311) );
  OAI21_X1 U495 ( .B1(n1386), .B2(n306), .A(n315), .ZN(n305) );
  INV_X1 U496 ( .A(n1391), .ZN(n315) );
  INV_X1 U497 ( .A(n313), .ZN(n306) );
  INV_X1 U498 ( .A(n310), .ZN(n307) );
  NOR2_X1 U499 ( .A1(n1390), .A2(n532), .ZN(n313) );
  INV_X1 U500 ( .A(n1387), .ZN(n314) );
  INV_X1 U501 ( .A(n327), .ZN(n323) );
  OR2_X1 U502 ( .A1(n1636), .A2(n92), .ZN(n1678) );
  INV_X1 U503 ( .A(n1017), .ZN(n382) );
  NOR2_X1 U504 ( .A1(n437), .A2(n1585), .ZN(n434) );
  AND2_X1 U505 ( .A1(n1731), .A2(n92), .ZN(n399) );
  INV_X1 U506 ( .A(n1535), .ZN(n216) );
  AND2_X1 U507 ( .A1(n289), .A2(n1702), .ZN(n1818) );
  INV_X1 U508 ( .A(n522), .ZN(n299) );
  INV_X1 U509 ( .A(n1317), .ZN(n414) );
  AND2_X1 U510 ( .A1(n2604), .A2(n2695), .ZN(n2595) );
  OR2_X1 U511 ( .A1(n373), .A2(n73), .ZN(n371) );
  OAI21_X1 U512 ( .B1(n4286), .B2(n317), .A(n3637), .ZN(n316) );
  NOR2_X1 U513 ( .A1(n4310), .A2(n3608), .ZN(n317) );
  AND2_X1 U514 ( .A1(n3179), .A2(n451), .ZN(n3180) );
  AND2_X1 U515 ( .A1(n4117), .A2(operand_c_i[7]), .ZN(n232) );
  OAI21_X1 U516 ( .B1(n4286), .B2(n188), .A(n3754), .ZN(n360) );
  NOR2_X1 U517 ( .A1(n3757), .A2(n457), .ZN(n3758) );
  AND2_X1 U518 ( .A1(n1636), .A2(n2013), .ZN(n293) );
  INV_X1 U519 ( .A(n1940), .ZN(n2320) );
  OAI211_X1 U520 ( .C1(n440), .C2(n1776), .A(n1559), .B(n439), .ZN(n1908) );
  NOR2_X1 U521 ( .A1(n82), .A2(vector_mode_i[1]), .ZN(n505) );
  OAI21_X1 U522 ( .B1(n157), .B2(n2160), .A(n340), .ZN(n1900) );
  AOI21_X1 U523 ( .B1(n3827), .B2(n3826), .A(n3825), .ZN(n3828) );
  INV_X1 U524 ( .A(n3495), .ZN(n3496) );
  OAI21_X1 U525 ( .B1(n4286), .B2(n189), .A(n547), .ZN(n367) );
  AND2_X1 U526 ( .A1(n3210), .A2(n3209), .ZN(n3211) );
  NAND4_X1 U527 ( .A1(n225), .A2(n2843), .A3(n462), .A4(n223), .ZN(
        result_o[29]) );
  NOR2_X1 U528 ( .A1(n3880), .A2(n179), .ZN(n226) );
  NOR2_X1 U529 ( .A1(n178), .A2(n3935), .ZN(n220) );
  NOR2_X1 U530 ( .A1(n3254), .A2(n3253), .ZN(n3255) );
  OAI21_X1 U531 ( .B1(n4286), .B2(n190), .A(n554), .ZN(n441) );
  AND2_X1 U532 ( .A1(n303), .A2(n302), .ZN(n2002) );
  OAI21_X1 U533 ( .B1(n2228), .B2(n2106), .A(n106), .ZN(n302) );
  OR2_X1 U534 ( .A1(n1838), .A2(n1620), .ZN(n418) );
  INV_X1 U535 ( .A(n2074), .ZN(n2075) );
  AND2_X1 U536 ( .A1(n2269), .A2(n2103), .ZN(n2034) );
  OR2_X1 U537 ( .A1(n1894), .A2(n1933), .ZN(n361) );
  INV_X1 U538 ( .A(n2304), .ZN(n2175) );
  NOR2_X1 U539 ( .A1(n1510), .A2(n1509), .ZN(n1511) );
  AND2_X1 U540 ( .A1(n1826), .A2(n4294), .ZN(n1509) );
  NOR2_X1 U541 ( .A1(n349), .A2(n347), .ZN(n346) );
  OAI211_X1 U542 ( .C1(n2188), .C2(n2023), .A(n1954), .B(n1953), .ZN(n2399) );
  AND4_X1 U543 ( .A1(n1949), .A2(n1950), .A3(n1952), .A4(n1951), .ZN(n1953) );
  NAND4_X1 U544 ( .A1(n2147), .A2(n2167), .A3(n2168), .A4(n329), .ZN(n2404) );
  AND2_X1 U545 ( .A1(n2166), .A2(n2165), .ZN(n2167) );
  NOR2_X1 U546 ( .A1(n2054), .A2(n443), .ZN(n2062) );
  OR2_X1 U547 ( .A1(n1912), .A2(n2280), .ZN(n429) );
  AND2_X1 U548 ( .A1(n1762), .A2(n238), .ZN(n237) );
  OR2_X2 U550 ( .A1(n2667), .A2(n3683), .ZN(n4038) );
  INV_X1 U551 ( .A(n1355), .ZN(n417) );
  INV_X1 U552 ( .A(n2000), .ZN(n1933) );
  INV_X1 U554 ( .A(n3350), .ZN(n398) );
  INV_X1 U555 ( .A(operand_a_i[7]), .ZN(n2543) );
  OR2_X2 U556 ( .A1(n2703), .A2(n3394), .ZN(n3228) );
  INV_X1 U560 ( .A(n2012), .ZN(n426) );
  NAND2_X1 U561 ( .A1(n669), .A2(vector_mode_i[0]), .ZN(n174) );
  INV_X1 U562 ( .A(vector_mode_i[1]), .ZN(n2695) );
  AND2_X1 U563 ( .A1(n296), .A2(n522), .ZN(n175) );
  OR2_X1 U564 ( .A1(div_valid), .A2(n3479), .ZN(n176) );
  AND2_X1 U565 ( .A1(n1296), .A2(n1295), .ZN(n177) );
  AND2_X1 U566 ( .A1(n3887), .A2(n3919), .ZN(n178) );
  AND2_X1 U567 ( .A1(n3850), .A2(n3855), .ZN(n179) );
  AND2_X1 U568 ( .A1(n1491), .A2(n1490), .ZN(n180) );
  AND2_X1 U569 ( .A1(n2369), .A2(n2352), .ZN(n181) );
  AND2_X1 U570 ( .A1(n1560), .A2(n92), .ZN(n182) );
  OR2_X1 U571 ( .A1(n4310), .A2(n3565), .ZN(n183) );
  XNOR2_X1 U573 ( .A(n1395), .B(n1380), .ZN(n185) );
  AND2_X1 U574 ( .A1(n307), .A2(n1387), .ZN(n186) );
  NOR2_X1 U575 ( .A1(n4310), .A2(n3768), .ZN(n187) );
  AND2_X1 U576 ( .A1(n514), .A2(n4091), .ZN(n2844) );
  NOR2_X1 U577 ( .A1(n4310), .A2(n3728), .ZN(n188) );
  NOR2_X1 U578 ( .A1(n4310), .A2(n3417), .ZN(n189) );
  NOR2_X1 U579 ( .A1(n4310), .A2(n3682), .ZN(n190) );
  AND2_X1 U580 ( .A1(n372), .A2(n3361), .ZN(n191) );
  AND2_X1 U581 ( .A1(n1564), .A2(n1565), .ZN(n192) );
  NAND2_X1 U582 ( .A1(n3521), .A2(n4012), .ZN(n193) );
  INV_X1 U583 ( .A(n425), .ZN(n424) );
  AND2_X1 U584 ( .A1(n1303), .A2(n1302), .ZN(n194) );
  AND2_X1 U585 ( .A1(n4301), .A2(n1331), .ZN(n195) );
  AND2_X1 U586 ( .A1(n1308), .A2(n1307), .ZN(n196) );
  AND2_X1 U587 ( .A1(n2918), .A2(n3119), .ZN(n197) );
  OR2_X1 U588 ( .A1(n4163), .A2(n3380), .ZN(n198) );
  OR2_X1 U589 ( .A1(n2313), .A2(n2260), .ZN(n199) );
  OR2_X1 U590 ( .A1(n1561), .A2(n1884), .ZN(n200) );
  INV_X1 U591 ( .A(n385), .ZN(int_div_div_op_a_signed) );
  NOR2_X1 U592 ( .A1(n4310), .A2(n3655), .ZN(n201) );
  AND2_X1 U593 ( .A1(n88), .A2(n1341), .ZN(n202) );
  OR2_X1 U594 ( .A1(n3762), .A2(n187), .ZN(n203) );
  AND2_X1 U595 ( .A1(n2647), .A2(n2651), .ZN(n2496) );
  OAI21_X1 U597 ( .B1(n206), .B2(n208), .A(n204), .ZN(n207) );
  AOI21_X1 U598 ( .B1(n2516), .B2(n205), .A(n2515), .ZN(n204) );
  INV_X1 U599 ( .A(n2513), .ZN(n205) );
  INV_X1 U600 ( .A(n2516), .ZN(n206) );
  NAND2_X1 U601 ( .A1(n207), .A2(n197), .ZN(n2519) );
  NAND2_X1 U602 ( .A1(n2512), .A2(n2511), .ZN(n208) );
  MUX2_X2 U603 ( .A(n2405), .B(n2406), .S(n91), .Z(n2968) );
  MUX2_X1 U604 ( .A(n2405), .B(n2406), .S(n2376), .Z(n2994) );
  NAND2_X1 U605 ( .A1(n2042), .A2(n476), .ZN(n2405) );
  OAI21_X1 U607 ( .B1(n999), .B2(n979), .A(n980), .ZN(n209) );
  NAND2_X1 U608 ( .A1(n210), .A2(n636), .ZN(n999) );
  NAND2_X1 U609 ( .A1(n633), .A2(n632), .ZN(n1009) );
  NAND2_X1 U610 ( .A1(n594), .A2(n479), .ZN(n637) );
  OAI21_X1 U611 ( .B1(n75), .B2(n3846), .A(n595), .ZN(n638) );
  NAND2_X1 U612 ( .A1(n593), .A2(n211), .ZN(n210) );
  OAI21_X1 U613 ( .B1(n58), .B2(n215), .A(n1471), .ZN(n1459) );
  NAND2_X1 U614 ( .A1(n1541), .A2(n216), .ZN(n1542) );
  NAND2_X1 U616 ( .A1(n217), .A2(n540), .ZN(n587) );
  INV_X1 U618 ( .A(n504), .ZN(n218) );
  AND2_X1 U619 ( .A1(n69), .A2(n2750), .ZN(n2890) );
  OAI211_X1 U620 ( .C1(n2618), .C2(vector_mode_i[1]), .A(n69), .B(n2617), .ZN(
        n3357) );
  INV_X1 U621 ( .A(n2615), .ZN(n2747) );
  NAND2_X1 U622 ( .A1(n2337), .A2(n181), .ZN(n2338) );
  AND2_X1 U623 ( .A1(n2652), .A2(n2651), .ZN(n219) );
  AOI22_X1 U624 ( .A1(n359), .A2(n356), .B1(n1298), .B2(n1619), .ZN(n355) );
  MUX2_X1 U625 ( .A(n2396), .B(n2415), .S(n91), .Z(n4015) );
  MUX2_X1 U626 ( .A(n1978), .B(n1977), .S(n2290), .Z(n2275) );
  NAND2_X1 U627 ( .A1(n2759), .A2(n191), .ZN(n2760) );
  INV_X1 U628 ( .A(n2751), .ZN(n372) );
  AND2_X1 U629 ( .A1(n2643), .A2(n4160), .ZN(n3361) );
  OAI211_X1 U630 ( .C1(n1681), .C2(n1984), .A(n1639), .B(n1678), .ZN(n1640) );
  OAI22_X1 U631 ( .A1(n1818), .A2(n437), .B1(n1814), .B2(n2178), .ZN(n1686) );
  AOI21_X2 U633 ( .B1(n2422), .B2(n2626), .A(n2499), .ZN(n4017) );
  INV_X2 U634 ( .A(n4006), .ZN(n4151) );
  NOR2_X2 U635 ( .A1(n2024), .A2(n4231), .ZN(n2321) );
  AND2_X1 U636 ( .A1(n375), .A2(n374), .ZN(n2619) );
  NAND2_X1 U637 ( .A1(n1632), .A2(n92), .ZN(n289) );
  OAI21_X1 U641 ( .B1(n4286), .B2(n464), .A(n4150), .ZN(n4191) );
  NAND2_X1 U642 ( .A1(n3177), .A2(n2368), .ZN(n252) );
  NAND2_X1 U643 ( .A1(n242), .A2(n1926), .ZN(n2411) );
  XNOR2_X1 U644 ( .A(n1309), .B(n196), .ZN(n452) );
  NAND2_X1 U645 ( .A1(n2766), .A2(n224), .ZN(n223) );
  NAND2_X1 U646 ( .A1(n2765), .A2(n2773), .ZN(n225) );
  NOR2_X1 U647 ( .A1(n1859), .A2(n1635), .ZN(n1685) );
  XNOR2_X1 U650 ( .A(n1333), .B(n195), .ZN(n228) );
  NOR2_X1 U653 ( .A1(n3976), .A2(n3652), .ZN(n2602) );
  NAND2_X1 U654 ( .A1(operand_a_i[7]), .A2(n231), .ZN(n2554) );
  NOR2_X1 U655 ( .A1(n4286), .A2(n232), .ZN(n4005) );
  NAND2_X1 U657 ( .A1(n235), .A2(n233), .ZN(result_o[25]) );
  NAND2_X1 U658 ( .A1(n4010), .A2(n4018), .ZN(n235) );
  NAND2_X1 U659 ( .A1(n280), .A2(n2600), .ZN(n273) );
  NAND2_X1 U660 ( .A1(n362), .A2(n363), .ZN(n3010) );
  OAI21_X1 U661 ( .B1(n1960), .B2(n1884), .A(n236), .ZN(n1894) );
  AOI21_X1 U662 ( .B1(n2725), .B2(n3463), .A(n401), .ZN(n2344) );
  OAI21_X1 U663 ( .B1(n4277), .B2(n2290), .A(n1750), .ZN(n2267) );
  NAND2_X1 U664 ( .A1(n1763), .A2(n237), .ZN(n2421) );
  NAND2_X1 U665 ( .A1(n1737), .A2(n239), .ZN(n238) );
  INV_X1 U666 ( .A(n2217), .ZN(n239) );
  NOR2_X1 U667 ( .A1(n405), .A2(n2347), .ZN(n402) );
  OAI21_X1 U668 ( .B1(n4286), .B2(n3461), .A(n3462), .ZN(n3497) );
  NAND2_X1 U669 ( .A1(operand_a_i[27]), .A2(n2848), .ZN(n2528) );
  NAND3_X1 U670 ( .A1(n255), .A2(n263), .A3(n2350), .ZN(n250) );
  NAND2_X1 U671 ( .A1(n1630), .A2(n1631), .ZN(n1632) );
  AOI21_X1 U673 ( .B1(n2887), .B2(n2604), .A(n2597), .ZN(n2614) );
  NOR2_X1 U674 ( .A1(n276), .A2(n278), .ZN(n275) );
  INV_X1 U675 ( .A(n3142), .ZN(n240) );
  INV_X1 U676 ( .A(n1663), .ZN(n241) );
  INV_X1 U677 ( .A(n243), .ZN(n242) );
  OAI21_X1 U678 ( .B1(n2334), .B2(n2207), .A(n1925), .ZN(n243) );
  INV_X1 U680 ( .A(n4130), .ZN(n295) );
  OAI22_X1 U681 ( .A1(n4226), .A2(n4127), .B1(n4229), .B2(n4115), .ZN(
        ff_input[0]) );
  AOI21_X2 U682 ( .B1(n1401), .B2(n82), .A(n1400), .ZN(n2161) );
  NAND2_X1 U683 ( .A1(n247), .A2(n244), .ZN(result_o[31]) );
  NAND2_X1 U684 ( .A1(n3942), .A2(n3941), .ZN(n247) );
  NAND4_X1 U685 ( .A1(n254), .A2(n253), .A3(n2354), .A4(n2355), .ZN(n248) );
  NAND2_X1 U688 ( .A1(n3217), .A2(n2372), .ZN(n253) );
  AOI21_X1 U689 ( .B1(n2968), .B2(n2368), .A(n2353), .ZN(n254) );
  AOI22_X1 U690 ( .A1(n3321), .A2(n2368), .B1(n3320), .B2(n2725), .ZN(n255) );
  AOI22_X1 U691 ( .A1(n2885), .A2(n261), .B1(n260), .B2(n2886), .ZN(n256) );
  OAI21_X1 U694 ( .B1(n2256), .B2(n2115), .A(n265), .ZN(n1947) );
  NAND2_X1 U695 ( .A1(n267), .A2(n266), .ZN(n265) );
  NAND2_X1 U696 ( .A1(n1354), .A2(n82), .ZN(n267) );
  NAND2_X1 U697 ( .A1(n267), .A2(n1355), .ZN(n2009) );
  NAND2_X1 U698 ( .A1(n2621), .A2(n2518), .ZN(n2506) );
  NOR2_X1 U700 ( .A1(n272), .A2(n268), .ZN(n2603) );
  INV_X1 U701 ( .A(n285), .ZN(n268) );
  NAND2_X1 U702 ( .A1(n2599), .A2(n2601), .ZN(n269) );
  NAND2_X1 U703 ( .A1(n282), .A2(n2602), .ZN(n270) );
  NOR2_X1 U704 ( .A1(n2564), .A2(n278), .ZN(n2639) );
  NAND4_X1 U705 ( .A1(n277), .A2(n275), .A3(n271), .A4(n274), .ZN(n2637) );
  NOR2_X1 U706 ( .A1(n4145), .A2(n3689), .ZN(n280) );
  NAND3_X1 U707 ( .A1(n2603), .A2(n2604), .A3(vector_mode_i[1]), .ZN(n281) );
  NAND3_X1 U708 ( .A1(n286), .A2(n2099), .A3(n456), .ZN(n4224) );
  NAND2_X1 U709 ( .A1(n2089), .A2(n2292), .ZN(n286) );
  NAND2_X1 U710 ( .A1(n1890), .A2(n1933), .ZN(n287) );
  AOI21_X1 U711 ( .B1(n288), .B2(n289), .A(n1634), .ZN(n1959) );
  NAND2_X1 U712 ( .A1(n1959), .A2(n1884), .ZN(n291) );
  NAND2_X1 U713 ( .A1(n2293), .A2(n1892), .ZN(n1907) );
  NAND2_X1 U714 ( .A1(n290), .A2(n1891), .ZN(n2293) );
  NAND2_X1 U715 ( .A1(n1890), .A2(n2000), .ZN(n290) );
  NAND2_X1 U716 ( .A1(n292), .A2(n291), .ZN(n1890) );
  AOI21_X1 U717 ( .B1(n1776), .B2(n2009), .A(n293), .ZN(n1708) );
  NAND2_X1 U718 ( .A1(n4100), .A2(n294), .ZN(ff_input[17]) );
  NAND2_X1 U719 ( .A1(n3882), .A2(operand_a_i[17]), .ZN(n294) );
  NAND2_X1 U722 ( .A1(div_shift[1]), .A2(div_valid), .ZN(n296) );
  NAND2_X1 U723 ( .A1(n1937), .A2(n383), .ZN(n1938) );
  NOR2_X1 U724 ( .A1(n1947), .A2(n1948), .ZN(n300) );
  NAND2_X1 U725 ( .A1(n301), .A2(n3681), .ZN(result_o[6]) );
  OAI21_X1 U726 ( .B1(n4286), .B2(n201), .A(n3677), .ZN(n301) );
  NAND2_X1 U727 ( .A1(n2002), .A2(n2108), .ZN(n2021) );
  NAND2_X1 U728 ( .A1(n2084), .A2(n2230), .ZN(n303) );
  OAI211_X1 U729 ( .C1(n1395), .C2(n312), .A(n308), .B(n304), .ZN(n2158) );
  NAND2_X1 U730 ( .A1(n1395), .A2(n309), .ZN(n308) );
  NAND2_X1 U731 ( .A1(n1390), .A2(n82), .ZN(n310) );
  NAND2_X1 U732 ( .A1(n314), .A2(n313), .ZN(n312) );
  NAND2_X1 U733 ( .A1(n316), .A2(n3641), .ZN(result_o[11]) );
  NAND2_X1 U734 ( .A1(n4191), .A2(n318), .ZN(result_o[0]) );
  NAND3_X1 U735 ( .A1(n2132), .A2(n2104), .A3(n92), .ZN(n320) );
  NAND2_X1 U736 ( .A1(n2105), .A2(n92), .ZN(n321) );
  NAND2_X1 U737 ( .A1(n323), .A2(n322), .ZN(n1741) );
  NAND2_X1 U738 ( .A1(n1716), .A2(n1619), .ZN(n322) );
  NAND3_X1 U740 ( .A1(n1716), .A2(n4294), .A3(n1619), .ZN(n324) );
  NAND2_X1 U741 ( .A1(n2176), .A2(n1620), .ZN(n325) );
  NAND2_X1 U742 ( .A1(n327), .A2(n4294), .ZN(n326) );
  NAND2_X1 U743 ( .A1(n331), .A2(n328), .ZN(n3788) );
  NAND2_X1 U744 ( .A1(n2404), .A2(n91), .ZN(n328) );
  NAND2_X1 U745 ( .A1(n2407), .A2(n2376), .ZN(n331) );
  NAND2_X1 U746 ( .A1(n1814), .A2(n4294), .ZN(n332) );
  NAND4_X1 U747 ( .A1(n332), .A2(n333), .A3(n1884), .A4(n1288), .ZN(n1319) );
  NAND2_X1 U748 ( .A1(n2004), .A2(n4282), .ZN(n333) );
  NAND2_X1 U749 ( .A1(n334), .A2(n3791), .ZN(result_o[16]) );
  OAI21_X1 U750 ( .B1(n4118), .B2(n203), .A(n3761), .ZN(n334) );
  NAND2_X1 U751 ( .A1(n335), .A2(operator_i[4]), .ZN(n2495) );
  INV_X1 U752 ( .A(operator_i[5]), .ZN(n335) );
  NAND2_X1 U753 ( .A1(n344), .A2(n343), .ZN(n2003) );
  NAND2_X1 U754 ( .A1(n338), .A2(n336), .ZN(n1927) );
  NAND2_X1 U755 ( .A1(n344), .A2(n337), .ZN(n336) );
  NAND2_X1 U756 ( .A1(n1944), .A2(n1619), .ZN(n338) );
  NAND2_X1 U757 ( .A1(n2003), .A2(n339), .ZN(n1799) );
  NAND2_X1 U758 ( .A1(n2003), .A2(n341), .ZN(n340) );
  MUX2_X1 U759 ( .A(n157), .B(n342), .S(n2262), .Z(n2242) );
  NAND2_X1 U760 ( .A1(n359), .A2(n82), .ZN(n344) );
  INV_X1 U761 ( .A(n2274), .ZN(n348) );
  NAND4_X1 U762 ( .A1(n348), .A2(n351), .A3(n346), .A4(n345), .ZN(n2397) );
  NAND2_X1 U763 ( .A1(n350), .A2(n4288), .ZN(n345) );
  NAND3_X1 U764 ( .A1(n2272), .A2(n199), .A3(n2273), .ZN(n349) );
  INV_X1 U765 ( .A(n2275), .ZN(n350) );
  INV_X1 U766 ( .A(n2266), .ZN(n351) );
  NAND2_X1 U767 ( .A1(n355), .A2(n2194), .ZN(n353) );
  NAND2_X1 U768 ( .A1(n355), .A2(n1619), .ZN(n354) );
  XNOR2_X1 U769 ( .A(n1297), .B(n177), .ZN(n359) );
  XNOR2_X1 U770 ( .A(n1304), .B(n194), .ZN(n358) );
  NAND2_X1 U771 ( .A1(n360), .A2(n3758), .ZN(result_o[5]) );
  NAND2_X1 U772 ( .A1(n4224), .A2(n2376), .ZN(n362) );
  NAND2_X1 U773 ( .A1(n2403), .A2(n91), .ZN(n363) );
  NAND2_X1 U774 ( .A1(n364), .A2(n1026), .ZN(n1494) );
  AOI21_X1 U775 ( .B1(n3628), .B2(n364), .A(n3054), .ZN(n3059) );
  XNOR2_X1 U776 ( .A(n861), .B(n455), .ZN(n364) );
  NAND2_X1 U777 ( .A1(n421), .A2(n366), .ZN(n1629) );
  INV_X1 U778 ( .A(n1587), .ZN(n1585) );
  NAND2_X1 U779 ( .A1(n367), .A2(n3460), .ZN(result_o[2]) );
  NAND2_X1 U780 ( .A1(n368), .A2(n2583), .ZN(n374) );
  NAND2_X1 U781 ( .A1(n2565), .A2(vector_mode_i[1]), .ZN(n368) );
  AOI21_X1 U782 ( .B1(n2755), .B2(n2754), .A(n369), .ZN(n2757) );
  NOR2_X1 U783 ( .A1(n73), .A2(n373), .ZN(n2753) );
  OAI21_X1 U784 ( .B1(n377), .B2(n376), .A(n2582), .ZN(n375) );
  NAND2_X1 U785 ( .A1(n3079), .A2(n2581), .ZN(n376) );
  NAND2_X1 U786 ( .A1(n2580), .A2(n2579), .ZN(n378) );
  INV_X1 U788 ( .A(n2770), .ZN(n2759) );
  NAND2_X1 U789 ( .A1(n379), .A2(n82), .ZN(n1364) );
  NAND2_X1 U790 ( .A1(n1358), .A2(n381), .ZN(n380) );
  NAND2_X1 U791 ( .A1(n202), .A2(n1322), .ZN(n381) );
  NAND2_X1 U792 ( .A1(n382), .A2(n1445), .ZN(n1446) );
  INV_X1 U793 ( .A(n2156), .ZN(n384) );
  NAND2_X1 U794 ( .A1(n2013), .A2(n384), .ZN(n383) );
  NAND2_X1 U795 ( .A1(n4274), .A2(n80), .ZN(n3353) );
  NAND2_X1 U796 ( .A1(n489), .A2(n490), .ZN(n513) );
  NOR2_X1 U797 ( .A1(n386), .A2(n385), .ZN(n3832) );
  NAND2_X1 U798 ( .A1(operand_a_i[31]), .A2(operator_i[0]), .ZN(n385) );
  MUX2_X1 U800 ( .A(n4228), .B(n4085), .S(n53), .Z(n4086) );
  MUX2_X1 U801 ( .A(n4099), .B(n4085), .S(n2522), .Z(n4081) );
  AND2_X2 U802 ( .A1(n391), .A2(n389), .ZN(n2329) );
  NAND2_X1 U803 ( .A1(n388), .A2(n387), .ZN(n2299) );
  NAND2_X1 U804 ( .A1(n2130), .A2(n86), .ZN(n387) );
  NAND3_X1 U805 ( .A1(n391), .A2(n389), .A3(n1884), .ZN(n388) );
  INV_X1 U806 ( .A(n1320), .ZN(n391) );
  MUX2_X1 U807 ( .A(n4228), .B(n4113), .S(n4095), .Z(n4096) );
  MUX2_X1 U808 ( .A(n4229), .B(n4113), .S(n4101), .Z(n4102) );
  MUX2_X1 U809 ( .A(n4099), .B(n4113), .S(n2561), .Z(n4104) );
  MUX2_X1 U810 ( .A(n4228), .B(n4113), .S(n2570), .Z(n3881) );
  MUX2_X1 U811 ( .A(n4099), .B(n4113), .S(n4071), .Z(n3845) );
  MUX2_X1 U812 ( .A(n4099), .B(n4113), .S(n4072), .Z(n4073) );
  MUX2_X1 U813 ( .A(n4099), .B(n4085), .S(n2521), .Z(n4080) );
  MUX2_X1 U814 ( .A(n4229), .B(n4085), .S(n585), .Z(n4077) );
  MUX2_X1 U815 ( .A(n4099), .B(n4085), .S(n4075), .Z(n4076) );
  MUX2_X1 U816 ( .A(n4228), .B(n4085), .S(n4067), .Z(n4068) );
  MUX2_X1 U817 ( .A(n4085), .B(n4229), .S(operand_a_i[11]), .Z(n3884) );
  MUX2_X1 U818 ( .A(n4085), .B(n4229), .S(operand_a_i[26]), .Z(n4078) );
  NAND3_X1 U819 ( .A1(n514), .A2(n393), .A3(n4091), .ZN(n392) );
  NAND3_X1 U820 ( .A1(n514), .A2(n4091), .A3(div_valid), .ZN(n394) );
  INV_X1 U821 ( .A(n219), .ZN(n2745) );
  AOI22_X1 U822 ( .A1(n1636), .A2(n182), .B1(n1629), .B2(n399), .ZN(n435) );
  NAND2_X1 U823 ( .A1(n435), .A2(n1702), .ZN(n1770) );
  NAND2_X1 U824 ( .A1(n1461), .A2(n400), .ZN(n1462) );
  NAND2_X1 U825 ( .A1(n405), .A2(n406), .ZN(n4123) );
  OAI21_X1 U826 ( .B1(n406), .B2(n2347), .A(n404), .ZN(n403) );
  AND2_X1 U827 ( .A1(n2342), .A2(bmask_a_i[4]), .ZN(n404) );
  NAND2_X1 U828 ( .A1(n2390), .A2(n2376), .ZN(n406) );
  NAND2_X1 U830 ( .A1(n2063), .A2(n2292), .ZN(n407) );
  OAI21_X1 U831 ( .B1(n4281), .B2(n410), .A(n408), .ZN(n411) );
  INV_X1 U832 ( .A(n2072), .ZN(n410) );
  NAND2_X1 U833 ( .A1(n412), .A2(n1317), .ZN(n2256) );
  NAND2_X1 U834 ( .A1(n1316), .A2(n82), .ZN(n412) );
  NAND2_X1 U835 ( .A1(n1317), .A2(n532), .ZN(n413) );
  NAND2_X1 U836 ( .A1(n1355), .A2(n532), .ZN(n416) );
  NAND3_X1 U837 ( .A1(n1571), .A2(n418), .A3(n1570), .ZN(n2306) );
  NAND2_X1 U838 ( .A1(n419), .A2(n420), .ZN(n1838) );
  NAND2_X1 U839 ( .A1(n1258), .A2(n427), .ZN(n421) );
  NAND2_X1 U840 ( .A1(n1257), .A2(n426), .ZN(n425) );
  INV_X1 U841 ( .A(n493), .ZN(n489) );
  OAI21_X1 U842 ( .B1(n492), .B2(ff_no_one), .A(n385), .ZN(n493) );
  NAND4_X1 U843 ( .A1(n1671), .A2(n430), .A3(n1672), .A4(n429), .ZN(n428) );
  NAND2_X1 U844 ( .A1(n518), .A2(n517), .ZN(n1584) );
  INV_X1 U845 ( .A(n2169), .ZN(n1635) );
  NAND2_X1 U846 ( .A1(n435), .A2(n434), .ZN(n436) );
  NAND3_X1 U847 ( .A1(n438), .A2(n200), .A3(n436), .ZN(n1935) );
  NAND2_X1 U848 ( .A1(n1635), .A2(n87), .ZN(n437) );
  NAND2_X1 U849 ( .A1(n1908), .A2(n1884), .ZN(n438) );
  OR2_X1 U850 ( .A1(n1775), .A2(n1764), .ZN(n439) );
  NOR2_X1 U851 ( .A1(n1556), .A2(n2106), .ZN(n440) );
  NAND2_X1 U852 ( .A1(n441), .A2(n3716), .ZN(result_o[1]) );
  OAI21_X1 U853 ( .B1(n4366), .B2(n3531), .A(n477), .ZN(result_o[24]) );
  NOR2_X1 U854 ( .A1(n4307), .A2(operator_i[4]), .ZN(n2502) );
  NOR2_X1 U855 ( .A1(n1043), .A2(n1044), .ZN(n1369) );
  XNOR2_X1 U856 ( .A(n875), .B(n442), .ZN(n3779) );
  AND2_X1 U857 ( .A1(n874), .A2(n873), .ZN(n442) );
  AND2_X1 U858 ( .A1(n2296), .A2(n2053), .ZN(n443) );
  AND2_X1 U859 ( .A1(n846), .A2(n845), .ZN(n444) );
  AND2_X1 U860 ( .A1(n727), .A2(n744), .ZN(n445) );
  AND2_X1 U861 ( .A1(n1061), .A2(n1091), .ZN(n446) );
  AND2_X1 U862 ( .A1(n797), .A2(n810), .ZN(n449) );
  OR2_X1 U863 ( .A1(n83), .A2(n4198), .ZN(n450) );
  OR2_X1 U864 ( .A1(n3178), .A2(n4192), .ZN(n451) );
  AND2_X1 U865 ( .A1(n750), .A2(n749), .ZN(n453) );
  AND2_X1 U866 ( .A1(n709), .A2(n777), .ZN(n454) );
  AND2_X1 U867 ( .A1(n860), .A2(n859), .ZN(n455) );
  OR2_X1 U868 ( .A1(n2098), .A2(n86), .ZN(n456) );
  AND2_X1 U869 ( .A1(n3756), .A2(n3755), .ZN(n457) );
  OR2_X1 U870 ( .A1(n83), .A2(n4194), .ZN(n458) );
  OR2_X1 U871 ( .A1(n83), .A2(operand_b_i[16]), .ZN(n459) );
  OR2_X1 U872 ( .A1(n3965), .A2(n4192), .ZN(n460) );
  OR2_X1 U873 ( .A1(n3753), .A2(n4182), .ZN(n461) );
  OR2_X1 U874 ( .A1(n3490), .A2(n4192), .ZN(n462) );
  NAND2_X1 U875 ( .A1(n2060), .A2(n2108), .ZN(n463) );
  INV_X1 U876 ( .A(n1729), .ZN(n1560) );
  AND2_X1 U877 ( .A1(n4117), .A2(operand_c_i[0]), .ZN(n464) );
  OR2_X1 U878 ( .A1(n83), .A2(operand_b_i[17]), .ZN(n465) );
  OR2_X1 U879 ( .A1(n83), .A2(operand_b_i[29]), .ZN(n466) );
  OR2_X1 U880 ( .A1(n83), .A2(operand_b_i[30]), .ZN(n467) );
  OR2_X1 U881 ( .A1(n83), .A2(operand_b_i[20]), .ZN(n468) );
  OR2_X1 U883 ( .A1(n83), .A2(n64), .ZN(n469) );
  INV_X1 U884 ( .A(operand_b_i[7]), .ZN(n588) );
  OR2_X1 U885 ( .A1(n83), .A2(operand_b_i[23]), .ZN(n470) );
  OR2_X1 U886 ( .A1(n83), .A2(operand_b_i[31]), .ZN(n471) );
  OR2_X1 U887 ( .A1(n2356), .A2(bmask_a_i[4]), .ZN(n472) );
  OR2_X1 U888 ( .A1(n83), .A2(operand_b_i[28]), .ZN(n473) );
  OR2_X1 U889 ( .A1(n83), .A2(operand_b_i[22]), .ZN(n474) );
  OR2_X1 U890 ( .A1(n1818), .A2(n1817), .ZN(n475) );
  OR2_X1 U891 ( .A1(n2275), .A2(n2254), .ZN(n476) );
  AND2_X1 U892 ( .A1(n3555), .A2(n3554), .ZN(n477) );
  OR2_X1 U893 ( .A1(n83), .A2(operand_b_i[25]), .ZN(n479) );
  AND2_X1 U894 ( .A1(n3345), .A2(n3344), .ZN(n480) );
  AND4_X1 U895 ( .A1(n2732), .A2(n2731), .A3(n2730), .A4(n2729), .ZN(n481) );
  NOR2_X1 U896 ( .A1(n83), .A2(operand_b_i[24]), .ZN(n591) );
  AND2_X1 U897 ( .A1(n2576), .A2(n2575), .ZN(n2577) );
  INV_X1 U898 ( .A(n3364), .ZN(n2640) );
  INV_X1 U899 ( .A(operand_b_i[23]), .ZN(n2505) );
  OR2_X1 U900 ( .A1(operand_a_i[31]), .A2(operand_b_i[31]), .ZN(n2524) );
  NOR2_X1 U901 ( .A1(n627), .A2(n628), .ZN(n956) );
  INV_X1 U902 ( .A(operand_a_i[17]), .ZN(n538) );
  INV_X1 U903 ( .A(operand_b_i[17]), .ZN(n2508) );
  NOR2_X1 U905 ( .A1(n624), .A2(n623), .ZN(n933) );
  NOR2_X1 U907 ( .A1(n931), .A2(n933), .ZN(n949) );
  AOI21_X1 U908 ( .B1(n2994), .B2(n2372), .A(n472), .ZN(n2361) );
  MUX2_X1 U909 ( .A(n2407), .B(n2404), .S(n2376), .Z(n2967) );
  INV_X1 U910 ( .A(n3754), .ZN(n3755) );
  AND2_X1 U911 ( .A1(n3835), .A2(n498), .ZN(n3837) );
  OAI22_X1 U912 ( .A1(n3753), .A2(n4184), .B1(n3552), .B2(n3551), .ZN(n3553)
         );
  INV_X1 U913 ( .A(operand_b_i[2]), .ZN(n3438) );
  NOR2_X1 U914 ( .A1(n335), .A2(operator_i[4]), .ZN(n502) );
  NOR2_X1 U915 ( .A1(n2944), .A2(n4337), .ZN(n4006) );
  INV_X1 U916 ( .A(n2875), .ZN(n2876) );
  OAI21_X1 U917 ( .B1(n3207), .B2(n3206), .A(n461), .ZN(n3208) );
  INV_X1 U918 ( .A(n3553), .ZN(n3554) );
  INV_X1 U919 ( .A(n3000), .ZN(n3001) );
  INV_X1 U920 ( .A(n3066), .ZN(n3067) );
  INV_X1 U921 ( .A(n3103), .ZN(n3108) );
  AND2_X1 U922 ( .A1(n3638), .A2(n3624), .ZN(n3639) );
  AND2_X1 U923 ( .A1(n4117), .A2(operand_c_i[3]), .ZN(n3461) );
  INV_X1 U924 ( .A(n3454), .ZN(n3459) );
  AOI21_X1 U925 ( .B1(n3715), .B2(n3714), .A(n3713), .ZN(n3716) );
  OR2_X1 U926 ( .A1(div_valid), .A2(n3438), .ZN(n517) );
  INV_X1 U927 ( .A(vector_mode_i[0]), .ZN(n2641) );
  INV_X1 U928 ( .A(bmask_b_i[4]), .ZN(n1196) );
  OAI21_X1 U929 ( .B1(n2420), .B2(n2376), .A(n2341), .ZN(n4193) );
  OAI211_X1 U930 ( .C1(n3965), .C2(n2386), .A(n2340), .B(n2339), .ZN(n2384) );
  INV_X1 U931 ( .A(n3313), .ZN(n3314) );
  AND2_X1 U932 ( .A1(n2877), .A2(n2876), .ZN(n2878) );
  INV_X1 U933 ( .A(n3208), .ZN(n3209) );
  AND2_X1 U934 ( .A1(n2884), .A2(n2946), .ZN(n2963) );
  AND2_X1 U935 ( .A1(n3009), .A2(n3026), .ZN(n3038) );
  AND2_X1 U936 ( .A1(n3002), .A2(n3001), .ZN(n3003) );
  AND2_X1 U937 ( .A1(n3108), .A2(n3107), .ZN(n3109) );
  AND2_X1 U938 ( .A1(n3252), .A2(n3251), .ZN(n3253) );
  NOR2_X1 U939 ( .A1(n3640), .A2(n3639), .ZN(n3641) );
  AND2_X1 U940 ( .A1(n3459), .A2(n3458), .ZN(n3460) );
  AND2_X1 U941 ( .A1(n2741), .A2(n2740), .ZN(n2742) );
  INV_X1 U943 ( .A(n525), .ZN(n526) );
  AND2_X1 U944 ( .A1(n3524), .A2(n3523), .ZN(n3525) );
  INV_X1 U945 ( .A(n3312), .ZN(n3317) );
  NOR2_X1 U946 ( .A1(n2879), .A2(n2878), .ZN(n2880) );
  NOR2_X1 U947 ( .A1(n2963), .A2(n2962), .ZN(n2964) );
  NOR2_X1 U948 ( .A1(n3038), .A2(n3037), .ZN(n3039) );
  NOR2_X1 U950 ( .A1(n3004), .A2(n3003), .ZN(n3005) );
  NOR2_X1 U951 ( .A1(n3070), .A2(n3069), .ZN(n3071) );
  INV_X1 U952 ( .A(n3589), .ZN(n3594) );
  AND2_X1 U953 ( .A1(n2162), .A2(n2025), .ZN(n1853) );
  NOR2_X1 U954 ( .A1(n3526), .A2(n3525), .ZN(n3527) );
  AND2_X1 U955 ( .A1(n481), .A2(n2737), .ZN(n2738) );
  OAI21_X1 U956 ( .B1(n3213), .B2(n3212), .A(n3211), .ZN(result_o[26]) );
  NOR2_X1 U957 ( .A1(n1853), .A2(n1852), .ZN(n1854) );
  AOI21_X1 U958 ( .B1(n1995), .B2(n2170), .A(n1994), .ZN(n1996) );
  AND2_X1 U959 ( .A1(n1552), .A2(n2230), .ZN(n1553) );
  NOR2_X1 U960 ( .A1(enable_i_BAR), .A2(n4306), .ZN(n488) );
  AOI21_X1 U961 ( .B1(n2060), .B2(n4288), .A(n1707), .ZN(n1726) );
  AOI21_X1 U962 ( .B1(n2233), .B2(n4233), .A(n2075), .ZN(n2088) );
  AND3_X1 U963 ( .A1(n1998), .A2(n1997), .A3(n1996), .ZN(n1999) );
  AOI21_X1 U964 ( .B1(n2291), .B2(n1884), .A(n1553), .ZN(n1554) );
  OAI21_X1 U965 ( .B1(n2289), .B2(n2023), .A(n2022), .ZN(n2398) );
  INV_X1 U966 ( .A(ff1_result[2]), .ZN(n482) );
  INV_X1 U967 ( .A(n513), .ZN(n483) );
  NAND2_X1 U968 ( .A1(n3464), .A2(n112), .ZN(n511) );
  NAND2_X1 U969 ( .A1(n483), .A2(n511), .ZN(n4091) );
  NOR2_X1 U970 ( .A1(n4274), .A2(ff1_result[3]), .ZN(n486) );
  INV_X1 U971 ( .A(ff1_result[4]), .ZN(n485) );
  NAND2_X1 U972 ( .A1(n486), .A2(n485), .ZN(n3717) );
  OAI21_X1 U973 ( .B1(n486), .B2(n485), .A(n3717), .ZN(n3797) );
  OR2_X1 U974 ( .A1(n3797), .A2(ff_no_one), .ZN(n4089) );
  XNOR2_X1 U975 ( .A(n4089), .B(n4091), .ZN(div_shift[4]) );
  NAND2_X1 U977 ( .A1(operator_i[4]), .A2(n4307), .ZN(n3350) );
  XNOR2_X1 U978 ( .A(n490), .B(n493), .ZN(div_shift[2]) );
  NAND2_X1 U980 ( .A1(n494), .A2(n385), .ZN(n495) );
  AND2_X1 U981 ( .A1(ff1_result[0]), .A2(ff1_result[1]), .ZN(n491) );
  INV_X1 U983 ( .A(operand_a_i[0]), .ZN(n2463) );
  OR2_X1 U984 ( .A1(n494), .A2(n385), .ZN(n496) );
  AND2_X1 U985 ( .A1(n496), .A2(n495), .ZN(div_shift[0]) );
  INV_X1 U986 ( .A(div_valid), .ZN(n515) );
  INV_X1 U987 ( .A(operator_i[3]), .ZN(n497) );
  INV_X1 U988 ( .A(operator_i[6]), .ZN(n2651) );
  INV_X1 U989 ( .A(n502), .ZN(n2500) );
  INV_X1 U991 ( .A(operator_i[0]), .ZN(n4131) );
  NOR2_X1 U992 ( .A1(n4131), .A2(operator_i[1]), .ZN(n2740) );
  NAND2_X1 U993 ( .A1(n2740), .A2(n4160), .ZN(n2646) );
  INV_X1 U994 ( .A(n487), .ZN(n500) );
  INV_X1 U995 ( .A(operator_i[2]), .ZN(n498) );
  NAND2_X1 U996 ( .A1(n498), .A2(n4306), .ZN(n499) );
  OR2_X1 U997 ( .A1(operator_i[6]), .A2(operator_i[3]), .ZN(n2642) );
  NOR2_X1 U998 ( .A1(n3350), .A2(n2642), .ZN(n3835) );
  OAI21_X1 U999 ( .B1(n52), .B2(n498), .A(n4290), .ZN(n3833) );
  AND2_X1 U1000 ( .A1(n3833), .A2(n2726), .ZN(n503) );
  NAND2_X1 U1002 ( .A1(n2651), .A2(n487), .ZN(n504) );
  NAND3_X1 U1003 ( .A1(n2660), .A2(n502), .A3(n498), .ZN(n2733) );
  NAND2_X1 U1004 ( .A1(n4131), .A2(operator_i[1]), .ZN(n4130) );
  OAI211_X1 U1005 ( .C1(n1267), .C2(n3683), .A(n503), .B(n4009), .ZN(n575) );
  OAI21_X1 U1006 ( .B1(div_valid), .B2(operand_b_i[4]), .A(n1871), .ZN(n506)
         );
  INV_X1 U1007 ( .A(n506), .ZN(n507) );
  OAI21_X1 U1008 ( .B1(div_shift[4]), .B2(n515), .A(n507), .ZN(n510) );
  INV_X1 U1009 ( .A(n579), .ZN(n508) );
  NAND2_X1 U1010 ( .A1(n508), .A2(bmask_b_i[4]), .ZN(n509) );
  NAND2_X1 U1011 ( .A1(n510), .A2(n509), .ZN(n1320) );
  INV_X1 U1012 ( .A(n511), .ZN(n512) );
  NAND2_X1 U1013 ( .A1(n513), .A2(n512), .ZN(n514) );
  INV_X1 U1014 ( .A(operand_b_i[3]), .ZN(n3479) );
  NAND2_X1 U1015 ( .A1(n1605), .A2(n515), .ZN(n582) );
  INV_X1 U1016 ( .A(n582), .ZN(n519) );
  NOR2_X1 U1017 ( .A1(n579), .A2(n1109), .ZN(n1579) );
  AOI21_X1 U1018 ( .B1(n519), .B2(operand_b_i[19]), .A(n1579), .ZN(n516) );
  INV_X1 U1019 ( .A(n2784), .ZN(n2668) );
  NOR2_X1 U1020 ( .A1(n2000), .A2(n2668), .ZN(n2130) );
  NAND2_X1 U1021 ( .A1(div_shift[2]), .A2(div_valid), .ZN(n518) );
  NOR2_X1 U1023 ( .A1(n1594), .A2(div_valid), .ZN(n1872) );
  INV_X1 U1024 ( .A(n1872), .ZN(n1603) );
  NAND2_X1 U1025 ( .A1(n519), .A2(n4194), .ZN(n520) );
  OR2_X1 U1026 ( .A1(n579), .A2(n1076), .ZN(n1868) );
  OAI211_X1 U1027 ( .C1(n3186), .C2(n1603), .A(n520), .B(n1868), .ZN(n521) );
  INV_X1 U1028 ( .A(operand_b_i[1]), .ZN(n2464) );
  NAND2_X1 U1029 ( .A1(n1872), .A2(n110), .ZN(n524) );
  INV_X1 U1030 ( .A(bmask_b_i[1]), .ZN(n729) );
  OR2_X1 U1031 ( .A1(n579), .A2(n729), .ZN(n1873) );
  NAND3_X1 U1032 ( .A1(n82), .A2(is_clpx_i), .A3(clpx_shift_i[1]), .ZN(n523)
         );
  AND2_X1 U1033 ( .A1(n1873), .A2(n523), .ZN(n1596) );
  OAI211_X1 U1034 ( .C1(n2508), .C2(n582), .A(n524), .B(n1596), .ZN(n525) );
  OR2_X1 U1035 ( .A1(n2217), .A2(n2178), .ZN(n1810) );
  NAND2_X1 U1037 ( .A1(n2632), .A2(n540), .ZN(n558) );
  NAND2_X1 U1039 ( .A1(n1205), .A2(n4198), .ZN(n529) );
  NAND2_X1 U1040 ( .A1(n2949), .A2(n4127), .ZN(n528) );
  NAND2_X1 U1041 ( .A1(n529), .A2(n528), .ZN(n531) );
  NAND2_X1 U1042 ( .A1(n77), .A2(is_subrot_i), .ZN(n679) );
  INV_X1 U1043 ( .A(operand_a_i[16]), .ZN(n4097) );
  NAND2_X1 U1044 ( .A1(n531), .A2(n530), .ZN(n537) );
  INV_X1 U1045 ( .A(n1181), .ZN(n1207) );
  MUX2_X1 U1046 ( .A(n1207), .B(n1128), .S(operand_b_i[0]), .Z(n533) );
  NAND2_X1 U1047 ( .A1(n533), .A2(n459), .ZN(n536) );
  NOR2_X1 U1048 ( .A1(n537), .A2(n536), .ZN(n548) );
  OR2_X1 U1050 ( .A1(n2495), .A2(n52), .ZN(n535) );
  OAI21_X1 U1051 ( .B1(n2745), .B2(n535), .A(n1180), .ZN(n634) );
  INV_X1 U1052 ( .A(n634), .ZN(n551) );
  NAND2_X1 U1053 ( .A1(n537), .A2(n536), .ZN(n549) );
  OAI21_X1 U1054 ( .B1(n548), .B2(n551), .A(n549), .ZN(n619) );
  INV_X1 U1055 ( .A(n619), .ZN(n557) );
  INV_X1 U1056 ( .A(operand_a_i[1]), .ZN(n2546) );
  MUX2_X1 U1057 ( .A(n74), .B(n2949), .S(n2546), .Z(n539) );
  OAI21_X1 U1058 ( .B1(n75), .B2(n538), .A(n539), .ZN(n543) );
  INV_X1 U1059 ( .A(n1181), .ZN(n1247) );
  MUX2_X1 U1060 ( .A(n1207), .B(n775), .S(operand_b_i[1]), .Z(n541) );
  NOR2_X1 U1062 ( .A1(n543), .A2(n542), .ZN(n614) );
  INV_X1 U1063 ( .A(n614), .ZN(n544) );
  NAND2_X1 U1065 ( .A1(n544), .A2(n616), .ZN(n545) );
  XOR2_X1 U1066 ( .A(n557), .B(n545), .Z(n3704) );
  INV_X1 U1068 ( .A(n2368), .ZN(n2358) );
  OAI21_X1 U1069 ( .B1(bmask_a_i[1]), .B2(bmask_b_i[0]), .A(n2358), .ZN(n735)
         );
  INV_X1 U1070 ( .A(bmask_a_i[2]), .ZN(n2348) );
  AND2_X1 U1071 ( .A1(n735), .A2(n2348), .ZN(n688) );
  NAND2_X1 U1072 ( .A1(n688), .A2(n729), .ZN(n1072) );
  NOR2_X1 U1073 ( .A1(bmask_a_i[4]), .A2(bmask_a_i[3]), .ZN(n732) );
  INV_X1 U1074 ( .A(n732), .ZN(n553) );
  INV_X1 U1075 ( .A(bmask_b_i[0]), .ZN(n719) );
  OAI22_X1 U1076 ( .A1(n1072), .A2(n553), .B1(n729), .B2(n719), .ZN(n1078) );
  OR2_X1 U1077 ( .A1(bmask_b_i[3]), .A2(bmask_b_i[2]), .ZN(n822) );
  OR2_X1 U1078 ( .A1(n1078), .A2(n822), .ZN(n741) );
  NOR2_X1 U1079 ( .A1(n741), .A2(bmask_b_i[4]), .ZN(n3456) );
  INV_X1 U1080 ( .A(n3456), .ZN(n547) );
  NAND2_X1 U1081 ( .A1(n2660), .A2(n2648), .ZN(n2662) );
  INV_X1 U1082 ( .A(n546), .ZN(n918) );
  NOR2_X1 U1083 ( .A1(n547), .A2(n546), .ZN(n555) );
  OR2_X1 U1084 ( .A1(n3704), .A2(n555), .ZN(n571) );
  INV_X1 U1085 ( .A(n548), .ZN(n550) );
  NAND2_X1 U1086 ( .A1(n550), .A2(n549), .ZN(n552) );
  XOR2_X1 U1087 ( .A(n552), .B(n551), .Z(n4176) );
  NOR2_X1 U1088 ( .A1(n2358), .A2(bmask_b_i[0]), .ZN(n753) );
  NAND2_X1 U1089 ( .A1(n753), .A2(n2348), .ZN(n711) );
  OAI21_X1 U1090 ( .B1(n711), .B2(n553), .A(n729), .ZN(n878) );
  NOR2_X1 U1091 ( .A1(n1218), .A2(bmask_b_i[2]), .ZN(n4120) );
  INV_X1 U1092 ( .A(n4120), .ZN(n1217) );
  NOR2_X1 U1093 ( .A1(n878), .A2(n1217), .ZN(n3715) );
  INV_X1 U1094 ( .A(n3715), .ZN(n554) );
  NOR2_X1 U1095 ( .A1(n554), .A2(n546), .ZN(n1262) );
  NAND2_X1 U1096 ( .A1(n4176), .A2(n1262), .ZN(n1263) );
  INV_X1 U1097 ( .A(n1263), .ZN(n572) );
  NAND2_X1 U1098 ( .A1(n3704), .A2(n555), .ZN(n570) );
  INV_X1 U1099 ( .A(n570), .ZN(n556) );
  AOI21_X1 U1100 ( .B1(n571), .B2(n572), .A(n556), .ZN(n944) );
  OAI21_X1 U1101 ( .B1(n557), .B2(n614), .A(n616), .ZN(n563) );
  INV_X1 U1103 ( .A(operand_a_i[2]), .ZN(n2547) );
  MUX2_X1 U1104 ( .A(n704), .B(n169), .S(n4087), .Z(n559) );
  OAI21_X1 U1105 ( .B1(n76), .B2(n71), .A(n559), .ZN(n612) );
  INV_X1 U1106 ( .A(n1181), .ZN(n817) );
  MUX2_X1 U1107 ( .A(n1207), .B(n1128), .S(operand_b_i[2]), .Z(n560) );
  NAND2_X1 U1108 ( .A1(n560), .A2(n458), .ZN(n613) );
  OR2_X1 U1109 ( .A1(n612), .A2(n613), .ZN(n561) );
  NAND2_X1 U1110 ( .A1(n612), .A2(n613), .ZN(n615) );
  NAND2_X1 U1111 ( .A1(n561), .A2(n615), .ZN(n562) );
  XNOR2_X1 U1112 ( .A(n563), .B(n562), .ZN(n3430) );
  OAI21_X1 U1113 ( .B1(n753), .B2(n729), .A(n732), .ZN(n564) );
  OR2_X1 U1114 ( .A1(bmask_a_i[0]), .A2(bmask_b_i[0]), .ZN(n718) );
  NAND2_X1 U1115 ( .A1(n718), .A2(bmask_a_i[1]), .ZN(n712) );
  NAND2_X1 U1116 ( .A1(n712), .A2(n2348), .ZN(n762) );
  NOR2_X1 U1117 ( .A1(n564), .A2(n762), .ZN(n1107) );
  NOR2_X1 U1118 ( .A1(n1107), .A2(n1217), .ZN(n3491) );
  INV_X1 U1119 ( .A(n3491), .ZN(n3462) );
  NOR2_X1 U1120 ( .A1(n3462), .A2(n546), .ZN(n565) );
  NOR2_X1 U1121 ( .A1(n3430), .A2(n565), .ZN(n943) );
  INV_X1 U1122 ( .A(n943), .ZN(n566) );
  NAND2_X1 U1123 ( .A1(n3430), .A2(n565), .ZN(n942) );
  NAND2_X1 U1124 ( .A1(n566), .A2(n942), .ZN(n567) );
  XOR2_X1 U1125 ( .A(n944), .B(n567), .Z(n569) );
  OAI22_X1 U1127 ( .A1(n1545), .A2(n4087), .B1(n1544), .B2(n53), .ZN(n568) );
  AOI21_X1 U1128 ( .B1(n569), .B2(n82), .A(n568), .ZN(n1766) );
  NAND2_X1 U1129 ( .A1(n571), .A2(n570), .ZN(n573) );
  XNOR2_X1 U1130 ( .A(n573), .B(n572), .ZN(n574) );
  NAND2_X1 U1131 ( .A1(n574), .A2(n82), .ZN(n577) );
  AOI22_X1 U1132 ( .A1(n1532), .A2(n4225), .B1(operand_a_i[30]), .B2(n91), 
        .ZN(n576) );
  NAND2_X1 U1133 ( .A1(n577), .A2(n576), .ZN(n1731) );
  INV_X1 U1134 ( .A(n1731), .ZN(n584) );
  INV_X1 U1135 ( .A(operand_b_i[0]), .ZN(n2661) );
  NAND2_X1 U1136 ( .A1(div_shift[0]), .A2(div_valid), .ZN(n578) );
  OAI21_X1 U1137 ( .B1(n2661), .B2(div_valid), .A(n578), .ZN(n1606) );
  INV_X1 U1138 ( .A(operand_b_i[16]), .ZN(n3765) );
  NAND2_X1 U1139 ( .A1(n1872), .A2(n4340), .ZN(n581) );
  OR2_X1 U1140 ( .A1(n579), .A2(n719), .ZN(n1589) );
  NAND3_X1 U1141 ( .A1(n82), .A2(is_clpx_i), .A3(clpx_shift_i[0]), .ZN(n580)
         );
  AND2_X1 U1142 ( .A1(n1589), .A2(n580), .ZN(n1601) );
  OAI211_X1 U1143 ( .C1(n3765), .C2(n582), .A(n581), .B(n1601), .ZN(n583) );
  AOI21_X1 U1144 ( .B1(n1606), .B2(n1871), .A(n583), .ZN(n1261) );
  MUX2_X1 U1145 ( .A(n1766), .B(n584), .S(n1657), .Z(n1408) );
  OR2_X1 U1146 ( .A1(n634), .A2(n2695), .ZN(n660) );
  MUX2_X1 U1147 ( .A(n704), .B(n2949), .S(n2543), .Z(n586) );
  OAI211_X1 U1149 ( .C1(n1207), .C2(operand_b_i[7]), .A(n589), .B(n470), .ZN(
        n632) );
  NOR2_X1 U1150 ( .A1(n633), .A2(n632), .ZN(n1008) );
  NOR2_X1 U1151 ( .A1(n635), .A2(n1008), .ZN(n995) );
  INV_X1 U1152 ( .A(operand_a_i[24]), .ZN(n3844) );
  INV_X1 U1153 ( .A(operand_a_i[8]), .ZN(n4106) );
  MUX2_X1 U1154 ( .A(n704), .B(n2949), .S(n4106), .Z(n590) );
  OAI21_X1 U1155 ( .B1(n75), .B2(n3844), .A(n590), .ZN(n636) );
  MUX2_X1 U1156 ( .A(n1247), .B(n775), .S(n4195), .Z(n594) );
  INV_X1 U1157 ( .A(operand_a_i[25]), .ZN(n3846) );
  MUX2_X1 U1158 ( .A(n169), .B(n704), .S(operand_a_i[9]), .Z(n595) );
  NAND2_X1 U1159 ( .A1(n995), .A2(n639), .ZN(n988) );
  INV_X1 U1160 ( .A(operand_a_i[26]), .ZN(n3848) );
  INV_X1 U1161 ( .A(operand_a_i[10]), .ZN(n2570) );
  MUX2_X1 U1162 ( .A(n1205), .B(n169), .S(n2570), .Z(n596) );
  OAI21_X1 U1163 ( .B1(n76), .B2(n3848), .A(n596), .ZN(n641) );
  MUX2_X1 U1164 ( .A(n1207), .B(n775), .S(operand_b_i[10]), .Z(n597) );
  OAI21_X1 U1165 ( .B1(n170), .B2(n83), .A(n597), .ZN(n640) );
  NOR2_X1 U1166 ( .A1(n641), .A2(n640), .ZN(n903) );
  MUX2_X1 U1167 ( .A(n2949), .B(n74), .S(operand_a_i[11]), .Z(n598) );
  OAI21_X1 U1168 ( .B1(n75), .B2(n2521), .A(n598), .ZN(n643) );
  MUX2_X1 U1169 ( .A(n775), .B(n1247), .S(n2562), .Z(n599) );
  NAND2_X1 U1170 ( .A1(n599), .A2(n469), .ZN(n642) );
  NOR2_X1 U1171 ( .A1(n903), .A2(n907), .ZN(n888) );
  INV_X1 U1173 ( .A(operand_a_i[12]), .ZN(n2561) );
  MUX2_X1 U1174 ( .A(n1205), .B(n2949), .S(n2561), .Z(n600) );
  OAI21_X1 U1175 ( .B1(n76), .B2(n2522), .A(n600), .ZN(n645) );
  MUX2_X1 U1176 ( .A(n1247), .B(n1128), .S(operand_b_i[12]), .Z(n601) );
  NAND2_X1 U1177 ( .A1(n601), .A2(n473), .ZN(n644) );
  MUX2_X1 U1178 ( .A(n1207), .B(n1128), .S(operand_b_i[13]), .Z(n602) );
  NAND2_X1 U1179 ( .A1(n602), .A2(n466), .ZN(n646) );
  MUX2_X1 U1180 ( .A(n704), .B(n2949), .S(n4101), .Z(n603) );
  OAI21_X1 U1181 ( .B1(n75), .B2(n53), .A(n603), .ZN(n647) );
  NOR2_X1 U1182 ( .A1(n923), .A2(n897), .ZN(n649) );
  NOR2_X1 U1184 ( .A1(n988), .A2(n651), .ZN(n653) );
  INV_X1 U1185 ( .A(operand_a_i[19]), .ZN(n4105) );
  MUX2_X1 U1186 ( .A(n169), .B(n1205), .S(n48), .Z(n604) );
  OAI21_X1 U1187 ( .B1(n75), .B2(n4105), .A(n604), .ZN(n622) );
  MUX2_X1 U1188 ( .A(n817), .B(n775), .S(operand_b_i[3]), .Z(n605) );
  OAI21_X1 U1189 ( .B1(operand_b_i[19]), .B2(n83), .A(n605), .ZN(n621) );
  NOR2_X1 U1190 ( .A1(n622), .A2(n621), .ZN(n931) );
  INV_X1 U1191 ( .A(operand_a_i[20]), .ZN(n4067) );
  INV_X1 U1192 ( .A(operand_a_i[4]), .ZN(n4108) );
  OAI21_X1 U1193 ( .B1(n75), .B2(n4067), .A(n606), .ZN(n624) );
  INV_X1 U1194 ( .A(operand_b_i[4]), .ZN(n3812) );
  MUX2_X1 U1195 ( .A(n1128), .B(n1247), .S(n3812), .Z(n607) );
  NAND2_X1 U1196 ( .A1(n607), .A2(n468), .ZN(n623) );
  INV_X1 U1198 ( .A(operand_a_i[5]), .ZN(n4079) );
  MUX2_X1 U1199 ( .A(n1205), .B(n2949), .S(n4079), .Z(n608) );
  OAI21_X1 U1200 ( .B1(n76), .B2(n4075), .A(n608), .ZN(n626) );
  MUX2_X1 U1201 ( .A(n817), .B(n775), .S(operand_b_i[5]), .Z(n609) );
  OAI21_X1 U1202 ( .B1(operand_b_i[21]), .B2(n83), .A(n609), .ZN(n625) );
  MUX2_X1 U1204 ( .A(n1207), .B(n775), .S(operand_b_i[6]), .Z(n610) );
  NAND2_X1 U1205 ( .A1(n610), .A2(n474), .ZN(n627) );
  INV_X1 U1206 ( .A(operand_a_i[22]), .ZN(n2514) );
  INV_X1 U1207 ( .A(operand_a_i[6]), .ZN(n2553) );
  MUX2_X1 U1208 ( .A(n74), .B(n169), .S(n4071), .Z(n611) );
  OAI21_X1 U1209 ( .B1(n75), .B2(n4072), .A(n611), .ZN(n628) );
  NOR2_X1 U1210 ( .A1(n950), .A2(n956), .ZN(n630) );
  NOR2_X1 U1211 ( .A1(n612), .A2(n613), .ZN(n617) );
  NOR2_X1 U1212 ( .A1(n614), .A2(n617), .ZN(n620) );
  OAI21_X1 U1213 ( .B1(n617), .B2(n616), .A(n615), .ZN(n618) );
  AOI21_X1 U1214 ( .B1(n620), .B2(n619), .A(n618), .ZN(n930) );
  NAND2_X1 U1215 ( .A1(n622), .A2(n621), .ZN(n937) );
  NAND2_X1 U1216 ( .A1(n624), .A2(n623), .ZN(n934) );
  OAI21_X1 U1217 ( .B1(n933), .B2(n937), .A(n934), .ZN(n952) );
  NAND2_X1 U1218 ( .A1(n626), .A2(n625), .ZN(n965) );
  NAND2_X1 U1219 ( .A1(n628), .A2(n627), .ZN(n957) );
  OAI21_X1 U1220 ( .B1(n956), .B2(n965), .A(n957), .ZN(n629) );
  AOI21_X1 U1221 ( .B1(n630), .B2(n952), .A(n629), .ZN(n631) );
  AND2_X1 U1222 ( .A1(n634), .A2(vector_mode_i[1]), .ZN(n669) );
  NAND2_X1 U1223 ( .A1(n638), .A2(n637), .ZN(n980) );
  NAND2_X1 U1224 ( .A1(n641), .A2(n640), .ZN(n989) );
  NAND2_X1 U1225 ( .A1(n643), .A2(n642), .ZN(n908) );
  OAI21_X1 U1226 ( .B1(n907), .B2(n989), .A(n908), .ZN(n891) );
  NAND2_X1 U1227 ( .A1(n645), .A2(n644), .ZN(n924) );
  NAND2_X1 U1228 ( .A1(n647), .A2(n646), .ZN(n898) );
  OAI21_X1 U1229 ( .B1(n897), .B2(n924), .A(n898), .ZN(n648) );
  AOI21_X1 U1230 ( .B1(n649), .B2(n891), .A(n648), .ZN(n650) );
  OAI21_X1 U1231 ( .B1(n890), .B2(n651), .A(n650), .ZN(n652) );
  INV_X1 U1233 ( .A(operand_a_i[30]), .ZN(n4112) );
  INV_X1 U1234 ( .A(operand_a_i[14]), .ZN(n4098) );
  OAI21_X1 U1235 ( .B1(n76), .B2(n4112), .A(n654), .ZN(n665) );
  MUX2_X1 U1236 ( .A(n1247), .B(n775), .S(operand_b_i[14]), .Z(n655) );
  NAND2_X1 U1237 ( .A1(n655), .A2(n467), .ZN(n666) );
  NOR2_X1 U1238 ( .A1(n665), .A2(n65), .ZN(n856) );
  MUX2_X1 U1239 ( .A(n1207), .B(n775), .S(operand_b_i[15]), .Z(n656) );
  NAND2_X1 U1240 ( .A1(n656), .A2(n471), .ZN(n667) );
  INV_X1 U1242 ( .A(operand_a_i[15]), .ZN(n4095) );
  MUX2_X1 U1243 ( .A(n74), .B(n2949), .S(n4095), .Z(n657) );
  OAI21_X1 U1244 ( .B1(n76), .B2(n4115), .A(n657), .ZN(n668) );
  NOR2_X1 U1245 ( .A1(n856), .A2(n858), .ZN(n864) );
  MUX2_X1 U1246 ( .A(n775), .B(n1247), .S(n3765), .Z(n658) );
  NAND2_X1 U1247 ( .A1(n658), .A2(n450), .ZN(n670) );
  MUX2_X1 U1248 ( .A(n2949), .B(n74), .S(operand_a_i[16]), .Z(n659) );
  OAI21_X1 U1249 ( .B1(n76), .B2(n2661), .A(n659), .ZN(n671) );
  INV_X1 U1250 ( .A(n660), .ZN(n868) );
  NAND2_X1 U1251 ( .A1(n864), .A2(n672), .ZN(n771) );
  INV_X1 U1252 ( .A(n771), .ZN(n726) );
  MUX2_X1 U1253 ( .A(n2949), .B(n1205), .S(operand_a_i[17]), .Z(n661) );
  OAI21_X1 U1254 ( .B1(n75), .B2(n2464), .A(n661), .ZN(n674) );
  MUX2_X1 U1255 ( .A(n1207), .B(n775), .S(operand_b_i[17]), .Z(n662) );
  OAI21_X1 U1256 ( .B1(n4225), .B2(n83), .A(n662), .ZN(n673) );
  NOR2_X1 U1257 ( .A1(n674), .A2(n673), .ZN(n745) );
  MUX2_X1 U1258 ( .A(n1205), .B(n169), .S(n71), .Z(n663) );
  OAI21_X1 U1259 ( .B1(n76), .B2(n3438), .A(n663), .ZN(n676) );
  MUX2_X1 U1260 ( .A(n1247), .B(n775), .S(n4194), .Z(n664) );
  OAI21_X1 U1261 ( .B1(operand_a_i[2]), .B2(n83), .A(n664), .ZN(n675) );
  NOR2_X1 U1262 ( .A1(n676), .A2(n675), .ZN(n748) );
  NAND2_X1 U1263 ( .A1(n726), .A2(n770), .ZN(n700) );
  INV_X1 U1264 ( .A(n700), .ZN(n678) );
  NAND2_X1 U1265 ( .A1(n666), .A2(n665), .ZN(n885) );
  NAND2_X1 U1266 ( .A1(n668), .A2(n667), .ZN(n859) );
  INV_X1 U1267 ( .A(n669), .ZN(n867) );
  NAND2_X1 U1268 ( .A1(n671), .A2(n670), .ZN(n873) );
  INV_X1 U1269 ( .A(n783), .ZN(n725) );
  NAND2_X1 U1270 ( .A1(n674), .A2(n673), .ZN(n744) );
  NAND2_X1 U1271 ( .A1(n676), .A2(n675), .ZN(n749) );
  OAI21_X1 U1272 ( .B1(n748), .B2(n744), .A(n749), .ZN(n781) );
  AOI21_X1 U1273 ( .B1(n725), .B2(n770), .A(n781), .ZN(n701) );
  INV_X1 U1274 ( .A(n701), .ZN(n677) );
  AOI21_X1 U1275 ( .B1(n4291), .B2(n678), .A(n677), .ZN(n686) );
  MUX2_X1 U1276 ( .A(n74), .B(n169), .S(n4105), .Z(n680) );
  OAI21_X1 U1277 ( .B1(n76), .B2(n3479), .A(n680), .ZN(n683) );
  MUX2_X1 U1278 ( .A(n1247), .B(n775), .S(operand_b_i[19]), .Z(n681) );
  OAI21_X1 U1279 ( .B1(n48), .B2(n83), .A(n681), .ZN(n682) );
  NOR2_X1 U1280 ( .A1(n683), .A2(n682), .ZN(n769) );
  INV_X1 U1281 ( .A(n769), .ZN(n684) );
  NAND2_X1 U1282 ( .A1(n683), .A2(n682), .ZN(n778) );
  NAND2_X1 U1283 ( .A1(n711), .A2(bmask_a_i[3]), .ZN(n720) );
  OR2_X1 U1284 ( .A1(n720), .A2(n729), .ZN(n764) );
  INV_X1 U1285 ( .A(n2372), .ZN(n2347) );
  NOR2_X1 U1286 ( .A1(n2347), .A2(n719), .ZN(n731) );
  AND2_X1 U1287 ( .A1(bmask_a_i[3]), .A2(bmask_a_i[2]), .ZN(n2342) );
  AOI21_X1 U1288 ( .B1(n731), .B2(bmask_a_i[3]), .A(n2342), .ZN(n687) );
  OAI21_X1 U1289 ( .B1(n764), .B2(n688), .A(n687), .ZN(n1135) );
  OR2_X1 U1290 ( .A1(n1135), .A2(bmask_a_i[4]), .ZN(n799) );
  INV_X1 U1291 ( .A(n731), .ZN(n738) );
  AOI21_X1 U1292 ( .B1(n729), .B2(n738), .A(n735), .ZN(n694) );
  AND2_X1 U1293 ( .A1(n694), .A2(bmask_a_i[2]), .ZN(n692) );
  INV_X1 U1294 ( .A(n692), .ZN(n689) );
  INV_X1 U1295 ( .A(bmask_a_i[3]), .ZN(n2345) );
  AND2_X1 U1296 ( .A1(n689), .A2(n2345), .ZN(n805) );
  NOR2_X1 U1297 ( .A1(n805), .A2(n1076), .ZN(n690) );
  NOR2_X1 U1298 ( .A1(n799), .A2(n690), .ZN(n912) );
  INV_X1 U1299 ( .A(n720), .ZN(n691) );
  AOI21_X1 U1300 ( .B1(n692), .B2(n691), .A(bmask_a_i[4]), .ZN(n800) );
  NOR2_X1 U1301 ( .A1(bmask_a_i[3]), .A2(bmask_a_i[2]), .ZN(n2352) );
  INV_X1 U1302 ( .A(n2352), .ZN(n693) );
  OAI21_X1 U1303 ( .B1(n694), .B2(n693), .A(bmask_a_i[4]), .ZN(n803) );
  OAI21_X1 U1304 ( .B1(n800), .B2(n1076), .A(n803), .ZN(n1139) );
  INV_X1 U1305 ( .A(n694), .ZN(n695) );
  NAND3_X1 U1306 ( .A1(n695), .A2(n732), .A3(n2348), .ZN(n914) );
  NOR2_X1 U1307 ( .A1(bmask_b_i[1]), .A2(bmask_b_i[0]), .ZN(n4119) );
  AND2_X1 U1308 ( .A1(n4119), .A2(bmask_b_i[2]), .ZN(n696) );
  AOI21_X1 U1309 ( .B1(n914), .B2(n1076), .A(n696), .ZN(n940) );
  AND2_X1 U1310 ( .A1(bmask_b_i[3]), .A2(bmask_b_i[4]), .ZN(n1173) );
  AOI21_X1 U1311 ( .B1(n940), .B2(bmask_b_i[4]), .A(n1173), .ZN(n697) );
  OAI21_X1 U1312 ( .B1(n1139), .B2(n1218), .A(n697), .ZN(n698) );
  AOI21_X1 U1313 ( .B1(bmask_b_i[3]), .B2(n912), .A(n698), .ZN(n3919) );
  INV_X1 U1314 ( .A(n3919), .ZN(n699) );
  NOR2_X1 U1316 ( .A1(n699), .A2(n1223), .ZN(n1045) );
  NOR2_X1 U1317 ( .A1(n700), .A2(n769), .ZN(n703) );
  OAI21_X1 U1318 ( .B1(n701), .B2(n769), .A(n778), .ZN(n702) );
  AOI21_X1 U1319 ( .B1(n1126), .B2(n703), .A(n702), .ZN(n710) );
  MUX2_X1 U1320 ( .A(n704), .B(n169), .S(n4067), .Z(n705) );
  OAI21_X1 U1321 ( .B1(n75), .B2(n3812), .A(n705), .ZN(n708) );
  MUX2_X1 U1322 ( .A(n1207), .B(n775), .S(operand_b_i[20]), .Z(n706) );
  OAI21_X1 U1323 ( .B1(operand_a_i[4]), .B2(n83), .A(n706), .ZN(n707) );
  INV_X1 U1324 ( .A(n779), .ZN(n709) );
  NAND2_X1 U1325 ( .A1(n708), .A2(n707), .ZN(n777) );
  XNOR2_X1 U1326 ( .A(n710), .B(n454), .ZN(n3922) );
  OR2_X1 U1327 ( .A1(n711), .A2(bmask_a_i[3]), .ZN(n757) );
  OAI21_X1 U1328 ( .B1(n757), .B2(bmask_b_i[1]), .A(bmask_a_i[4]), .ZN(n714)
         );
  INV_X1 U1329 ( .A(n2342), .ZN(n2356) );
  NOR2_X1 U1330 ( .A1(n2356), .A2(n712), .ZN(n755) );
  NAND2_X1 U1331 ( .A1(n755), .A2(bmask_b_i[1]), .ZN(n713) );
  AND2_X1 U1332 ( .A1(n714), .A2(n713), .ZN(n879) );
  AOI22_X1 U1333 ( .A1(n4119), .A2(n2368), .B1(n729), .B2(n2348), .ZN(n715) );
  NAND2_X1 U1334 ( .A1(n762), .A2(n715), .ZN(n722) );
  AND2_X1 U1335 ( .A1(n722), .A2(n2345), .ZN(n716) );
  OR2_X1 U1336 ( .A1(n716), .A2(n2369), .ZN(n827) );
  OAI21_X1 U1337 ( .B1(n879), .B2(n1076), .A(n827), .ZN(n1177) );
  NAND2_X1 U1338 ( .A1(n716), .A2(n2369), .ZN(n1004) );
  NAND2_X1 U1339 ( .A1(n878), .A2(bmask_b_i[2]), .ZN(n717) );
  OAI21_X1 U1340 ( .B1(n1004), .B2(bmask_b_i[2]), .A(n717), .ZN(n1174) );
  AOI21_X1 U1341 ( .B1(n1174), .B2(bmask_b_i[4]), .A(n1173), .ZN(n724) );
  AND2_X1 U1342 ( .A1(bmask_a_i[1]), .A2(bmask_a_i[2]), .ZN(n759) );
  AOI21_X1 U1343 ( .B1(n759), .B2(n718), .A(bmask_a_i[3]), .ZN(n721) );
  OAI21_X1 U1344 ( .B1(n759), .B2(n719), .A(bmask_b_i[1]), .ZN(n733) );
  OAI21_X1 U1345 ( .B1(n721), .B2(n733), .A(n720), .ZN(n1168) );
  NOR2_X1 U1346 ( .A1(n1168), .A2(bmask_a_i[4]), .ZN(n880) );
  NOR2_X1 U1347 ( .A1(n722), .A2(n2345), .ZN(n1169) );
  NOR2_X1 U1348 ( .A1(n1169), .A2(bmask_a_i[4]), .ZN(n877) );
  OAI21_X1 U1349 ( .B1(n880), .B2(n1076), .A(n877), .ZN(n928) );
  OR2_X1 U1350 ( .A1(n928), .A2(n1109), .ZN(n723) );
  OAI211_X1 U1351 ( .C1(n1177), .C2(n1218), .A(n724), .B(n723), .ZN(n3270) );
  NOR2_X1 U1352 ( .A1(n3270), .A2(n1223), .ZN(n1046) );
  NOR2_X1 U1353 ( .A1(n1382), .A2(n1388), .ZN(n1048) );
  AOI21_X1 U1354 ( .B1(n1126), .B2(n726), .A(n725), .ZN(n728) );
  INV_X1 U1355 ( .A(n745), .ZN(n727) );
  XNOR2_X1 U1356 ( .A(n728), .B(n445), .ZN(n2987) );
  OAI21_X1 U1357 ( .B1(n735), .B2(n2348), .A(n729), .ZN(n730) );
  OAI21_X1 U1358 ( .B1(n731), .B2(bmask_a_i[2]), .A(n730), .ZN(n1190) );
  AND2_X1 U1359 ( .A1(n1190), .A2(n732), .ZN(n1083) );
  OAI21_X1 U1360 ( .B1(n738), .B2(n733), .A(n2345), .ZN(n1073) );
  AOI21_X1 U1361 ( .B1(n1073), .B2(n1072), .A(bmask_a_i[4]), .ZN(n1080) );
  OAI21_X1 U1362 ( .B1(n1083), .B2(n1076), .A(n1080), .ZN(n986) );
  NAND2_X1 U1363 ( .A1(n2342), .A2(bmask_b_i[1]), .ZN(n739) );
  OR2_X1 U1364 ( .A1(bmask_b_i[1]), .A2(bmask_a_i[3]), .ZN(n734) );
  OR2_X1 U1365 ( .A1(n762), .A2(n734), .ZN(n758) );
  INV_X1 U1366 ( .A(n735), .ZN(n736) );
  OAI21_X1 U1367 ( .B1(n758), .B2(n736), .A(bmask_a_i[4]), .ZN(n737) );
  OAI21_X1 U1368 ( .B1(n739), .B2(n738), .A(n737), .ZN(n1075) );
  OAI21_X1 U1369 ( .B1(n1190), .B2(n2345), .A(n2369), .ZN(n1081) );
  OR2_X1 U1370 ( .A1(n1076), .A2(bmask_b_i[3]), .ZN(n823) );
  OAI22_X1 U1371 ( .A1(n1075), .A2(n1217), .B1(n1081), .B2(n823), .ZN(n740) );
  INV_X1 U1372 ( .A(n740), .ZN(n743) );
  NAND2_X1 U1373 ( .A1(n741), .A2(bmask_b_i[4]), .ZN(n742) );
  OAI211_X1 U1374 ( .C1(n986), .C2(n1109), .A(n743), .B(n742), .ZN(n3174) );
  NOR2_X1 U1375 ( .A1(n3174), .A2(n546), .ZN(n1042) );
  NOR2_X1 U1376 ( .A1(n2987), .A2(n1042), .ZN(n1377) );
  NOR2_X1 U1377 ( .A1(n771), .A2(n745), .ZN(n747) );
  OAI21_X1 U1378 ( .B1(n783), .B2(n745), .A(n744), .ZN(n746) );
  AOI21_X1 U1379 ( .B1(n1126), .B2(n747), .A(n746), .ZN(n751) );
  INV_X1 U1380 ( .A(n748), .ZN(n750) );
  XNOR2_X1 U1381 ( .A(n751), .B(n453), .ZN(n1043) );
  OAI21_X1 U1382 ( .B1(bmask_a_i[1]), .B2(bmask_b_i[1]), .A(bmask_a_i[2]), 
        .ZN(n752) );
  OR2_X1 U1383 ( .A1(n4119), .A2(n752), .ZN(n754) );
  OR2_X1 U1384 ( .A1(n754), .A2(n753), .ZN(n761) );
  INV_X1 U1385 ( .A(n755), .ZN(n756) );
  OAI21_X1 U1386 ( .B1(n764), .B2(n761), .A(n756), .ZN(n1216) );
  NOR2_X1 U1387 ( .A1(n1216), .A2(bmask_a_i[4]), .ZN(n848) );
  NAND3_X1 U1388 ( .A1(n758), .A2(bmask_a_i[4]), .A3(n757), .ZN(n851) );
  OAI21_X1 U1389 ( .B1(n848), .B2(n1076), .A(n851), .ZN(n1114) );
  NAND2_X1 U1390 ( .A1(n1114), .A2(n1171), .ZN(n767) );
  AOI21_X1 U1391 ( .B1(n759), .B2(bmask_a_i[0]), .A(bmask_a_i[3]), .ZN(n760)
         );
  AND2_X1 U1392 ( .A1(n761), .A2(n760), .ZN(n849) );
  NAND2_X1 U1393 ( .A1(n762), .A2(bmask_a_i[3]), .ZN(n763) );
  AND2_X1 U1394 ( .A1(n764), .A2(n763), .ZN(n1104) );
  OAI211_X1 U1395 ( .C1(n849), .C2(n1076), .A(n1104), .B(n2369), .ZN(n1110) );
  OR2_X1 U1396 ( .A1(n1109), .A2(bmask_b_i[4]), .ZN(n1214) );
  INV_X1 U1397 ( .A(n1214), .ZN(n1193) );
  NOR2_X1 U1398 ( .A1(n822), .A2(n1196), .ZN(n1079) );
  INV_X1 U1399 ( .A(n1107), .ZN(n765) );
  AOI22_X1 U1400 ( .A1(n1110), .A2(n1193), .B1(n1079), .B2(n765), .ZN(n766) );
  NAND2_X1 U1401 ( .A1(n767), .A2(n766), .ZN(n3026) );
  INV_X1 U1402 ( .A(n3026), .ZN(n768) );
  NOR2_X1 U1403 ( .A1(n768), .A2(n1223), .ZN(n1044) );
  NAND2_X1 U1404 ( .A1(n1392), .A2(n1048), .ZN(n1335) );
  NOR2_X1 U1405 ( .A1(n769), .A2(n779), .ZN(n782) );
  NOR2_X1 U1406 ( .A1(n784), .A2(n771), .ZN(n1147) );
  INV_X1 U1407 ( .A(n1147), .ZN(n1116) );
  INV_X1 U1408 ( .A(operand_b_i[5]), .ZN(n3738) );
  MUX2_X1 U1409 ( .A(n74), .B(n2949), .S(n4075), .Z(n772) );
  OAI21_X1 U1410 ( .B1(n75), .B2(n3738), .A(n772), .ZN(n786) );
  MUX2_X1 U1411 ( .A(n1247), .B(n1128), .S(operand_b_i[21]), .Z(n773) );
  OAI21_X1 U1412 ( .B1(operand_a_i[5]), .B2(n83), .A(n773), .ZN(n785) );
  NOR2_X1 U1413 ( .A1(n786), .A2(n785), .ZN(n841) );
  INV_X1 U1414 ( .A(operand_b_i[6]), .ZN(n3663) );
  MUX2_X1 U1415 ( .A(n1205), .B(n169), .S(n4072), .Z(n774) );
  OAI21_X1 U1416 ( .B1(n75), .B2(n3663), .A(n774), .ZN(n788) );
  MUX2_X1 U1417 ( .A(n1207), .B(n1128), .S(operand_b_i[22]), .Z(n776) );
  OAI21_X1 U1418 ( .B1(operand_a_i[6]), .B2(n83), .A(n776), .ZN(n787) );
  NOR2_X1 U1419 ( .A1(n788), .A2(n787), .ZN(n844) );
  NOR2_X1 U1420 ( .A1(n841), .A2(n844), .ZN(n809) );
  INV_X1 U1421 ( .A(n809), .ZN(n790) );
  NOR2_X1 U1422 ( .A1(n1116), .A2(n790), .ZN(n792) );
  OAI21_X1 U1423 ( .B1(n779), .B2(n778), .A(n777), .ZN(n780) );
  NAND2_X1 U1424 ( .A1(n786), .A2(n785), .ZN(n840) );
  NAND2_X1 U1425 ( .A1(n788), .A2(n787), .ZN(n845) );
  OAI21_X1 U1426 ( .B1(n844), .B2(n840), .A(n845), .ZN(n812) );
  INV_X1 U1427 ( .A(n812), .ZN(n789) );
  OAI21_X1 U1428 ( .B1(n1123), .B2(n790), .A(n789), .ZN(n791) );
  AOI21_X1 U1429 ( .B1(n1126), .B2(n792), .A(n791), .ZN(n798) );
  MUX2_X1 U1430 ( .A(n1205), .B(n169), .S(n585), .Z(n793) );
  OAI21_X1 U1431 ( .B1(n76), .B2(n588), .A(n793), .ZN(n796) );
  MUX2_X1 U1432 ( .A(n817), .B(n1128), .S(operand_b_i[23]), .Z(n794) );
  OAI21_X1 U1433 ( .B1(operand_a_i[7]), .B2(n83), .A(n794), .ZN(n795) );
  NOR2_X1 U1434 ( .A1(n796), .A2(n795), .ZN(n808) );
  INV_X1 U1435 ( .A(n808), .ZN(n797) );
  NAND2_X1 U1436 ( .A1(n796), .A2(n795), .ZN(n810) );
  XNOR2_X1 U1437 ( .A(n798), .B(n449), .ZN(n2952) );
  NAND2_X1 U1438 ( .A1(n799), .A2(bmask_b_i[2]), .ZN(n801) );
  NAND2_X1 U1439 ( .A1(n801), .A2(n800), .ZN(n863) );
  INV_X1 U1440 ( .A(n805), .ZN(n802) );
  NAND2_X1 U1441 ( .A1(n802), .A2(bmask_a_i[4]), .ZN(n1136) );
  AOI22_X1 U1442 ( .A1(n1136), .A2(n4120), .B1(n1171), .B2(n803), .ZN(n807) );
  AOI21_X1 U1443 ( .B1(n914), .B2(bmask_b_i[2]), .A(bmask_a_i[4]), .ZN(n804)
         );
  AND2_X1 U1444 ( .A1(n805), .A2(n804), .ZN(n1013) );
  NOR2_X1 U1445 ( .A1(n1109), .A2(bmask_b_i[2]), .ZN(n984) );
  NAND2_X1 U1446 ( .A1(n984), .A2(n4119), .ZN(n1012) );
  OAI211_X1 U1447 ( .C1(n1013), .C2(bmask_b_i[3]), .A(bmask_b_i[4]), .B(n1012), 
        .ZN(n806) );
  OAI211_X1 U1448 ( .C1(n863), .C2(n1214), .A(n807), .B(n806), .ZN(n3552) );
  NOR2_X1 U1449 ( .A1(n3552), .A2(n1223), .ZN(n1052) );
  NOR2_X1 U1450 ( .A1(n635), .A2(n808), .ZN(n813) );
  NAND2_X1 U1451 ( .A1(n813), .A2(n809), .ZN(n1146) );
  NOR2_X1 U1452 ( .A1(n1116), .A2(n1146), .ZN(n815) );
  OAI21_X1 U1453 ( .B1(n635), .B2(n810), .A(n174), .ZN(n811) );
  AOI21_X1 U1454 ( .B1(n813), .B2(n812), .A(n811), .ZN(n1156) );
  AOI21_X1 U1455 ( .B1(n1126), .B2(n815), .A(n814), .ZN(n821) );
  MUX2_X1 U1456 ( .A(n2949), .B(n1205), .S(operand_a_i[24]), .Z(n816) );
  OAI21_X1 U1457 ( .B1(n76), .B2(n2566), .A(n816), .ZN(n820) );
  MUX2_X1 U1458 ( .A(n1247), .B(n1128), .S(n4340), .Z(n818) );
  OAI21_X1 U1459 ( .B1(n149), .B2(n540), .A(n818), .ZN(n819) );
  NOR2_X1 U1460 ( .A1(n820), .A2(n819), .ZN(n1089) );
  INV_X1 U1461 ( .A(n1089), .ZN(n1061) );
  NAND2_X1 U1462 ( .A1(n820), .A2(n819), .ZN(n1091) );
  XNOR2_X1 U1463 ( .A(n821), .B(n446), .ZN(n3542) );
  INV_X1 U1464 ( .A(n984), .ZN(n1106) );
  OAI22_X1 U1465 ( .A1(n880), .A2(n822), .B1(n878), .B2(n1106), .ZN(n1003) );
  INV_X1 U1466 ( .A(n823), .ZN(n824) );
  NAND2_X1 U1467 ( .A1(n1004), .A2(n824), .ZN(n825) );
  NAND2_X1 U1468 ( .A1(n825), .A2(bmask_b_i[4]), .ZN(n830) );
  INV_X1 U1469 ( .A(n1168), .ZN(n826) );
  AOI22_X1 U1470 ( .A1(n1171), .A2(n827), .B1(n826), .B2(n4120), .ZN(n829) );
  OAI211_X1 U1471 ( .C1(n877), .C2(n1076), .A(n879), .B(n1193), .ZN(n828) );
  OAI211_X1 U1472 ( .C1(n1003), .C2(n830), .A(n829), .B(n828), .ZN(n4018) );
  NOR2_X1 U1473 ( .A1(n4018), .A2(n1223), .ZN(n1053) );
  NOR2_X1 U1474 ( .A1(n3542), .A2(n1053), .ZN(n1349) );
  NOR2_X1 U1475 ( .A1(n1359), .A2(n1349), .ZN(n1055) );
  AOI21_X1 U1476 ( .B1(n4291), .B2(n1147), .A(n4308), .ZN(n832) );
  INV_X1 U1477 ( .A(n841), .ZN(n831) );
  AOI21_X1 U1478 ( .B1(n1190), .B2(n2345), .A(n2369), .ZN(n1084) );
  AOI21_X1 U1479 ( .B1(n1075), .B2(bmask_b_i[2]), .A(n1084), .ZN(n1194) );
  NAND2_X1 U1480 ( .A1(n1078), .A2(bmask_b_i[2]), .ZN(n834) );
  NAND2_X1 U1481 ( .A1(n1083), .A2(n1076), .ZN(n833) );
  AND2_X1 U1482 ( .A1(n834), .A2(n833), .ZN(n969) );
  INV_X1 U1483 ( .A(n969), .ZN(n835) );
  MUX2_X1 U1484 ( .A(n1194), .B(n835), .S(bmask_b_i[4]), .Z(n838) );
  INV_X1 U1485 ( .A(n1081), .ZN(n836) );
  OAI21_X1 U1486 ( .B1(n1080), .B2(n1076), .A(n836), .ZN(n902) );
  NAND2_X1 U1487 ( .A1(n902), .A2(n1193), .ZN(n837) );
  OAI21_X1 U1488 ( .B1(n838), .B2(bmask_b_i[3]), .A(n837), .ZN(n3131) );
  INV_X1 U1489 ( .A(n3131), .ZN(n839) );
  NOR2_X1 U1490 ( .A1(n839), .A2(n1223), .ZN(n1049) );
  NOR2_X1 U1491 ( .A1(n3274), .A2(n1049), .ZN(n1324) );
  NOR2_X1 U1492 ( .A1(n1116), .A2(n841), .ZN(n843) );
  OAI21_X1 U1493 ( .B1(n1123), .B2(n841), .A(n840), .ZN(n842) );
  AOI21_X1 U1494 ( .B1(n1126), .B2(n843), .A(n842), .ZN(n847) );
  INV_X1 U1495 ( .A(n844), .ZN(n846) );
  XNOR2_X1 U1496 ( .A(n847), .B(n444), .ZN(n1050) );
  OAI21_X1 U1497 ( .B1(n1104), .B2(n1076), .A(n848), .ZN(n887) );
  NAND2_X1 U1498 ( .A1(n887), .A2(n1196), .ZN(n854) );
  OAI211_X1 U1499 ( .C1(n1107), .C2(n1076), .A(n849), .B(n2369), .ZN(n961) );
  NAND2_X1 U1500 ( .A1(n961), .A2(n1109), .ZN(n853) );
  NOR2_X1 U1501 ( .A1(n849), .A2(n2369), .ZN(n1105) );
  INV_X1 U1502 ( .A(n1105), .ZN(n850) );
  OAI21_X1 U1503 ( .B1(n851), .B2(n1076), .A(n850), .ZN(n1215) );
  NOR2_X1 U1504 ( .A1(n1215), .A2(n1218), .ZN(n852) );
  AOI21_X1 U1505 ( .B1(n854), .B2(n853), .A(n852), .ZN(n2946) );
  INV_X1 U1506 ( .A(n2946), .ZN(n855) );
  NOR2_X1 U1507 ( .A1(n855), .A2(n1223), .ZN(n1051) );
  NAND2_X1 U1508 ( .A1(n1055), .A2(n1341), .ZN(n1057) );
  NOR2_X1 U1509 ( .A1(n1335), .A2(n1057), .ZN(n1059) );
  INV_X1 U1510 ( .A(n856), .ZN(n886) );
  INV_X1 U1511 ( .A(n885), .ZN(n857) );
  AOI21_X1 U1512 ( .B1(n4291), .B2(n886), .A(n857), .ZN(n861) );
  INV_X1 U1513 ( .A(n858), .ZN(n860) );
  INV_X1 U1514 ( .A(n1013), .ZN(n862) );
  AOI222_X1 U1515 ( .A1(n863), .A2(n1171), .B1(n4119), .B2(n1079), .C1(n862), 
        .C2(n1193), .ZN(n3767) );
  NOR2_X1 U1516 ( .A1(n3767), .A2(n546), .ZN(n1026) );
  INV_X1 U1517 ( .A(n864), .ZN(n865) );
  NOR2_X1 U1518 ( .A1(n865), .A2(n868), .ZN(n871) );
  INV_X1 U1519 ( .A(n866), .ZN(n869) );
  OAI21_X1 U1520 ( .B1(n869), .B2(n868), .A(n867), .ZN(n870) );
  AOI21_X1 U1521 ( .B1(n4291), .B2(n871), .A(n870), .ZN(n875) );
  INV_X1 U1522 ( .A(n872), .ZN(n874) );
  NAND2_X1 U1523 ( .A1(n1004), .A2(bmask_b_i[3]), .ZN(n876) );
  OAI211_X1 U1524 ( .C1(n877), .C2(n1218), .A(n876), .B(bmask_b_i[2]), .ZN(
        n884) );
  AOI21_X1 U1525 ( .B1(n878), .B2(bmask_b_i[4]), .A(n1173), .ZN(n883) );
  NAND2_X1 U1526 ( .A1(n879), .A2(n4120), .ZN(n882) );
  NAND2_X1 U1527 ( .A1(n880), .A2(n984), .ZN(n881) );
  NOR2_X1 U1529 ( .A1(n3000), .A2(n546), .ZN(n1027) );
  NOR2_X1 U1530 ( .A1(n3779), .A2(n1027), .ZN(n1484) );
  NOR2_X1 U1531 ( .A1(n1493), .A2(n1484), .ZN(n1038) );
  OAI21_X1 U1532 ( .B1(n887), .B2(bmask_b_i[3]), .A(n961), .ZN(n1222) );
  OR2_X1 U1533 ( .A1(n1222), .A2(bmask_b_i[4]), .ZN(n3066) );
  NOR2_X1 U1534 ( .A1(n3066), .A2(n546), .ZN(n1033) );
  INV_X1 U1535 ( .A(n888), .ZN(n889) );
  NOR2_X1 U1536 ( .A1(n889), .A2(n923), .ZN(n894) );
  INV_X1 U1537 ( .A(n988), .ZN(n919) );
  NAND2_X1 U1538 ( .A1(n894), .A2(n919), .ZN(n896) );
  INV_X1 U1539 ( .A(n890), .ZN(n920) );
  INV_X1 U1540 ( .A(n891), .ZN(n892) );
  OAI21_X1 U1541 ( .B1(n892), .B2(n923), .A(n924), .ZN(n893) );
  AOI21_X1 U1542 ( .B1(n894), .B2(n920), .A(n893), .ZN(n895) );
  OAI21_X1 U1543 ( .B1(n1011), .B2(n896), .A(n895), .ZN(n901) );
  NAND2_X1 U1545 ( .A1(n4293), .A2(n898), .ZN(n900) );
  XNOR2_X1 U1546 ( .A(n901), .B(n900), .ZN(n3581) );
  MUX2_X1 U1547 ( .A(n902), .B(n969), .S(bmask_b_i[3]), .Z(n1197) );
  NAND2_X1 U1548 ( .A1(n1197), .A2(n1196), .ZN(n3105) );
  NOR2_X1 U1549 ( .A1(n3105), .A2(n1223), .ZN(n1032) );
  NAND2_X1 U1550 ( .A1(n1461), .A2(n1472), .ZN(n1037) );
  INV_X1 U1551 ( .A(n903), .ZN(n990) );
  NAND2_X1 U1552 ( .A1(n919), .A2(n990), .ZN(n906) );
  INV_X1 U1553 ( .A(n989), .ZN(n904) );
  AOI21_X1 U1554 ( .B1(n920), .B2(n990), .A(n904), .ZN(n905) );
  OAI21_X1 U1555 ( .B1(n1011), .B2(n906), .A(n905), .ZN(n911) );
  INV_X1 U1556 ( .A(n907), .ZN(n909) );
  NAND2_X1 U1557 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1558 ( .A(n911), .B(n910), .ZN(n3627) );
  NAND2_X1 U1559 ( .A1(n912), .A2(n1109), .ZN(n917) );
  NAND2_X1 U1560 ( .A1(bmask_b_i[2]), .A2(bmask_b_i[3]), .ZN(n913) );
  OAI22_X1 U1561 ( .A1(n914), .A2(n1106), .B1(n4119), .B2(n913), .ZN(n915) );
  INV_X1 U1562 ( .A(n915), .ZN(n916) );
  NAND2_X1 U1563 ( .A1(n917), .A2(n916), .ZN(n1141) );
  NOR2_X1 U1564 ( .A1(n1141), .A2(bmask_b_i[4]), .ZN(n3251) );
  AND2_X1 U1565 ( .A1(n3251), .A2(n918), .ZN(n1029) );
  OR2_X1 U1566 ( .A1(n3627), .A2(n1029), .ZN(n1541) );
  NAND2_X1 U1567 ( .A1(n919), .A2(n888), .ZN(n922) );
  AOI21_X1 U1568 ( .B1(n920), .B2(n888), .A(n891), .ZN(n921) );
  OAI21_X1 U1569 ( .B1(n1011), .B2(n922), .A(n921), .ZN(n927) );
  INV_X1 U1570 ( .A(n923), .ZN(n925) );
  NAND2_X1 U1571 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1572 ( .A(n927), .B(n926), .ZN(n3242) );
  OR2_X1 U1573 ( .A1(n928), .A2(bmask_b_i[3]), .ZN(n1175) );
  AOI21_X1 U1574 ( .B1(n1174), .B2(bmask_b_i[3]), .A(bmask_b_i[4]), .ZN(n929)
         );
  NAND2_X1 U1575 ( .A1(n1175), .A2(n929), .ZN(n3591) );
  NOR2_X1 U1576 ( .A1(n3591), .A2(n1223), .ZN(n1030) );
  NAND2_X1 U1577 ( .A1(n1541), .A2(n1536), .ZN(n1467) );
  NAND2_X1 U1578 ( .A1(n1038), .A2(n1492), .ZN(n1041) );
  INV_X1 U1579 ( .A(n930), .ZN(n964) );
  INV_X1 U1580 ( .A(n931), .ZN(n938) );
  INV_X1 U1581 ( .A(n937), .ZN(n932) );
  AOI21_X1 U1582 ( .B1(n964), .B2(n938), .A(n932), .ZN(n936) );
  NAND2_X1 U1583 ( .A1(n166), .A2(n934), .ZN(n935) );
  XOR2_X1 U1584 ( .A(n936), .B(n935), .Z(n3811) );
  OR2_X1 U1585 ( .A1(n1174), .A2(n1218), .ZN(n3754) );
  NOR2_X1 U1586 ( .A1(n3754), .A2(n546), .ZN(n946) );
  NOR2_X1 U1587 ( .A1(n3811), .A2(n946), .ZN(n1410) );
  NAND2_X1 U1588 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1589 ( .A(n964), .B(n939), .ZN(n3466) );
  NOR2_X1 U1590 ( .A1(n940), .A2(n1218), .ZN(n3827) );
  INV_X1 U1591 ( .A(n3827), .ZN(n941) );
  NOR2_X1 U1592 ( .A1(n941), .A2(n546), .ZN(n945) );
  NOR2_X1 U1593 ( .A1(n3466), .A2(n945), .ZN(n1417) );
  NOR2_X1 U1594 ( .A1(n1410), .A2(n1417), .ZN(n948) );
  OAI21_X1 U1595 ( .B1(n944), .B2(n943), .A(n942), .ZN(n1409) );
  NAND2_X1 U1596 ( .A1(n3466), .A2(n945), .ZN(n1418) );
  NAND2_X1 U1597 ( .A1(n3811), .A2(n946), .ZN(n1411) );
  OAI21_X1 U1598 ( .B1(n1410), .B2(n1418), .A(n1411), .ZN(n947) );
  AOI21_X1 U1599 ( .B1(n948), .B2(n1409), .A(n947), .ZN(n1427) );
  INV_X1 U1600 ( .A(n949), .ZN(n951) );
  NOR2_X1 U1601 ( .A1(n951), .A2(n4297), .ZN(n955) );
  INV_X1 U1602 ( .A(n952), .ZN(n953) );
  OAI21_X1 U1603 ( .B1(n953), .B2(n4297), .A(n965), .ZN(n954) );
  AOI21_X1 U1604 ( .B1(n955), .B2(n964), .A(n954), .ZN(n960) );
  INV_X1 U1605 ( .A(n956), .ZN(n958) );
  NAND2_X1 U1606 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1607 ( .A(n960), .B(n959), .Z(n3643) );
  AND2_X1 U1608 ( .A1(n961), .A2(n1171), .ZN(n4004) );
  INV_X1 U1609 ( .A(n4004), .ZN(n962) );
  NOR2_X1 U1610 ( .A1(n962), .A2(n1223), .ZN(n971) );
  OR2_X1 U1611 ( .A1(n3643), .A2(n971), .ZN(n1430) );
  AOI21_X1 U1612 ( .B1(n964), .B2(n165), .A(n952), .ZN(n968) );
  INV_X1 U1613 ( .A(n950), .ZN(n966) );
  NAND2_X1 U1614 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1615 ( .A(n968), .B(n967), .Z(n3719) );
  AND2_X1 U1616 ( .A1(n969), .A2(n1171), .ZN(n3664) );
  INV_X1 U1617 ( .A(n3664), .ZN(n3677) );
  NOR2_X1 U1618 ( .A1(n3677), .A2(n546), .ZN(n970) );
  OR2_X1 U1619 ( .A1(n3719), .A2(n970), .ZN(n1437) );
  NAND2_X1 U1620 ( .A1(n1430), .A2(n1437), .ZN(n974) );
  NAND2_X1 U1621 ( .A1(n3719), .A2(n970), .ZN(n1436) );
  INV_X1 U1622 ( .A(n1436), .ZN(n1428) );
  NAND2_X1 U1623 ( .A1(n3643), .A2(n971), .ZN(n1429) );
  INV_X1 U1624 ( .A(n1429), .ZN(n972) );
  AOI21_X1 U1625 ( .B1(n1430), .B2(n1428), .A(n972), .ZN(n973) );
  OAI21_X1 U1626 ( .B1(n1427), .B2(n974), .A(n973), .ZN(n1443) );
  INV_X1 U1627 ( .A(n975), .ZN(n1000) );
  NAND2_X1 U1628 ( .A1(n995), .A2(n1000), .ZN(n978) );
  INV_X1 U1629 ( .A(n999), .ZN(n976) );
  AOI21_X1 U1630 ( .B1(n996), .B2(n1000), .A(n976), .ZN(n977) );
  OAI21_X1 U1631 ( .B1(n1011), .B2(n978), .A(n977), .ZN(n983) );
  INV_X1 U1632 ( .A(n979), .ZN(n981) );
  NAND2_X1 U1633 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1634 ( .A(n983), .B(n982), .ZN(n3512) );
  NAND2_X1 U1635 ( .A1(n984), .A2(n1196), .ZN(n993) );
  NOR2_X1 U1636 ( .A1(n1078), .A2(n993), .ZN(n985) );
  AOI21_X1 U1637 ( .B1(n986), .B2(n1171), .A(n985), .ZN(n3347) );
  NOR2_X1 U1638 ( .A1(n3347), .A2(n1223), .ZN(n1019) );
  OAI21_X1 U1639 ( .B1(n1011), .B2(n988), .A(n890), .ZN(n992) );
  NAND2_X1 U1640 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1641 ( .A(n992), .B(n991), .ZN(n3337) );
  NOR2_X1 U1642 ( .A1(n1107), .A2(n993), .ZN(n994) );
  AOI21_X1 U1643 ( .B1(n1110), .B2(n1171), .A(n994), .ZN(n3637) );
  NOR2_X1 U1644 ( .A1(n3637), .A2(n1223), .ZN(n1020) );
  OR2_X1 U1645 ( .A1(n3337), .A2(n1020), .ZN(n1519) );
  NAND2_X1 U1646 ( .A1(n1528), .A2(n1519), .ZN(n1023) );
  INV_X1 U1647 ( .A(n995), .ZN(n998) );
  INV_X1 U1648 ( .A(n996), .ZN(n997) );
  OAI21_X1 U1649 ( .B1(n1011), .B2(n998), .A(n997), .ZN(n1002) );
  NAND2_X1 U1650 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1651 ( .A(n1002), .B(n1001), .ZN(n2636) );
  NAND2_X1 U1652 ( .A1(n1003), .A2(n1196), .ZN(n1006) );
  NAND3_X1 U1653 ( .A1(n1004), .A2(bmask_b_i[2]), .A3(n1171), .ZN(n1005) );
  NAND2_X1 U1654 ( .A1(n1006), .A2(n1005), .ZN(n3523) );
  INV_X1 U1655 ( .A(n3523), .ZN(n1007) );
  NOR2_X1 U1656 ( .A1(n1007), .A2(n1223), .ZN(n1016) );
  INV_X1 U1657 ( .A(n1008), .ZN(n1010) );
  OAI22_X1 U1658 ( .A1(n1013), .A2(n1218), .B1(bmask_b_i[4]), .B2(n1012), .ZN(
        n2735) );
  INV_X1 U1659 ( .A(n2735), .ZN(n1014) );
  NOR2_X1 U1660 ( .A1(n1014), .A2(n1223), .ZN(n1015) );
  NOR2_X1 U1661 ( .A1(n3992), .A2(n1015), .ZN(n1444) );
  INV_X1 U1662 ( .A(n1444), .ZN(n1452) );
  NAND2_X1 U1663 ( .A1(n1445), .A2(n1452), .ZN(n1525) );
  NOR2_X1 U1664 ( .A1(n1023), .A2(n1525), .ZN(n1025) );
  NAND2_X1 U1668 ( .A1(n3512), .A2(n1019), .ZN(n1527) );
  INV_X1 U1669 ( .A(n1527), .ZN(n1514) );
  AOI21_X1 U1672 ( .B1(n1514), .B2(n1519), .A(n4273), .ZN(n1022) );
  OAI21_X1 U1673 ( .B1(n1023), .B2(n1524), .A(n1022), .ZN(n1024) );
  NAND2_X1 U1674 ( .A1(n3779), .A2(n1027), .ZN(n1485) );
  OAI21_X1 U1675 ( .B1(n1484), .B2(n1494), .A(n1485), .ZN(n1028) );
  INV_X1 U1676 ( .A(n1028), .ZN(n1040) );
  NAND2_X1 U1677 ( .A1(n3581), .A2(n1032), .ZN(n1471) );
  INV_X1 U1678 ( .A(n1471), .ZN(n1035) );
  AOI21_X1 U1679 ( .B1(n1461), .B2(n1035), .A(n1034), .ZN(n1036) );
  OAI21_X1 U1680 ( .B1(n1037), .B2(n1468), .A(n1036), .ZN(n1480) );
  NAND2_X1 U1681 ( .A1(n1480), .A2(n1038), .ZN(n1039) );
  NAND2_X1 U1683 ( .A1(n2987), .A2(n1042), .ZN(n1378) );
  NAND2_X1 U1684 ( .A1(n1043), .A2(n1044), .ZN(n1370) );
  OAI21_X1 U1685 ( .B1(n1369), .B2(n1378), .A(n1370), .ZN(n1383) );
  NAND2_X1 U1686 ( .A1(n3922), .A2(n1046), .ZN(n1389) );
  OAI21_X1 U1687 ( .B1(n1388), .B2(n1396), .A(n1389), .ZN(n1047) );
  AOI21_X1 U1688 ( .B1(n1383), .B2(n1048), .A(n1047), .ZN(n1325) );
  NAND2_X1 U1689 ( .A1(n3274), .A2(n1049), .ZN(n1336) );
  NAND2_X1 U1690 ( .A1(n3133), .A2(n1051), .ZN(n1331) );
  OAI21_X1 U1691 ( .B1(n1330), .B2(n1336), .A(n1331), .ZN(n1343) );
  NAND2_X1 U1692 ( .A1(n2952), .A2(n1052), .ZN(n1360) );
  NAND2_X1 U1693 ( .A1(n3542), .A2(n1053), .ZN(n1350) );
  OAI21_X1 U1694 ( .B1(n1349), .B2(n1360), .A(n1350), .ZN(n1054) );
  AOI21_X1 U1695 ( .B1(n1055), .B2(n1343), .A(n1054), .ZN(n1056) );
  OAI21_X1 U1696 ( .B1(n1325), .B2(n1057), .A(n1056), .ZN(n1058) );
  NAND2_X1 U1698 ( .A1(n89), .A2(n1061), .ZN(n1063) );
  NOR2_X1 U1699 ( .A1(n1116), .A2(n1063), .ZN(n1065) );
  INV_X1 U1700 ( .A(n1156), .ZN(n1120) );
  INV_X1 U1701 ( .A(n1091), .ZN(n1060) );
  AOI21_X1 U1702 ( .B1(n1120), .B2(n1061), .A(n1060), .ZN(n1062) );
  OAI21_X1 U1703 ( .B1(n1123), .B2(n1063), .A(n1062), .ZN(n1064) );
  AOI21_X1 U1704 ( .B1(n4291), .B2(n1065), .A(n1064), .ZN(n1071) );
  INV_X1 U1705 ( .A(operand_b_i[9]), .ZN(n2567) );
  MUX2_X1 U1706 ( .A(n169), .B(n1205), .S(operand_a_i[25]), .Z(n1066) );
  OAI21_X1 U1707 ( .B1(n76), .B2(n2567), .A(n1066), .ZN(n1069) );
  MUX2_X1 U1708 ( .A(n1247), .B(n1128), .S(operand_b_i[25]), .Z(n1067) );
  OAI21_X1 U1709 ( .B1(operand_a_i[9]), .B2(n540), .A(n1067), .ZN(n1068) );
  INV_X1 U1710 ( .A(n1092), .ZN(n1070) );
  NAND2_X1 U1711 ( .A1(n1069), .A2(n1068), .ZN(n1090) );
  NAND3_X1 U1712 ( .A1(n1073), .A2(bmask_a_i[4]), .A3(n1072), .ZN(n1074) );
  NAND2_X1 U1713 ( .A1(n1074), .A2(n1171), .ZN(n1188) );
  OAI21_X1 U1714 ( .B1(n1075), .B2(n1214), .A(n1188), .ZN(n1077) );
  NAND2_X1 U1715 ( .A1(n1077), .A2(n1076), .ZN(n1088) );
  AOI22_X1 U1716 ( .A1(n1080), .A2(n1079), .B1(n1078), .B2(n1173), .ZN(n1087)
         );
  NAND2_X1 U1717 ( .A1(n1081), .A2(n1196), .ZN(n1082) );
  OAI211_X1 U1718 ( .C1(bmask_b_i[3]), .C2(n1083), .A(n1082), .B(bmask_b_i[2]), 
        .ZN(n1086) );
  OR2_X1 U1719 ( .A1(n1084), .A2(n1218), .ZN(n1085) );
  NAND4_X1 U1720 ( .A1(n1088), .A2(n1087), .A3(n1086), .A4(n1085), .ZN(n3206)
         );
  NOR2_X1 U1721 ( .A1(n3206), .A2(n1223), .ZN(n1224) );
  NOR2_X1 U1722 ( .A1(n4051), .A2(n1224), .ZN(n1311) );
  NAND2_X1 U1723 ( .A1(n89), .A2(n1145), .ZN(n1094) );
  NOR2_X1 U1724 ( .A1(n1116), .A2(n1094), .ZN(n1096) );
  OAI21_X1 U1725 ( .B1(n1092), .B2(n1091), .A(n1090), .ZN(n1152) );
  AOI21_X1 U1726 ( .B1(n1120), .B2(n1145), .A(n1152), .ZN(n1093) );
  OAI21_X1 U1727 ( .B1(n1123), .B2(n1094), .A(n1093), .ZN(n1095) );
  AOI21_X1 U1728 ( .B1(n4291), .B2(n1096), .A(n1095), .ZN(n1103) );
  INV_X1 U1729 ( .A(operand_b_i[10]), .ZN(n2571) );
  MUX2_X1 U1731 ( .A(n2949), .B(n74), .S(operand_a_i[26]), .Z(n1098) );
  OAI21_X1 U1732 ( .B1(n76), .B2(n2571), .A(n1098), .ZN(n1101) );
  MUX2_X1 U1733 ( .A(n1207), .B(n587), .S(n170), .Z(n1099) );
  OAI21_X1 U1734 ( .B1(n168), .B2(n540), .A(n1099), .ZN(n1100) );
  NOR2_X1 U1735 ( .A1(n1101), .A2(n1100), .ZN(n1144) );
  INV_X1 U1736 ( .A(n1144), .ZN(n1102) );
  NAND2_X1 U1737 ( .A1(n1101), .A2(n1100), .ZN(n1149) );
  NOR2_X1 U1738 ( .A1(n1104), .A2(n2369), .ZN(n1219) );
  OAI22_X1 U1739 ( .A1(n1219), .A2(n1217), .B1(n1105), .B2(n1218), .ZN(n1112)
         );
  OAI21_X1 U1740 ( .B1(n1107), .B2(n1106), .A(bmask_b_i[4]), .ZN(n1108) );
  AOI21_X1 U1741 ( .B1(n1110), .B2(n1109), .A(n1108), .ZN(n1111) );
  NOR2_X1 U1742 ( .A1(n1112), .A2(n1111), .ZN(n1113) );
  OAI21_X1 U1743 ( .B1(n1114), .B2(n1214), .A(n1113), .ZN(n2875) );
  NOR2_X1 U1744 ( .A1(n2875), .A2(n1223), .ZN(n1225) );
  NOR2_X1 U1745 ( .A1(n3197), .A2(n1225), .ZN(n1306) );
  INV_X1 U1746 ( .A(n1145), .ZN(n1115) );
  NOR2_X1 U1747 ( .A1(n1115), .A2(n1144), .ZN(n1119) );
  NAND2_X1 U1748 ( .A1(n1119), .A2(n89), .ZN(n1122) );
  NOR2_X1 U1749 ( .A1(n1116), .A2(n1122), .ZN(n1125) );
  INV_X1 U1750 ( .A(n1152), .ZN(n1117) );
  OAI21_X1 U1751 ( .B1(n1117), .B2(n1144), .A(n1149), .ZN(n1118) );
  AOI21_X1 U1752 ( .B1(n1120), .B2(n1119), .A(n1118), .ZN(n1121) );
  OAI21_X1 U1753 ( .B1(n1123), .B2(n1122), .A(n1121), .ZN(n1124) );
  AOI21_X1 U1754 ( .B1(n4291), .B2(n1125), .A(n1124), .ZN(n1134) );
  MUX2_X1 U1755 ( .A(n704), .B(n169), .S(n2521), .Z(n1127) );
  OAI21_X1 U1756 ( .B1(n75), .B2(n2562), .A(n1127), .ZN(n1131) );
  MUX2_X1 U1757 ( .A(n817), .B(n1128), .S(n64), .Z(n1129) );
  OAI21_X1 U1758 ( .B1(operand_a_i[11]), .B2(n540), .A(n1129), .ZN(n1130) );
  NOR2_X1 U1759 ( .A1(n1131), .A2(n1130), .ZN(n1150) );
  INV_X1 U1760 ( .A(n1150), .ZN(n1132) );
  NAND2_X1 U1761 ( .A1(n1131), .A2(n1130), .ZN(n1148) );
  INV_X1 U1764 ( .A(n1135), .ZN(n1137) );
  AOI22_X1 U1765 ( .A1(n1137), .A2(n4120), .B1(n1136), .B2(n1171), .ZN(n1138)
         );
  OAI21_X1 U1766 ( .B1(n1214), .B2(n1139), .A(n1138), .ZN(n1140) );
  AOI21_X1 U1767 ( .B1(n1141), .B2(bmask_b_i[4]), .A(n1140), .ZN(n3855) );
  INV_X1 U1768 ( .A(n3855), .ZN(n1142) );
  NOR2_X1 U1769 ( .A1(n1142), .A2(n1223), .ZN(n1226) );
  NOR2_X1 U1770 ( .A1(n2864), .A2(n1226), .ZN(n1289) );
  NOR2_X1 U1771 ( .A1(n1144), .A2(n1150), .ZN(n1153) );
  NAND2_X1 U1772 ( .A1(n1145), .A2(n1153), .ZN(n1155) );
  NOR2_X1 U1773 ( .A1(n1146), .A2(n1155), .ZN(n1159) );
  NAND2_X1 U1774 ( .A1(n1159), .A2(n1147), .ZN(n1161) );
  OAI21_X1 U1775 ( .B1(n1150), .B2(n1149), .A(n1148), .ZN(n1151) );
  AOI21_X1 U1776 ( .B1(n1153), .B2(n1152), .A(n1151), .ZN(n1154) );
  OAI21_X1 U1777 ( .B1(n1156), .B2(n1155), .A(n1154), .ZN(n1157) );
  AOI21_X1 U1778 ( .B1(n1159), .B2(n4308), .A(n1157), .ZN(n1160) );
  OAI21_X1 U1779 ( .B1(n1162), .B2(n1161), .A(n1160), .ZN(n1244) );
  INV_X1 U1780 ( .A(operand_b_i[12]), .ZN(n3240) );
  MUX2_X1 U1781 ( .A(n1205), .B(n2949), .S(n2522), .Z(n1163) );
  OAI21_X1 U1782 ( .B1(n76), .B2(n3240), .A(n1163), .ZN(n1166) );
  MUX2_X1 U1783 ( .A(n1247), .B(n1128), .S(operand_b_i[28]), .Z(n1164) );
  OAI21_X1 U1784 ( .B1(operand_a_i[12]), .B2(n540), .A(n1164), .ZN(n1165) );
  OR2_X1 U1785 ( .A1(n1166), .A2(n1165), .ZN(n1198) );
  NAND2_X1 U1786 ( .A1(n1166), .A2(n1165), .ZN(n1178) );
  NAND2_X1 U1787 ( .A1(n1198), .A2(n1178), .ZN(n1167) );
  XNOR2_X1 U1788 ( .A(n1244), .B(n1167), .ZN(n3869) );
  AND2_X1 U1789 ( .A1(n1168), .A2(n1217), .ZN(n1170) );
  OAI21_X1 U1790 ( .B1(n1170), .B2(n1169), .A(bmask_a_i[4]), .ZN(n1172) );
  AOI22_X1 U1791 ( .A1(n1174), .A2(n1173), .B1(n1172), .B2(n1171), .ZN(n1176)
         );
  OAI211_X1 U1792 ( .C1(n1214), .C2(n1177), .A(n1176), .B(n1175), .ZN(n2773)
         );
  NOR2_X1 U1793 ( .A1(n2773), .A2(n1223), .ZN(n1227) );
  NOR2_X1 U1794 ( .A1(n3869), .A2(n1227), .ZN(n1294) );
  NOR2_X1 U1795 ( .A1(n1294), .A2(n1289), .ZN(n1229) );
  NAND2_X1 U1796 ( .A1(n1299), .A2(n1229), .ZN(n1283) );
  INV_X1 U1797 ( .A(n1178), .ZN(n1201) );
  AOI21_X1 U1798 ( .B1(n4295), .B2(n1198), .A(n1201), .ZN(n1187) );
  INV_X1 U1799 ( .A(operand_b_i[13]), .ZN(n3578) );
  MUX2_X1 U1800 ( .A(n74), .B(n169), .S(n53), .Z(n1179) );
  OAI21_X1 U1801 ( .B1(n75), .B2(n111), .A(n1179), .ZN(n1185) );
  MUX2_X1 U1802 ( .A(n1181), .B(n1180), .S(operand_b_i[29]), .Z(n1183) );
  NOR2_X1 U1803 ( .A1(n540), .A2(operand_a_i[13]), .ZN(n1182) );
  OR2_X1 U1804 ( .A1(n1183), .A2(n1182), .ZN(n1184) );
  OR2_X1 U1805 ( .A1(n1185), .A2(n1184), .ZN(n1202) );
  NAND2_X1 U1806 ( .A1(n1185), .A2(n1184), .ZN(n1199) );
  NAND2_X1 U1807 ( .A1(n1202), .A2(n1199), .ZN(n1186) );
  XOR2_X1 U1808 ( .A(n1187), .B(n1186), .Z(n2834) );
  NAND2_X1 U1809 ( .A1(n1188), .A2(n1217), .ZN(n1192) );
  NAND2_X1 U1810 ( .A1(bmask_a_i[4]), .A2(bmask_a_i[3]), .ZN(n1189) );
  OR2_X1 U1811 ( .A1(n1190), .A2(n1189), .ZN(n1191) );
  AOI22_X1 U1812 ( .A1(n1194), .A2(n1193), .B1(n1192), .B2(n1191), .ZN(n1195)
         );
  OAI21_X1 U1813 ( .B1(n1197), .B2(n1196), .A(n1195), .ZN(n3313) );
  NOR2_X1 U1814 ( .A1(n3313), .A2(n1223), .ZN(n1230) );
  NAND2_X1 U1815 ( .A1(n1198), .A2(n1202), .ZN(n1238) );
  INV_X1 U1816 ( .A(n1238), .ZN(n1204) );
  INV_X1 U1817 ( .A(n1199), .ZN(n1200) );
  AOI21_X1 U1818 ( .B1(n1202), .B2(n1201), .A(n1200), .ZN(n1241) );
  INV_X1 U1819 ( .A(n1241), .ZN(n1203) );
  AOI21_X1 U1820 ( .B1(n1244), .B2(n1204), .A(n1203), .ZN(n1213) );
  INV_X1 U1821 ( .A(operand_b_i[14]), .ZN(n3092) );
  MUX2_X1 U1822 ( .A(n1205), .B(n169), .S(n4112), .Z(n1206) );
  OAI21_X1 U1823 ( .B1(n75), .B2(n3092), .A(n1206), .ZN(n1210) );
  MUX2_X1 U1824 ( .A(n817), .B(n1128), .S(operand_b_i[30]), .Z(n1208) );
  OAI21_X1 U1825 ( .B1(n4300), .B2(n540), .A(n1208), .ZN(n1209) );
  NOR2_X1 U1826 ( .A1(n1210), .A2(n1209), .ZN(n1240) );
  INV_X1 U1827 ( .A(n1240), .ZN(n1211) );
  NAND2_X1 U1828 ( .A1(n1210), .A2(n1209), .ZN(n1239) );
  NAND2_X1 U1829 ( .A1(n1211), .A2(n1239), .ZN(n1212) );
  XOR2_X1 U1830 ( .A(n1213), .B(n1212), .Z(n3290) );
  NOR2_X1 U1831 ( .A1(n1215), .A2(n1214), .ZN(n1221) );
  OAI22_X1 U1832 ( .A1(n1219), .A2(n1218), .B1(n1217), .B2(n1216), .ZN(n1220)
         );
  OR3_X1 U1833 ( .A1(n1222), .A2(n1221), .A3(n1220), .ZN(n3941) );
  NOR2_X1 U1834 ( .A1(n3941), .A2(n1223), .ZN(n1231) );
  OR2_X1 U1835 ( .A1(n3290), .A2(n1231), .ZN(n1278) );
  NAND2_X1 U1836 ( .A1(n1285), .A2(n1278), .ZN(n1234) );
  OR2_X1 U1837 ( .A1(n1283), .A2(n1234), .ZN(n1237) );
  NAND2_X1 U1838 ( .A1(n4051), .A2(n1224), .ZN(n1312) );
  NAND2_X1 U1839 ( .A1(n3197), .A2(n1225), .ZN(n1307) );
  NAND2_X1 U1840 ( .A1(n2864), .A2(n1226), .ZN(n1302) );
  NAND2_X1 U1841 ( .A1(n3869), .A2(n1227), .ZN(n1295) );
  OAI21_X1 U1842 ( .B1(n1294), .B2(n1302), .A(n1295), .ZN(n1228) );
  AOI21_X1 U1843 ( .B1(n1229), .B2(n1290), .A(n1228), .ZN(n1272) );
  NAND2_X1 U1844 ( .A1(n2834), .A2(n1230), .ZN(n1284) );
  INV_X1 U1845 ( .A(n1284), .ZN(n1273) );
  NAND2_X1 U1846 ( .A1(n3290), .A2(n1231), .ZN(n1277) );
  INV_X1 U1847 ( .A(n1277), .ZN(n1232) );
  AOI21_X1 U1848 ( .B1(n1278), .B2(n1273), .A(n1232), .ZN(n1233) );
  OAI21_X1 U1849 ( .B1(n1272), .B2(n1234), .A(n1233), .ZN(n1235) );
  INV_X1 U1850 ( .A(n1235), .ZN(n1236) );
  OAI21_X1 U1851 ( .B1(n1270), .B2(n1237), .A(n1236), .ZN(n1256) );
  NOR2_X1 U1852 ( .A1(n1238), .A2(n1240), .ZN(n1243) );
  OAI21_X1 U1853 ( .B1(n1241), .B2(n1240), .A(n1239), .ZN(n1242) );
  AOI21_X1 U1854 ( .B1(n4295), .B2(n1243), .A(n1242), .ZN(n2408) );
  INV_X1 U1855 ( .A(operand_b_i[15]), .ZN(n3055) );
  MUX2_X1 U1856 ( .A(n74), .B(n2949), .S(n4115), .Z(n1245) );
  OAI21_X1 U1857 ( .B1(n3055), .B2(n76), .A(n1245), .ZN(n1246) );
  INV_X1 U1858 ( .A(n1246), .ZN(n1252) );
  MUX2_X1 U1859 ( .A(n1207), .B(n1128), .S(operand_b_i[31]), .Z(n1248) );
  OAI21_X1 U1860 ( .B1(operand_a_i[15]), .B2(n540), .A(n1248), .ZN(n1250) );
  INV_X1 U1861 ( .A(n1250), .ZN(n1251) );
  NOR2_X1 U1862 ( .A1(n1252), .A2(n1251), .ZN(n2388) );
  INV_X1 U1863 ( .A(n2388), .ZN(n1253) );
  NAND2_X1 U1864 ( .A1(n1252), .A2(n1251), .ZN(n2387) );
  NAND2_X1 U1865 ( .A1(n1253), .A2(n2387), .ZN(n1254) );
  XOR2_X1 U1866 ( .A(n2408), .B(n1254), .Z(n3959) );
  INV_X1 U1867 ( .A(n3959), .ZN(n1255) );
  XNOR2_X1 U1868 ( .A(n1256), .B(n1255), .ZN(n1258) );
  NAND2_X1 U1870 ( .A1(n1267), .A2(n532), .ZN(n2728) );
  INV_X1 U1871 ( .A(n2733), .ZN(n2351) );
  AOI21_X1 U1872 ( .B1(n532), .B2(n52), .A(n4337), .ZN(n1259) );
  OAI21_X1 U1873 ( .B1(n2728), .B2(n2351), .A(n1259), .ZN(n2012) );
  INV_X1 U1874 ( .A(n1261), .ZN(n1619) );
  OR2_X1 U1876 ( .A1(n4176), .A2(n1262), .ZN(n1264) );
  AND2_X1 U1877 ( .A1(n1264), .A2(n1263), .ZN(n1266) );
  OAI22_X1 U1878 ( .A1(n1545), .A2(n4127), .B1(n1544), .B2(n4115), .ZN(n1265)
         );
  AOI21_X1 U1879 ( .B1(n1266), .B2(n82), .A(n1265), .ZN(n1729) );
  OR2_X1 U1880 ( .A1(n1267), .A2(n4130), .ZN(n2106) );
  OR2_X1 U1881 ( .A1(n1729), .A2(n2106), .ZN(n1268) );
  NOR2_X1 U1882 ( .A1(n1730), .A2(n1268), .ZN(n1269) );
  INV_X1 U1883 ( .A(n1283), .ZN(n1271) );
  NAND2_X1 U1884 ( .A1(n1271), .A2(n1285), .ZN(n1276) );
  INV_X1 U1885 ( .A(n1272), .ZN(n1274) );
  AOI21_X1 U1886 ( .B1(n1274), .B2(n1285), .A(n1273), .ZN(n1275) );
  OAI21_X1 U1887 ( .B1(n1315), .B2(n1276), .A(n1275), .ZN(n1280) );
  NAND2_X1 U1888 ( .A1(n1278), .A2(n1277), .ZN(n1279) );
  XNOR2_X1 U1889 ( .A(n1280), .B(n1279), .ZN(n1282) );
  AOI22_X1 U1890 ( .A1(n1532), .A2(n4112), .B1(n91), .B2(n2546), .ZN(n1281) );
  OAI21_X1 U1891 ( .B1(n1282), .B2(n532), .A(n1281), .ZN(n1607) );
  NAND2_X1 U1892 ( .A1(n4272), .A2(n1647), .ZN(n1288) );
  NOR2_X1 U1893 ( .A1(n1788), .A2(n1619), .ZN(n1562) );
  OAI21_X1 U1894 ( .B1(n1315), .B2(n1283), .A(n4296), .ZN(n1286) );
  OAI22_X1 U1895 ( .A1(n1545), .A2(n54), .B1(n2376), .B2(operand_a_i[2]), .ZN(
        n1287) );
  INV_X1 U1896 ( .A(n1944), .ZN(n2004) );
  AND2_X1 U1897 ( .A1(n2290), .A2(n4294), .ZN(n1749) );
  INV_X1 U1898 ( .A(n1289), .ZN(n1303) );
  NAND2_X1 U1899 ( .A1(n1299), .A2(n1303), .ZN(n1293) );
  INV_X1 U1900 ( .A(n1302), .ZN(n1291) );
  AOI21_X1 U1901 ( .B1(n1290), .B2(n1303), .A(n1291), .ZN(n1292) );
  OAI21_X1 U1902 ( .B1(n1315), .B2(n1293), .A(n1292), .ZN(n1297) );
  INV_X1 U1903 ( .A(n1294), .ZN(n1296) );
  OAI22_X1 U1904 ( .A1(n1545), .A2(operand_a_i[28]), .B1(n1544), .B2(n48), 
        .ZN(n1298) );
  INV_X1 U1905 ( .A(n1299), .ZN(n1301) );
  INV_X1 U1906 ( .A(n1290), .ZN(n1300) );
  OAI21_X1 U1907 ( .B1(n1315), .B2(n1301), .A(n1300), .ZN(n1304) );
  OAI22_X1 U1908 ( .A1(n1545), .A2(operand_a_i[27]), .B1(n1544), .B2(
        operand_a_i[4]), .ZN(n1305) );
  OAI21_X1 U1909 ( .B1(n1315), .B2(n1311), .A(n1312), .ZN(n1309) );
  INV_X1 U1910 ( .A(n1306), .ZN(n1308) );
  OAI22_X1 U1911 ( .A1(n1545), .A2(operand_a_i[26]), .B1(n1544), .B2(
        operand_a_i[5]), .ZN(n1310) );
  INV_X1 U1913 ( .A(n1311), .ZN(n1313) );
  NAND2_X1 U1914 ( .A1(n1313), .A2(n1312), .ZN(n1314) );
  XOR2_X1 U1915 ( .A(n1315), .B(n1314), .Z(n1316) );
  AOI22_X1 U1916 ( .A1(n1532), .A2(operand_a_i[25]), .B1(operand_a_i[6]), .B2(
        n91), .ZN(n1317) );
  AOI22_X1 U1918 ( .A1(n1749), .A2(n1713), .B1(n2174), .B2(n1824), .ZN(n1318)
         );
  NAND2_X1 U1919 ( .A1(n1319), .A2(n1318), .ZN(n2192) );
  INV_X1 U1922 ( .A(n1324), .ZN(n1337) );
  NAND2_X1 U1923 ( .A1(n88), .A2(n1337), .ZN(n1329) );
  INV_X1 U1925 ( .A(n1325), .ZN(n1357) );
  INV_X1 U1926 ( .A(n1336), .ZN(n1327) );
  AOI21_X1 U1927 ( .B1(n1357), .B2(n1337), .A(n1327), .ZN(n1328) );
  OAI21_X1 U1928 ( .B1(n1395), .B2(n1329), .A(n1328), .ZN(n1333) );
  OAI22_X1 U1930 ( .A1(n1545), .A2(operand_a_i[22]), .B1(n2376), .B2(
        operand_a_i[9]), .ZN(n1334) );
  INV_X1 U1931 ( .A(n1895), .ZN(n2076) );
  NAND2_X1 U1932 ( .A1(n4272), .A2(n2076), .ZN(n1368) );
  AOI22_X1 U1933 ( .A1(n1532), .A2(operand_a_i[21]), .B1(n168), .B2(n91), .ZN(
        n1339) );
  NAND2_X1 U1934 ( .A1(n1340), .A2(n1339), .ZN(n2117) );
  INV_X1 U1935 ( .A(n2117), .ZN(n2077) );
  NAND2_X1 U1936 ( .A1(n1821), .A2(n2077), .ZN(n1367) );
  INV_X1 U1937 ( .A(n1341), .ZN(n1342) );
  NOR2_X1 U1938 ( .A1(n1342), .A2(n1359), .ZN(n1346) );
  NAND2_X1 U1939 ( .A1(n1346), .A2(n88), .ZN(n1348) );
  INV_X1 U1940 ( .A(n1356), .ZN(n1344) );
  OAI21_X1 U1941 ( .B1(n1344), .B2(n1359), .A(n1360), .ZN(n1345) );
  AOI21_X1 U1942 ( .B1(n1346), .B2(n1357), .A(n1345), .ZN(n1347) );
  OAI21_X1 U1943 ( .B1(n1395), .B2(n1348), .A(n1347), .ZN(n1353) );
  INV_X1 U1944 ( .A(n1349), .ZN(n1351) );
  NAND2_X1 U1945 ( .A1(n1351), .A2(n1350), .ZN(n1352) );
  XNOR2_X1 U1946 ( .A(n1353), .B(n1352), .ZN(n1354) );
  AOI22_X1 U1947 ( .A1(n1532), .A2(operand_a_i[24]), .B1(operand_a_i[7]), .B2(
        n91), .ZN(n1355) );
  OR2_X1 U1948 ( .A1(n1764), .A2(n2009), .ZN(n1366) );
  AOI21_X1 U1949 ( .B1(n1357), .B2(n1341), .A(n1356), .ZN(n1358) );
  INV_X1 U1950 ( .A(n1359), .ZN(n1361) );
  NAND2_X1 U1951 ( .A1(n1361), .A2(n1360), .ZN(n1362) );
  AOI22_X1 U1952 ( .A1(n1532), .A2(operand_a_i[23]), .B1(n149), .B2(n91), .ZN(
        n1363) );
  OR2_X1 U1953 ( .A1(n1751), .A2(n2013), .ZN(n1365) );
  NAND4_X1 U1954 ( .A1(n1368), .A2(n1367), .A3(n1366), .A4(n1365), .ZN(n2205)
         );
  INV_X1 U1956 ( .A(n1369), .ZN(n1371) );
  NAND2_X1 U1957 ( .A1(n1371), .A2(n1370), .ZN(n1372) );
  XNOR2_X1 U1958 ( .A(n1373), .B(n1372), .ZN(n1374) );
  NAND2_X1 U1959 ( .A1(n1374), .A2(n82), .ZN(n1376) );
  AOI22_X1 U1960 ( .A1(n1532), .A2(n72), .B1(operand_a_i[13]), .B2(n91), .ZN(
        n1375) );
  NAND2_X1 U1961 ( .A1(n1376), .A2(n1375), .ZN(n2027) );
  INV_X1 U1962 ( .A(n2027), .ZN(n2157) );
  NAND2_X1 U1963 ( .A1(n1321), .A2(n2157), .ZN(n1405) );
  NAND2_X1 U1965 ( .A1(n4326), .A2(n1378), .ZN(n1380) );
  OAI22_X1 U1966 ( .A1(n1545), .A2(operand_a_i[17]), .B1(n2376), .B2(n4300), 
        .ZN(n1381) );
  AOI21_X1 U1967 ( .B1(n185), .B2(n82), .A(n1381), .ZN(n1716) );
  INV_X1 U1968 ( .A(n1716), .ZN(n2154) );
  NAND2_X1 U1969 ( .A1(n1821), .A2(n2154), .ZN(n1404) );
  INV_X1 U1970 ( .A(n1382), .ZN(n1397) );
  NAND2_X1 U1971 ( .A1(n1392), .A2(n1397), .ZN(n1387) );
  INV_X1 U1972 ( .A(n1396), .ZN(n1385) );
  AOI21_X1 U1973 ( .B1(n1384), .B2(n1397), .A(n1385), .ZN(n1386) );
  NAND2_X1 U1974 ( .A1(n155), .A2(n1389), .ZN(n1390) );
  OAI22_X1 U1975 ( .A1(n1545), .A2(operand_a_i[20]), .B1(n2376), .B2(
        operand_a_i[11]), .ZN(n1391) );
  OR2_X1 U1976 ( .A1(n1764), .A2(n2116), .ZN(n1403) );
  INV_X1 U1977 ( .A(n1392), .ZN(n1394) );
  INV_X1 U1978 ( .A(n1384), .ZN(n1393) );
  OAI21_X1 U1979 ( .B1(n1395), .B2(n1394), .A(n1393), .ZN(n1399) );
  NAND2_X1 U1980 ( .A1(n1397), .A2(n1396), .ZN(n1398) );
  XNOR2_X1 U1981 ( .A(n1399), .B(n1398), .ZN(n1401) );
  OAI22_X1 U1982 ( .A1(n1545), .A2(n4105), .B1(n2376), .B2(n2561), .ZN(n1400)
         );
  INV_X1 U1983 ( .A(n2161), .ZN(n2028) );
  MUX2_X1 U1986 ( .A(n2205), .B(n2294), .S(n1635), .Z(n2149) );
  AOI22_X1 U1988 ( .A1(n2192), .A2(n2108), .B1(n4233), .B2(n4331), .ZN(n1407)
         );
  OAI21_X1 U1989 ( .B1(n1810), .B2(n1408), .A(n1407), .ZN(n1426) );
  OR2_X1 U1990 ( .A1(n2217), .A2(n437), .ZN(n1809) );
  INV_X1 U1991 ( .A(n1409), .ZN(n1421) );
  OAI21_X1 U1992 ( .B1(n1421), .B2(n1417), .A(n1418), .ZN(n1414) );
  INV_X1 U1993 ( .A(n1410), .ZN(n1412) );
  NAND2_X1 U1994 ( .A1(n1412), .A2(n1411), .ZN(n1413) );
  XNOR2_X1 U1995 ( .A(n1414), .B(n1413), .ZN(n1416) );
  OAI22_X1 U1996 ( .A1(n1545), .A2(n4108), .B1(n1544), .B2(n2521), .ZN(n1415)
         );
  AOI21_X1 U1997 ( .B1(n1416), .B2(n82), .A(n1415), .ZN(n1676) );
  INV_X1 U1998 ( .A(n1417), .ZN(n1419) );
  NAND2_X1 U1999 ( .A1(n1419), .A2(n1418), .ZN(n1420) );
  XOR2_X1 U2000 ( .A(n1421), .B(n1420), .Z(n1422) );
  NAND2_X1 U2001 ( .A1(n1422), .A2(n82), .ZN(n1424) );
  AOI22_X1 U2002 ( .A1(n1532), .A2(n48), .B1(operand_a_i[28]), .B2(n91), .ZN(
        n1423) );
  NAND2_X1 U2003 ( .A1(n1424), .A2(n1423), .ZN(n1557) );
  INV_X1 U2004 ( .A(n1557), .ZN(n1658) );
  MUX2_X1 U2005 ( .A(n1676), .B(n1658), .S(n1730), .Z(n1811) );
  NOR2_X1 U2006 ( .A1(n1809), .A2(n1811), .ZN(n1425) );
  NOR2_X1 U2007 ( .A1(n1426), .A2(n1425), .ZN(n1555) );
  INV_X1 U2008 ( .A(n1427), .ZN(n1439) );
  AOI21_X1 U2009 ( .B1(n1439), .B2(n1437), .A(n1428), .ZN(n1432) );
  NAND2_X1 U2010 ( .A1(n1430), .A2(n1429), .ZN(n1431) );
  XOR2_X1 U2011 ( .A(n1432), .B(n1431), .Z(n1433) );
  NAND2_X1 U2012 ( .A1(n1433), .A2(n82), .ZN(n1435) );
  AOI22_X1 U2013 ( .A1(n1532), .A2(operand_a_i[6]), .B1(operand_a_i[25]), .B2(
        n91), .ZN(n1434) );
  NAND2_X1 U2014 ( .A1(n1435), .A2(n1434), .ZN(n1680) );
  INV_X1 U2015 ( .A(n1680), .ZN(n1661) );
  NAND2_X1 U2016 ( .A1(n1437), .A2(n1436), .ZN(n1438) );
  XNOR2_X1 U2017 ( .A(n1439), .B(n1438), .ZN(n1441) );
  OAI22_X1 U2018 ( .A1(n1545), .A2(n4079), .B1(n1544), .B2(n3848), .ZN(n1440)
         );
  AOI21_X1 U2019 ( .B1(n1441), .B2(n82), .A(n1440), .ZN(n1656) );
  MUX2_X1 U2020 ( .A(n1661), .B(n1656), .S(n1657), .Z(n1808) );
  NOR2_X1 U2021 ( .A1(n2217), .A2(n1808), .ZN(n1442) );
  NAND2_X1 U2022 ( .A1(n1442), .A2(n1620), .ZN(n1512) );
  INV_X1 U2023 ( .A(n1443), .ZN(n1526) );
  OAI21_X1 U2024 ( .B1(n1526), .B2(n1444), .A(n1451), .ZN(n1447) );
  XNOR2_X1 U2025 ( .A(n1447), .B(n1446), .ZN(n1448) );
  NAND2_X1 U2026 ( .A1(n1448), .A2(n82), .ZN(n1450) );
  AOI22_X1 U2027 ( .A1(n1532), .A2(n149), .B1(operand_a_i[23]), .B2(n91), .ZN(
        n1449) );
  NAND2_X1 U2028 ( .A1(n1450), .A2(n1449), .ZN(n1984) );
  NAND2_X1 U2029 ( .A1(n1452), .A2(n1451), .ZN(n1453) );
  XOR2_X1 U2030 ( .A(n1526), .B(n1453), .Z(n1454) );
  NAND2_X1 U2031 ( .A1(n1454), .A2(n82), .ZN(n1456) );
  AOI22_X1 U2032 ( .A1(n1532), .A2(operand_a_i[7]), .B1(operand_a_i[24]), .B2(
        n91), .ZN(n1455) );
  NAND2_X1 U2033 ( .A1(n1456), .A2(n1455), .ZN(n2171) );
  MUX2_X1 U2034 ( .A(n1984), .B(n2171), .S(n1657), .Z(n1457) );
  NAND3_X1 U2035 ( .A1(n2170), .A2(n4294), .A3(n1457), .ZN(n1507) );
  AOI21_X1 U2037 ( .B1(n1543), .B2(n1460), .A(n1459), .ZN(n1463) );
  XOR2_X1 U2038 ( .A(n1463), .B(n1462), .Z(n1464) );
  NAND2_X1 U2039 ( .A1(n1464), .A2(n82), .ZN(n1466) );
  AOI22_X1 U2040 ( .A1(n1532), .A2(n4300), .B1(operand_a_i[17]), .B2(n91), 
        .ZN(n1465) );
  NAND2_X1 U2041 ( .A1(n1466), .A2(n1465), .ZN(n1914) );
  NAND2_X1 U2042 ( .A1(n1321), .A2(n1914), .ZN(n1478) );
  INV_X1 U2043 ( .A(n1467), .ZN(n1470) );
  INV_X1 U2044 ( .A(n58), .ZN(n1469) );
  AOI21_X1 U2045 ( .B1(n1543), .B2(n1470), .A(n1469), .ZN(n1474) );
  NAND2_X1 U2046 ( .A1(n1472), .A2(n1471), .ZN(n1473) );
  XOR2_X1 U2047 ( .A(n1474), .B(n1473), .Z(n1476) );
  OAI22_X1 U2048 ( .A1(n1545), .A2(n4101), .B1(n1544), .B2(n71), .ZN(n1475) );
  AOI21_X1 U2049 ( .B1(n1476), .B2(n82), .A(n1475), .ZN(n1918) );
  INV_X1 U2050 ( .A(n1918), .ZN(n1757) );
  NAND2_X1 U2051 ( .A1(n1821), .A2(n1757), .ZN(n1477) );
  NAND2_X1 U2052 ( .A1(n1478), .A2(n1477), .ZN(n1504) );
  INV_X1 U2053 ( .A(n1492), .ZN(n1479) );
  NOR2_X1 U2054 ( .A1(n1479), .A2(n1493), .ZN(n1483) );
  INV_X1 U2055 ( .A(n1480), .ZN(n1481) );
  OAI21_X1 U2056 ( .B1(n1481), .B2(n1493), .A(n1494), .ZN(n1482) );
  AOI21_X1 U2057 ( .B1(n1483), .B2(n1543), .A(n1482), .ZN(n1488) );
  INV_X1 U2058 ( .A(n1484), .ZN(n1486) );
  NAND2_X1 U2059 ( .A1(n1486), .A2(n1485), .ZN(n1487) );
  XOR2_X1 U2060 ( .A(n1488), .B(n1487), .Z(n1489) );
  NAND2_X1 U2061 ( .A1(n1489), .A2(n82), .ZN(n1491) );
  AOI22_X1 U2062 ( .A1(n1532), .A2(operand_a_i[16]), .B1(operand_a_i[15]), 
        .B2(n91), .ZN(n1490) );
  AOI21_X1 U2063 ( .B1(n1543), .B2(n1492), .A(n57), .ZN(n1497) );
  INV_X1 U2064 ( .A(n1493), .ZN(n1495) );
  NAND2_X1 U2065 ( .A1(n1495), .A2(n1494), .ZN(n1496) );
  XOR2_X1 U2066 ( .A(n1497), .B(n1496), .Z(n1498) );
  NAND2_X1 U2067 ( .A1(n1498), .A2(n82), .ZN(n1500) );
  AOI22_X1 U2068 ( .A1(n1532), .A2(operand_a_i[15]), .B1(operand_a_i[16]), 
        .B2(n91), .ZN(n1499) );
  NAND2_X1 U2069 ( .A1(n1500), .A2(n1499), .ZN(n1915) );
  INV_X1 U2070 ( .A(n1915), .ZN(n1501) );
  MUX2_X1 U2071 ( .A(n180), .B(n1501), .S(n1730), .Z(n1715) );
  NOR2_X1 U2072 ( .A1(n1715), .A2(n1620), .ZN(n1502) );
  NOR2_X1 U2073 ( .A1(n1504), .A2(n1502), .ZN(n2143) );
  OR2_X1 U2074 ( .A1(n1657), .A2(n426), .ZN(n1508) );
  NAND2_X1 U2075 ( .A1(n1508), .A2(n1915), .ZN(n1827) );
  NOR2_X1 U2076 ( .A1(n1827), .A2(n1620), .ZN(n1503) );
  NOR2_X1 U2077 ( .A1(n1504), .A2(n1503), .ZN(n1955) );
  NAND2_X1 U2078 ( .A1(n2000), .A2(n2784), .ZN(n2280) );
  OAI22_X1 U2079 ( .A1(n2333), .A2(n2143), .B1(n1955), .B2(n2280), .ZN(n1505)
         );
  INV_X1 U2080 ( .A(n1505), .ZN(n1506) );
  NAND2_X1 U2081 ( .A1(n1507), .A2(n1506), .ZN(n1510) );
  NAND2_X1 U2082 ( .A1(n1508), .A2(n2171), .ZN(n2277) );
  INV_X1 U2083 ( .A(n3387), .ZN(n3363) );
  NOR2_X1 U2084 ( .A1(n2277), .A2(n3363), .ZN(n1826) );
  NAND2_X1 U2085 ( .A1(n1512), .A2(n1511), .ZN(n2291) );
  AND2_X1 U2086 ( .A1(n2333), .A2(n2280), .ZN(n2215) );
  INV_X1 U2087 ( .A(n1525), .ZN(n1513) );
  NAND2_X1 U2088 ( .A1(n1528), .A2(n1513), .ZN(n1517) );
  INV_X1 U2089 ( .A(n4271), .ZN(n1515) );
  AOI21_X1 U2090 ( .B1(n1515), .B2(n1528), .A(n1514), .ZN(n1516) );
  OAI21_X1 U2091 ( .B1(n1526), .B2(n1517), .A(n1516), .ZN(n1521) );
  NAND2_X1 U2092 ( .A1(n1519), .A2(n1518), .ZN(n1520) );
  XNOR2_X1 U2093 ( .A(n1521), .B(n1520), .ZN(n1523) );
  OAI22_X1 U2094 ( .A1(n1545), .A2(n2570), .B1(n1544), .B2(n4075), .ZN(n1522)
         );
  AOI21_X1 U2095 ( .B1(n1523), .B2(n82), .A(n1522), .ZN(n1966) );
  INV_X1 U2096 ( .A(n1966), .ZN(n1689) );
  NAND2_X1 U2097 ( .A1(n1321), .A2(n1689), .ZN(n1551) );
  OAI21_X1 U2098 ( .B1(n1526), .B2(n1525), .A(n4314), .ZN(n1530) );
  NAND2_X1 U2099 ( .A1(n1528), .A2(n1527), .ZN(n1529) );
  XNOR2_X1 U2100 ( .A(n1530), .B(n1529), .ZN(n1531) );
  NAND2_X1 U2101 ( .A1(n1531), .A2(n82), .ZN(n1534) );
  AOI22_X1 U2102 ( .A1(n1532), .A2(operand_a_i[9]), .B1(operand_a_i[22]), .B2(
        n91), .ZN(n1533) );
  NAND2_X1 U2103 ( .A1(n1534), .A2(n1533), .ZN(n1985) );
  NAND2_X1 U2104 ( .A1(n1821), .A2(n1985), .ZN(n1550) );
  AOI21_X1 U2105 ( .B1(n1543), .B2(n1541), .A(n1535), .ZN(n1538) );
  XOR2_X1 U2106 ( .A(n1538), .B(n1537), .Z(n1540) );
  OAI22_X1 U2107 ( .A1(n1545), .A2(n2561), .B1(n1544), .B2(n4105), .ZN(n1539)
         );
  AOI21_X1 U2108 ( .B1(n1540), .B2(n82), .A(n1539), .ZN(n1917) );
  OR2_X1 U2109 ( .A1(n1764), .A2(n1917), .ZN(n1549) );
  XNOR2_X1 U2110 ( .A(n1543), .B(n1542), .ZN(n1547) );
  INV_X1 U2111 ( .A(operand_a_i[11]), .ZN(n4069) );
  OAI22_X1 U2112 ( .A1(n1545), .A2(n4069), .B1(n1544), .B2(n4067), .ZN(n1546)
         );
  AOI21_X1 U2113 ( .B1(n1547), .B2(n82), .A(n1546), .ZN(n1919) );
  OR2_X1 U2114 ( .A1(n1751), .A2(n1919), .ZN(n1548) );
  NAND4_X1 U2115 ( .A1(n1551), .A2(n1550), .A3(n1549), .A4(n1548), .ZN(n2298)
         );
  INV_X1 U2116 ( .A(n2298), .ZN(n2142) );
  NOR2_X1 U2117 ( .A1(n2215), .A2(n2142), .ZN(n1552) );
  NAND2_X1 U2118 ( .A1(n1555), .A2(n1554), .ZN(n2420) );
  OAI21_X1 U2119 ( .B1(n1656), .B2(n2106), .A(n1566), .ZN(n1775) );
  MUX2_X1 U2120 ( .A(n1766), .B(n1676), .S(n4294), .Z(n1556) );
  NAND2_X1 U2121 ( .A1(n1557), .A2(n92), .ZN(n1558) );
  AND2_X1 U2122 ( .A1(n1566), .A2(n1558), .ZN(n1765) );
  NAND2_X1 U2123 ( .A1(n1765), .A2(n1321), .ZN(n1559) );
  AOI22_X1 U2124 ( .A1(n1260), .A2(n4272), .B1(n4282), .B2(n1647), .ZN(n1561)
         );
  INV_X1 U2125 ( .A(n1935), .ZN(n1568) );
  NOR2_X1 U2126 ( .A1(n1629), .A2(n1620), .ZN(n1767) );
  NAND2_X1 U2127 ( .A1(n1767), .A2(n2106), .ZN(n1768) );
  INV_X1 U2129 ( .A(n1562), .ZN(n1614) );
  OR2_X1 U2130 ( .A1(n1614), .A2(n1966), .ZN(n1565) );
  OR2_X1 U2131 ( .A1(n1764), .A2(n1918), .ZN(n1564) );
  OR2_X1 U2132 ( .A1(n1751), .A2(n1917), .ZN(n1563) );
  AOI21_X1 U2133 ( .B1(n2184), .B2(n92), .A(n2104), .ZN(n1567) );
  AOI21_X1 U2134 ( .B1(n1909), .B2(n1635), .A(n1567), .ZN(n1936) );
  MUX2_X1 U2135 ( .A(n1568), .B(n1936), .S(n2000), .Z(n2125) );
  INV_X1 U2136 ( .A(n2023), .ZN(n1892) );
  NAND2_X1 U2137 ( .A1(n2125), .A2(n1892), .ZN(n1627) );
  NOR2_X1 U2138 ( .A1(n2207), .A2(n2106), .ZN(n2309) );
  INV_X1 U2139 ( .A(n2013), .ZN(n1569) );
  NAND2_X1 U2140 ( .A1(n1569), .A2(n1321), .ZN(n1571) );
  OR2_X1 U2141 ( .A1(n1614), .A2(n1895), .ZN(n1570) );
  INV_X1 U2142 ( .A(n2306), .ZN(n1572) );
  NAND2_X1 U2143 ( .A1(n1587), .A2(n2230), .ZN(n2105) );
  NOR2_X1 U2144 ( .A1(n2207), .A2(n2305), .ZN(n2231) );
  AOI21_X1 U2145 ( .B1(n2309), .B2(n1572), .A(n2231), .ZN(n1624) );
  INV_X1 U2146 ( .A(n4276), .ZN(n1573) );
  OAI21_X1 U2147 ( .B1(n1573), .B2(n2106), .A(n106), .ZN(n1575) );
  NOR2_X1 U2148 ( .A1(n1635), .A2(n4294), .ZN(n1930) );
  INV_X1 U2149 ( .A(n1930), .ZN(n1815) );
  NAND2_X1 U2150 ( .A1(n1929), .A2(n92), .ZN(n1789) );
  NAND2_X1 U2151 ( .A1(n1789), .A2(n2206), .ZN(n1574) );
  AOI22_X1 U2152 ( .A1(n1575), .A2(n1815), .B1(n1574), .B2(n1620), .ZN(n1623)
         );
  INV_X1 U2153 ( .A(n1584), .ZN(n1578) );
  INV_X1 U2154 ( .A(n1868), .ZN(n1576) );
  AOI21_X1 U2155 ( .B1(n1871), .B2(n170), .A(n1576), .ZN(n1577) );
  OAI21_X1 U2156 ( .B1(n1578), .B2(n1594), .A(n1577), .ZN(n1595) );
  NAND2_X1 U2157 ( .A1(n1595), .A2(n3387), .ZN(n2314) );
  INV_X1 U2158 ( .A(n1605), .ZN(n1600) );
  AOI21_X1 U2159 ( .B1(n1871), .B2(operand_b_i[19]), .A(n1579), .ZN(n1580) );
  OAI21_X1 U2160 ( .B1(n1581), .B2(n1600), .A(n1580), .ZN(n1586) );
  OR2_X1 U2161 ( .A1(n1586), .A2(n2668), .ZN(n2024) );
  NAND2_X1 U2162 ( .A1(n1871), .A2(n4194), .ZN(n1582) );
  OAI211_X1 U2163 ( .C1(n1603), .C2(n2571), .A(n1582), .B(n1868), .ZN(n1583)
         );
  NAND2_X1 U2164 ( .A1(n2321), .A2(n1585), .ZN(n1588) );
  NAND2_X1 U2165 ( .A1(n1586), .A2(n2784), .ZN(n2017) );
  OAI211_X1 U2167 ( .C1(n2206), .C2(n2314), .A(n1588), .B(n4278), .ZN(n1803)
         );
  INV_X1 U2168 ( .A(n1606), .ZN(n1591) );
  INV_X1 U2169 ( .A(n1589), .ZN(n1864) );
  AOI21_X1 U2170 ( .B1(n1871), .B2(n4340), .A(n1864), .ZN(n1590) );
  OAI21_X1 U2171 ( .B1(n1591), .B2(n1594), .A(n1590), .ZN(n2262) );
  MUX2_X1 U2172 ( .A(n1647), .B(n1260), .S(n2262), .Z(n1787) );
  INV_X1 U2173 ( .A(n1873), .ZN(n1592) );
  AOI21_X1 U2174 ( .B1(n1871), .B2(n110), .A(n1592), .ZN(n1593) );
  OAI21_X1 U2175 ( .B1(n175), .B2(n1594), .A(n1593), .ZN(n2198) );
  MUX2_X1 U2176 ( .A(n1787), .B(n1702), .S(n2198), .Z(n2315) );
  OR2_X1 U2177 ( .A1(n1595), .A2(n3363), .ZN(n2199) );
  NOR2_X2 U2179 ( .A1(n2024), .A2(n2103), .ZN(n2323) );
  NAND2_X1 U2180 ( .A1(n1871), .A2(n4328), .ZN(n1597) );
  OAI211_X1 U2181 ( .C1(n1603), .C2(n2567), .A(n1597), .B(n1596), .ZN(n1598)
         );
  INV_X1 U2182 ( .A(n1598), .ZN(n1599) );
  NAND2_X1 U2184 ( .A1(n1702), .A2(n2120), .ZN(n1611) );
  INV_X1 U2185 ( .A(operand_b_i[8]), .ZN(n2566) );
  NAND2_X1 U2186 ( .A1(n1871), .A2(operand_b_i[16]), .ZN(n1602) );
  OAI211_X1 U2187 ( .C1(n1603), .C2(n2566), .A(n1602), .B(n1601), .ZN(n1604)
         );
  INV_X1 U2188 ( .A(n2115), .ZN(n1794) );
  INV_X1 U2189 ( .A(n1607), .ZN(n1796) );
  NOR2_X1 U2190 ( .A1(n2155), .A2(n1796), .ZN(n1609) );
  OR2_X1 U2191 ( .A1(n2120), .A2(n2115), .ZN(n2156) );
  NOR2_X1 U2192 ( .A1(n1609), .A2(n1608), .ZN(n1610) );
  NAND2_X1 U2193 ( .A1(n1611), .A2(n1610), .ZN(n1940) );
  NAND2_X1 U2194 ( .A1(n2323), .A2(n2320), .ZN(n1612) );
  OAI21_X1 U2195 ( .B1(n2315), .B2(n2199), .A(n1612), .ZN(n1613) );
  NOR2_X1 U2196 ( .A1(n1803), .A2(n1613), .ZN(n1622) );
  NAND2_X1 U2197 ( .A1(n1321), .A2(n2161), .ZN(n1618) );
  OR2_X1 U2198 ( .A1(n1614), .A2(n2027), .ZN(n1617) );
  OR2_X1 U2199 ( .A1(n1764), .A2(n2117), .ZN(n1616) );
  OR2_X1 U2200 ( .A1(n1751), .A2(n2116), .ZN(n1615) );
  MUX2_X1 U2201 ( .A(n1914), .B(n1915), .S(n1619), .Z(n2176) );
  NAND2_X1 U2202 ( .A1(n1943), .A2(n4233), .ZN(n1621) );
  OAI211_X1 U2203 ( .C1(n1624), .C2(n1623), .A(n1622), .B(n1621), .ZN(n1625)
         );
  INV_X1 U2204 ( .A(n1625), .ZN(n1626) );
  NAND2_X1 U2205 ( .A1(n1627), .A2(n1626), .ZN(n2391) );
  INV_X1 U2206 ( .A(n1766), .ZN(n1628) );
  NAND2_X1 U2207 ( .A1(n1629), .A2(n1628), .ZN(n1631) );
  NAND2_X1 U2208 ( .A1(n1636), .A2(n1731), .ZN(n1630) );
  OR2_X1 U2209 ( .A1(n1636), .A2(n1620), .ZN(n1681) );
  NOR2_X1 U2210 ( .A1(n1676), .A2(n2106), .ZN(n1777) );
  INV_X1 U2211 ( .A(n1751), .ZN(n1674) );
  NAND2_X1 U2212 ( .A1(n1765), .A2(n1674), .ZN(n1633) );
  OAI21_X1 U2213 ( .B1(n1681), .B2(n1777), .A(n1633), .ZN(n1634) );
  INV_X1 U2214 ( .A(n2171), .ZN(n1688) );
  NAND2_X1 U2215 ( .A1(n1767), .A2(n1688), .ZN(n1638) );
  NOR2_X1 U2216 ( .A1(n1636), .A2(n4294), .ZN(n1677) );
  NAND2_X1 U2217 ( .A1(n1677), .A2(n1661), .ZN(n1637) );
  NAND3_X1 U2218 ( .A1(n1768), .A2(n1638), .A3(n1637), .ZN(n1641) );
  NOR2_X1 U2219 ( .A1(n1641), .A2(n1640), .ZN(n1960) );
  NAND2_X1 U2220 ( .A1(n2089), .A2(n1892), .ZN(n1655) );
  OAI22_X1 U2221 ( .A1(n2143), .A2(n106), .B1(n2305), .B2(n2294), .ZN(n1642)
         );
  AOI21_X1 U2222 ( .B1(n1642), .B2(n92), .A(n1585), .ZN(n1893) );
  INV_X1 U2223 ( .A(n4232), .ZN(n2254) );
  NAND2_X1 U2224 ( .A1(n1930), .A2(n1824), .ZN(n1644) );
  NOR2_X1 U2225 ( .A1(n2290), .A2(n1620), .ZN(n1928) );
  NAND2_X1 U2226 ( .A1(n1928), .A2(n1713), .ZN(n1643) );
  OAI211_X1 U2227 ( .C1(n2205), .C2(n1884), .A(n1644), .B(n1643), .ZN(n2090)
         );
  NAND2_X1 U2228 ( .A1(n2090), .A2(n2309), .ZN(n1645) );
  OAI21_X1 U2229 ( .B1(n1893), .B2(n2254), .A(n1645), .ZN(n1653) );
  AND2_X1 U2230 ( .A1(n2262), .A2(n2012), .ZN(n1646) );
  OR2_X1 U2231 ( .A1(n1260), .A2(n1646), .ZN(n1703) );
  INV_X1 U2232 ( .A(n2262), .ZN(n2257) );
  MUX2_X1 U2233 ( .A(n1647), .B(n2004), .S(n2257), .Z(n2238) );
  INV_X1 U2234 ( .A(n2198), .ZN(n2193) );
  MUX2_X1 U2235 ( .A(n1703), .B(n2238), .S(n2193), .Z(n2196) );
  OR2_X1 U2236 ( .A1(n2207), .A2(n2206), .ZN(n1651) );
  INV_X1 U2237 ( .A(n2120), .ZN(n1948) );
  OAI22_X1 U2238 ( .A1(n2004), .A2(n2155), .B1(n1948), .B2(n1702), .ZN(n1649)
         );
  NAND2_X1 U2239 ( .A1(n2120), .A2(n2115), .ZN(n2160) );
  OAI22_X1 U2240 ( .A1(n1260), .A2(n2160), .B1(n2156), .B2(n1647), .ZN(n1648)
         );
  OR2_X1 U2241 ( .A1(n1649), .A2(n1648), .ZN(n2191) );
  NAND2_X1 U2242 ( .A1(n2323), .A2(n2191), .ZN(n1650) );
  OAI211_X1 U2243 ( .C1(n2196), .C2(n2199), .A(n1651), .B(n1650), .ZN(n1652)
         );
  NOR3_X1 U2244 ( .A1(n1653), .A2(n1803), .A3(n1652), .ZN(n1654) );
  NAND2_X1 U2245 ( .A1(n1655), .A2(n1654), .ZN(n2392) );
  MUX2_X1 U2246 ( .A(n1656), .B(n1676), .S(n1730), .Z(n1728) );
  MUX2_X1 U2247 ( .A(n1658), .B(n1766), .S(n1657), .Z(n1733) );
  OAI22_X1 U2248 ( .A1(n1728), .A2(n1809), .B1(n1810), .B2(n1733), .ZN(n1673)
         );
  MUX2_X1 U2249 ( .A(n2306), .B(n2304), .S(n2230), .Z(n2100) );
  NAND2_X1 U2250 ( .A1(n2171), .A2(n426), .ZN(n1659) );
  OR2_X1 U2251 ( .A1(n2290), .A2(n1659), .ZN(n2218) );
  INV_X1 U2252 ( .A(n2218), .ZN(n1660) );
  OR2_X1 U2253 ( .A1(n1660), .A2(n1930), .ZN(n1825) );
  MUX2_X1 U2254 ( .A(n1688), .B(n1661), .S(n1730), .Z(n2173) );
  NAND2_X1 U2255 ( .A1(n2173), .A2(n1620), .ZN(n1666) );
  NAND3_X1 U2256 ( .A1(n1825), .A2(n3387), .A3(n1666), .ZN(n1662) );
  OAI21_X1 U2257 ( .B1(n2254), .B2(n2100), .A(n1662), .ZN(n1665) );
  NAND2_X1 U2258 ( .A1(n1915), .A2(n426), .ZN(n2043) );
  NOR2_X1 U2259 ( .A1(n2290), .A2(n2043), .ZN(n2066) );
  OR2_X1 U2260 ( .A1(n1930), .A2(n2066), .ZN(n1828) );
  OAI21_X1 U2261 ( .B1(n2176), .B2(n4294), .A(n1828), .ZN(n1663) );
  AND2_X1 U2262 ( .A1(n2184), .A2(n1635), .ZN(n1910) );
  INV_X1 U2263 ( .A(n1910), .ZN(n1664) );
  INV_X1 U2264 ( .A(n2132), .ZN(n1669) );
  MUX2_X1 U2265 ( .A(n1985), .B(n1984), .S(n1730), .Z(n1667) );
  OAI211_X1 U2266 ( .C1(n1620), .C2(n1667), .A(n2170), .B(n1666), .ZN(n1668)
         );
  OAI21_X1 U2267 ( .B1(n1669), .B2(n2333), .A(n1668), .ZN(n2185) );
  NAND2_X1 U2268 ( .A1(n2185), .A2(n86), .ZN(n1672) );
  AOI22_X1 U2269 ( .A1(n4276), .A2(n1749), .B1(n2174), .B2(n1929), .ZN(n1670)
         );
  NAND2_X1 U2270 ( .A1(n2330), .A2(n2108), .ZN(n1671) );
  INV_X1 U2271 ( .A(n1775), .ZN(n1675) );
  AOI22_X1 U2272 ( .A1(n1675), .A2(n1674), .B1(n1765), .B2(n1821), .ZN(n1684)
         );
  NAND2_X1 U2273 ( .A1(n1677), .A2(n1676), .ZN(n1679) );
  OR2_X1 U2274 ( .A1(n1681), .A2(n1680), .ZN(n1682) );
  INV_X1 U2275 ( .A(n2329), .ZN(n2150) );
  INV_X1 U2276 ( .A(n1984), .ZN(n1687) );
  NAND2_X1 U2277 ( .A1(n1321), .A2(n1687), .ZN(n1693) );
  NAND2_X1 U2278 ( .A1(n1821), .A2(n1688), .ZN(n1692) );
  OR2_X1 U2279 ( .A1(n1764), .A2(n1689), .ZN(n1691) );
  OR2_X1 U2280 ( .A1(n1751), .A2(n1985), .ZN(n1690) );
  NAND4_X1 U2281 ( .A1(n1693), .A2(n1692), .A3(n1691), .A4(n1690), .ZN(n1860)
         );
  INV_X1 U2282 ( .A(n1917), .ZN(n1756) );
  INV_X1 U2284 ( .A(n1919), .ZN(n1694) );
  NAND2_X1 U2285 ( .A1(n1821), .A2(n1694), .ZN(n1697) );
  INV_X1 U2286 ( .A(n1914), .ZN(n1867) );
  OR2_X1 U2287 ( .A1(n1764), .A2(n1867), .ZN(n1696) );
  OR2_X1 U2288 ( .A1(n1751), .A2(n1918), .ZN(n1695) );
  NAND4_X1 U2289 ( .A1(n1698), .A2(n1697), .A3(n1696), .A4(n1695), .ZN(n1820)
         );
  NAND2_X1 U2290 ( .A1(n1820), .A2(n2105), .ZN(n1699) );
  OAI21_X1 U2291 ( .B1(n106), .B2(n1860), .A(n1699), .ZN(n1700) );
  NAND2_X1 U2292 ( .A1(n1700), .A2(n92), .ZN(n1701) );
  NAND2_X1 U2293 ( .A1(n1701), .A2(n2206), .ZN(n2060) );
  OAI21_X1 U2294 ( .B1(n2155), .B2(n1260), .A(n1702), .ZN(n2239) );
  OAI21_X1 U2295 ( .B1(n2323), .B2(n426), .A(n2239), .ZN(n1706) );
  INV_X1 U2296 ( .A(n2199), .ZN(n1704) );
  AOI21_X1 U2297 ( .B1(n1702), .B2(n2198), .A(n1703), .ZN(n2240) );
  NAND2_X1 U2298 ( .A1(n1704), .A2(n2240), .ZN(n1705) );
  NAND2_X1 U2299 ( .A1(n1706), .A2(n1705), .ZN(n1707) );
  INV_X1 U2300 ( .A(n1824), .ZN(n1709) );
  MUX2_X1 U2301 ( .A(n1709), .B(n1708), .S(n1620), .Z(n1710) );
  OAI21_X1 U2302 ( .B1(n1710), .B2(n2106), .A(n2206), .ZN(n2229) );
  OR2_X1 U2303 ( .A1(n1751), .A2(n1944), .ZN(n1712) );
  OR2_X1 U2304 ( .A1(n1764), .A2(n1796), .ZN(n1711) );
  OAI21_X1 U2305 ( .B1(n2052), .B2(n2106), .A(n106), .ZN(n1714) );
  OAI211_X1 U2306 ( .C1(n2229), .C2(n86), .A(n2108), .B(n1714), .ZN(n1725) );
  NAND2_X1 U2307 ( .A1(n1715), .A2(n1620), .ZN(n1719) );
  OR2_X1 U2308 ( .A1(n1751), .A2(n1716), .ZN(n1718) );
  OR2_X1 U2309 ( .A1(n1764), .A2(n2027), .ZN(n1717) );
  AND3_X1 U2310 ( .A1(n1719), .A2(n1718), .A3(n1717), .ZN(n2048) );
  AOI21_X1 U2311 ( .B1(n2048), .B2(n92), .A(n1585), .ZN(n2084) );
  NAND2_X1 U2312 ( .A1(n4272), .A2(n2158), .ZN(n1723) );
  NAND2_X1 U2313 ( .A1(n1821), .A2(n2161), .ZN(n1722) );
  OR2_X1 U2314 ( .A1(n1764), .A2(n1895), .ZN(n1721) );
  OR2_X1 U2315 ( .A1(n1751), .A2(n2117), .ZN(n1720) );
  NAND2_X1 U2316 ( .A1(n2002), .A2(n4233), .ZN(n1724) );
  NAND4_X1 U2317 ( .A1(n1727), .A2(n1726), .A3(n1725), .A4(n1724), .ZN(n2390)
         );
  MUX2_X1 U2318 ( .A(n2173), .B(n1728), .S(n1620), .Z(n2216) );
  MUX2_X1 U2319 ( .A(n1731), .B(n1560), .S(n1730), .Z(n1732) );
  NAND2_X1 U2320 ( .A1(n2174), .A2(n1732), .ZN(n1736) );
  INV_X1 U2321 ( .A(n1733), .ZN(n1734) );
  NAND2_X1 U2322 ( .A1(n1749), .A2(n1734), .ZN(n1735) );
  OAI211_X1 U2323 ( .C1(n2216), .C2(n2230), .A(n1736), .B(n1735), .ZN(n1737)
         );
  OR2_X1 U2324 ( .A1(n1751), .A2(n2027), .ZN(n1740) );
  INV_X1 U2325 ( .A(n1764), .ZN(n1738) );
  NAND2_X1 U2326 ( .A1(n1738), .A2(n2161), .ZN(n1739) );
  OAI211_X1 U2327 ( .C1(n1741), .C2(n4294), .A(n1740), .B(n1739), .ZN(n2270)
         );
  INV_X1 U2328 ( .A(n2270), .ZN(n2220) );
  NAND2_X1 U2329 ( .A1(n1321), .A2(n2077), .ZN(n1745) );
  NAND2_X1 U2330 ( .A1(n1821), .A2(n2158), .ZN(n1744) );
  OR2_X1 U2331 ( .A1(n1764), .A2(n2013), .ZN(n1743) );
  OR2_X1 U2332 ( .A1(n1751), .A2(n1895), .ZN(n1742) );
  INV_X1 U2333 ( .A(n164), .ZN(n1746) );
  OR2_X1 U2334 ( .A1(n1751), .A2(n1796), .ZN(n1748) );
  OR2_X1 U2335 ( .A1(n1764), .A2(n1795), .ZN(n1747) );
  OAI211_X1 U2336 ( .C1(n1927), .C2(n4294), .A(n1748), .B(n1747), .ZN(n1771)
         );
  AOI22_X1 U2337 ( .A1(n1929), .A2(n1749), .B1(n2174), .B2(n1838), .ZN(n1750)
         );
  AOI22_X1 U2338 ( .A1(n4233), .A2(n2033), .B1(n2108), .B2(n2267), .ZN(n1763)
         );
  INV_X1 U2339 ( .A(n2215), .ZN(n1761) );
  NAND2_X1 U2340 ( .A1(n1321), .A2(n1985), .ZN(n1755) );
  NAND2_X1 U2341 ( .A1(n1821), .A2(n1984), .ZN(n1754) );
  OR2_X1 U2342 ( .A1(n1764), .A2(n1919), .ZN(n1753) );
  OR2_X1 U2343 ( .A1(n1751), .A2(n1966), .ZN(n1752) );
  NAND4_X1 U2344 ( .A1(n1755), .A2(n1754), .A3(n1753), .A4(n1752), .ZN(n2221)
         );
  NAND2_X1 U2345 ( .A1(n1821), .A2(n1756), .ZN(n1760) );
  NAND2_X1 U2346 ( .A1(n1321), .A2(n1757), .ZN(n1759) );
  NAND2_X1 U2347 ( .A1(n2176), .A2(n4294), .ZN(n1758) );
  INV_X1 U2349 ( .A(n2214), .ZN(n2064) );
  MUX2_X1 U2350 ( .A(n2221), .B(n2064), .S(n86), .Z(n1995) );
  NAND2_X1 U2351 ( .A1(n1761), .A2(n1995), .ZN(n1762) );
  AOI22_X1 U2352 ( .A1(n1767), .A2(n1766), .B1(n1765), .B2(n1738), .ZN(n1769)
         );
  INV_X1 U2353 ( .A(n1977), .ZN(n1773) );
  NAND2_X1 U2354 ( .A1(n1771), .A2(n2290), .ZN(n1772) );
  OAI21_X1 U2355 ( .B1(n1773), .B2(n2230), .A(n1772), .ZN(n1842) );
  INV_X1 U2356 ( .A(n1776), .ZN(n1779) );
  NOR2_X1 U2357 ( .A1(n4294), .A2(n1777), .ZN(n1778) );
  NAND2_X1 U2358 ( .A1(n1779), .A2(n1778), .ZN(n1780) );
  AOI21_X1 U2359 ( .B1(n2221), .B2(n92), .A(n2104), .ZN(n1783) );
  AOI21_X1 U2360 ( .B1(n1978), .B2(n1635), .A(n1783), .ZN(n1843) );
  NAND2_X1 U2361 ( .A1(n1843), .A2(n2000), .ZN(n1784) );
  OAI21_X1 U2362 ( .B1(n2000), .B2(n1842), .A(n1784), .ZN(n2063) );
  NAND2_X1 U2363 ( .A1(n4281), .A2(n1892), .ZN(n1807) );
  OAI22_X1 U2364 ( .A1(n2214), .A2(n106), .B1(n2305), .B2(n2270), .ZN(n1785)
         );
  NAND2_X1 U2365 ( .A1(n1785), .A2(n92), .ZN(n1786) );
  NAND2_X1 U2366 ( .A1(n1786), .A2(n2206), .ZN(n1844) );
  AND2_X1 U2367 ( .A1(n1844), .A2(n4233), .ZN(n1805) );
  MUX2_X1 U2368 ( .A(n2003), .B(n2004), .S(n2262), .Z(n2316) );
  MUX2_X1 U2369 ( .A(n1787), .B(n2316), .S(n2193), .Z(n2265) );
  NAND3_X1 U2370 ( .A1(n106), .A2(n1789), .A3(n4294), .ZN(n1793) );
  OAI21_X1 U2371 ( .B1(n164), .B2(n2106), .A(n2305), .ZN(n1792) );
  NAND2_X1 U2372 ( .A1(n1838), .A2(n92), .ZN(n1790) );
  NAND3_X1 U2373 ( .A1(n1930), .A2(n2206), .A3(n1790), .ZN(n1791) );
  NAND4_X1 U2374 ( .A1(n2108), .A2(n1793), .A3(n1792), .A4(n1791), .ZN(n1802)
         );
  OR2_X1 U2375 ( .A1(n2156), .A2(n1944), .ZN(n1800) );
  NAND2_X1 U2376 ( .A1(n2120), .A2(n1794), .ZN(n2159) );
  OR2_X1 U2377 ( .A1(n2159), .A2(n1795), .ZN(n1798) );
  OR2_X1 U2378 ( .A1(n2160), .A2(n1796), .ZN(n1797) );
  NAND2_X1 U2379 ( .A1(n2323), .A2(n2269), .ZN(n1801) );
  OAI211_X1 U2380 ( .C1(n2265), .C2(n2199), .A(n1802), .B(n1801), .ZN(n1804)
         );
  NOR3_X1 U2381 ( .A1(n1805), .A2(n1804), .A3(n1803), .ZN(n1806) );
  NAND2_X1 U2382 ( .A1(n1807), .A2(n1806), .ZN(n2393) );
  OAI22_X1 U2383 ( .A1(n1811), .A2(n1810), .B1(n1809), .B2(n1808), .ZN(n1837)
         );
  INV_X1 U2384 ( .A(n2048), .ZN(n1885) );
  INV_X1 U2385 ( .A(n1860), .ZN(n1812) );
  NAND2_X1 U2386 ( .A1(n2170), .A2(n1812), .ZN(n1813) );
  OAI21_X1 U2387 ( .B1(n1885), .B2(n2333), .A(n1813), .ZN(n2285) );
  NAND2_X1 U2388 ( .A1(n2285), .A2(n1884), .ZN(n1835) );
  OAI22_X1 U2389 ( .A1(n2052), .A2(n1884), .B1(n1815), .B2(n1814), .ZN(n1816)
         );
  INV_X1 U2390 ( .A(n1816), .ZN(n1819) );
  INV_X1 U2391 ( .A(n1928), .ZN(n1817) );
  NAND2_X1 U2392 ( .A1(n1819), .A2(n475), .ZN(n2234) );
  NAND2_X1 U2393 ( .A1(n1820), .A2(n2290), .ZN(n1829) );
  INV_X1 U2394 ( .A(n1829), .ZN(n1863) );
  AOI22_X1 U2395 ( .A1(n2234), .A2(n2108), .B1(n4287), .B2(n1863), .ZN(n1834)
         );
  INV_X1 U2396 ( .A(n2009), .ZN(n2258) );
  NAND2_X1 U2397 ( .A1(n2258), .A2(n4272), .ZN(n1823) );
  NAND2_X1 U2398 ( .A1(n4282), .A2(n1569), .ZN(n1822) );
  OAI211_X1 U2399 ( .C1(n1824), .C2(n1620), .A(n1823), .B(n1822), .ZN(n2047)
         );
  MUX2_X1 U2400 ( .A(n2047), .B(n2228), .S(n2230), .Z(n1882) );
  INV_X1 U2401 ( .A(n1882), .ZN(n2082) );
  AOI22_X1 U2402 ( .A1(n2082), .A2(n4233), .B1(n1826), .B2(n1825), .ZN(n1833)
         );
  INV_X1 U2403 ( .A(n1827), .ZN(n2046) );
  NAND2_X1 U2404 ( .A1(n1828), .A2(n2046), .ZN(n1830) );
  NAND2_X1 U2405 ( .A1(n1830), .A2(n1829), .ZN(n1858) );
  INV_X1 U2406 ( .A(n2280), .ZN(n1831) );
  NAND2_X1 U2407 ( .A1(n1858), .A2(n1831), .ZN(n1832) );
  NAND2_X1 U2408 ( .A1(n1930), .A2(n1838), .ZN(n1840) );
  NAND2_X1 U2409 ( .A1(n1928), .A2(n1929), .ZN(n1839) );
  OAI211_X1 U2410 ( .C1(n164), .C2(n1884), .A(n1840), .B(n1839), .ZN(n1841) );
  NAND2_X1 U2412 ( .A1(n1843), .A2(n4233), .ZN(n1856) );
  NAND2_X1 U2413 ( .A1(n1844), .A2(n2108), .ZN(n1855) );
  AND2_X1 U2414 ( .A1(n4231), .A2(n3387), .ZN(n1845) );
  OAI22_X1 U2416 ( .A1(n1895), .A2(n2160), .B1(n2159), .B2(n2013), .ZN(n1847)
         );
  OAI22_X1 U2417 ( .A1(n2116), .A2(n2155), .B1(n2156), .B2(n2117), .ZN(n1846)
         );
  NOR2_X1 U2418 ( .A1(n1847), .A2(n1846), .ZN(n2025) );
  INV_X1 U2419 ( .A(n2236), .ZN(n1848) );
  NOR2_X1 U2420 ( .A1(n2012), .A2(n3363), .ZN(n2172) );
  NAND2_X1 U2421 ( .A1(n2013), .A2(n2172), .ZN(n1941) );
  NOR2_X1 U2422 ( .A1(n4231), .A2(n1941), .ZN(n2118) );
  AOI21_X1 U2423 ( .B1(n1848), .B2(n2103), .A(n2118), .ZN(n1949) );
  NOR2_X1 U2424 ( .A1(n2017), .A2(n2103), .ZN(n2146) );
  OAI22_X1 U2425 ( .A1(n4298), .A2(n2160), .B1(n2159), .B2(n2194), .ZN(n1850)
         );
  OAI22_X1 U2426 ( .A1(n2256), .A2(n2156), .B1(n2155), .B2(n2009), .ZN(n1849)
         );
  NOR2_X1 U2427 ( .A1(n1850), .A2(n1849), .ZN(n2268) );
  AOI22_X1 U2428 ( .A1(n2269), .A2(n2146), .B1(n2321), .B2(n2268), .ZN(n1851)
         );
  NAND2_X1 U2429 ( .A1(n1949), .A2(n1851), .ZN(n1852) );
  AND3_X1 U2430 ( .A1(n1855), .A2(n1856), .A3(n1854), .ZN(n1857) );
  OAI21_X1 U2431 ( .B1(n2227), .B2(n2023), .A(n1857), .ZN(n2401) );
  AOI22_X1 U2432 ( .A1(n2234), .A2(n4233), .B1(n2130), .B2(n1858), .ZN(n1889)
         );
  OAI21_X1 U2433 ( .B1(n1860), .B2(n2106), .A(n106), .ZN(n1861) );
  INV_X1 U2434 ( .A(n1861), .ZN(n1862) );
  AOI21_X1 U2435 ( .B1(n1859), .B2(n2290), .A(n1862), .ZN(n2233) );
  AOI22_X1 U2436 ( .A1(n2233), .A2(n2108), .B1(n2329), .B2(n1863), .ZN(n1888)
         );
  AOI21_X1 U2437 ( .B1(n1872), .B2(operand_b_i[16]), .A(n1864), .ZN(n1866) );
  NAND2_X1 U2438 ( .A1(n1871), .A2(n4196), .ZN(n1865) );
  AND2_X1 U2439 ( .A1(n1866), .A2(n1865), .ZN(n1983) );
  MUX2_X1 U2440 ( .A(n1867), .B(n1918), .S(n1983), .Z(n1964) );
  NAND2_X1 U2441 ( .A1(n1871), .A2(operand_b_i[10]), .ZN(n1870) );
  NAND2_X1 U2442 ( .A1(n1872), .A2(n4194), .ZN(n1869) );
  NAND3_X1 U2443 ( .A1(n1870), .A2(n1869), .A3(n1868), .ZN(n1878) );
  NOR2_X1 U2444 ( .A1(n1878), .A2(n3363), .ZN(n2129) );
  NAND2_X1 U2445 ( .A1(n1871), .A2(n4195), .ZN(n1875) );
  NAND2_X1 U2446 ( .A1(n1872), .A2(n4328), .ZN(n1874) );
  NAND3_X1 U2447 ( .A1(n1875), .A2(n1874), .A3(n1873), .ZN(n1963) );
  NAND2_X1 U2448 ( .A1(n2129), .A2(n1963), .ZN(n1989) );
  INV_X1 U2449 ( .A(n1983), .ZN(n1965) );
  MUX2_X1 U2450 ( .A(n1919), .B(n1917), .S(n1965), .Z(n1969) );
  INV_X1 U2451 ( .A(n1963), .ZN(n1982) );
  NAND2_X1 U2452 ( .A1(n2129), .A2(n1982), .ZN(n1987) );
  OAI22_X1 U2453 ( .A1(n1964), .A2(n1989), .B1(n1969), .B2(n1987), .ZN(n1880)
         );
  NAND2_X1 U2454 ( .A1(n2043), .A2(n1963), .ZN(n1877) );
  NAND2_X1 U2455 ( .A1(n1965), .A2(n2012), .ZN(n1876) );
  AND2_X1 U2456 ( .A1(n1915), .A2(n1876), .ZN(n1961) );
  NAND2_X1 U2457 ( .A1(n1877), .A2(n1961), .ZN(n2055) );
  NAND2_X1 U2458 ( .A1(n1878), .A2(n3387), .ZN(n1913) );
  NOR2_X1 U2459 ( .A1(n2055), .A2(n1913), .ZN(n1879) );
  NOR2_X1 U2460 ( .A1(n1880), .A2(n1879), .ZN(n1881) );
  OR2_X1 U2461 ( .A1(n2280), .A2(n2043), .ZN(n2219) );
  OAI211_X1 U2462 ( .C1(n1882), .C2(n2333), .A(n1881), .B(n2219), .ZN(n1883)
         );
  INV_X1 U2463 ( .A(n1883), .ZN(n1887) );
  NAND2_X1 U2464 ( .A1(n2329), .A2(n1884), .ZN(n2137) );
  OR2_X1 U2465 ( .A1(n2137), .A2(n1885), .ZN(n1886) );
  NAND4_X1 U2466 ( .A1(n1889), .A2(n1888), .A3(n1887), .A4(n1886), .ZN(n2410)
         );
  NAND2_X1 U2467 ( .A1(n2090), .A2(n1933), .ZN(n1891) );
  OAI22_X1 U2468 ( .A1(n4292), .A2(n2254), .B1(n1893), .B2(n2207), .ZN(n1905)
         );
  INV_X1 U2469 ( .A(n2017), .ZN(n2035) );
  MUX2_X1 U2470 ( .A(n1895), .B(n2117), .S(n2115), .Z(n1896) );
  NAND2_X1 U2471 ( .A1(n1896), .A2(n1948), .ZN(n1901) );
  OAI211_X1 U2472 ( .C1(n426), .C2(n2115), .A(n2120), .B(n2013), .ZN(n1897) );
  AOI21_X1 U2473 ( .B1(n1901), .B2(n1897), .A(n3363), .ZN(n1898) );
  AOI21_X1 U2474 ( .B1(n2035), .B2(n2191), .A(n1898), .ZN(n2152) );
  OAI22_X1 U2475 ( .A1(n4298), .A2(n2156), .B1(n2155), .B2(n2256), .ZN(n1899)
         );
  NOR2_X1 U2476 ( .A1(n1900), .A2(n1899), .ZN(n2190) );
  MUX2_X1 U2477 ( .A(n2258), .B(n1569), .S(n2115), .Z(n1902) );
  OAI21_X1 U2478 ( .B1(n1902), .B2(n1948), .A(n1901), .ZN(n2145) );
  AOI22_X1 U2479 ( .A1(n2321), .A2(n2190), .B1(n2323), .B2(n2145), .ZN(n1903)
         );
  OAI211_X1 U2480 ( .C1(n2152), .C2(n2103), .A(n1949), .B(n1903), .ZN(n1904)
         );
  NOR2_X1 U2481 ( .A1(n1905), .A2(n1904), .ZN(n1906) );
  NAND2_X1 U2482 ( .A1(n1907), .A2(n1906), .ZN(n2400) );
  MUX2_X1 U2483 ( .A(n1909), .B(n1908), .S(n1635), .Z(n2334) );
  INV_X1 U2484 ( .A(n2130), .ZN(n2068) );
  NAND2_X1 U2485 ( .A1(n2329), .A2(n1910), .ZN(n1911) );
  OAI21_X1 U2486 ( .B1(n1912), .B2(n2068), .A(n1911), .ZN(n1923) );
  INV_X1 U2487 ( .A(n1913), .ZN(n2044) );
  MUX2_X1 U2488 ( .A(n1915), .B(n1914), .S(n1983), .Z(n1981) );
  NAND2_X1 U2489 ( .A1(n1981), .A2(n1982), .ZN(n1916) );
  OAI21_X1 U2490 ( .B1(n1982), .B2(n2043), .A(n1916), .ZN(n2128) );
  MUX2_X1 U2491 ( .A(n1918), .B(n1917), .S(n1983), .Z(n1979) );
  MUX2_X1 U2492 ( .A(n1919), .B(n1966), .S(n1983), .Z(n1990) );
  OAI22_X1 U2493 ( .A1(n1979), .A2(n1989), .B1(n1990), .B2(n1987), .ZN(n1920)
         );
  AOI21_X1 U2494 ( .B1(n2044), .B2(n2128), .A(n1920), .ZN(n1921) );
  OAI211_X1 U2495 ( .C1(n2100), .C2(n2333), .A(n1921), .B(n2219), .ZN(n1922)
         );
  NOR2_X1 U2496 ( .A1(n1923), .A2(n1922), .ZN(n1926) );
  INV_X1 U2497 ( .A(n2137), .ZN(n1924) );
  AOI22_X1 U2498 ( .A1(n2330), .A2(n4233), .B1(n1924), .B2(n2132), .ZN(n1925)
         );
  NAND2_X1 U2499 ( .A1(n1928), .A2(n4276), .ZN(n1932) );
  OAI211_X1 U2501 ( .C1(n2306), .C2(n1884), .A(n1932), .B(n1931), .ZN(n2126)
         );
  INV_X1 U2502 ( .A(n2126), .ZN(n1934) );
  NAND2_X1 U2503 ( .A1(n1936), .A2(n4233), .ZN(n1954) );
  OR2_X1 U2504 ( .A1(n2155), .A2(n2076), .ZN(n1937) );
  NAND2_X1 U2505 ( .A1(n1938), .A2(n3387), .ZN(n1939) );
  OAI21_X1 U2506 ( .B1(n1940), .B2(n2017), .A(n1939), .ZN(n2102) );
  NOR2_X1 U2507 ( .A1(n1948), .A2(n1941), .ZN(n1942) );
  OAI21_X1 U2508 ( .B1(n2102), .B2(n1942), .A(n4231), .ZN(n1952) );
  NAND2_X1 U2509 ( .A1(n1943), .A2(n2108), .ZN(n1951) );
  OAI22_X1 U2510 ( .A1(n4298), .A2(n2155), .B1(n2156), .B2(n157), .ZN(n1945)
         );
  NOR2_X1 U2511 ( .A1(n1946), .A2(n1945), .ZN(n2322) );
  INV_X1 U2512 ( .A(n2143), .ZN(n1957) );
  INV_X1 U2513 ( .A(n1955), .ZN(n1956) );
  AOI22_X1 U2514 ( .A1(n2329), .A2(n1957), .B1(n1956), .B2(n2130), .ZN(n2098)
         );
  NAND2_X1 U2515 ( .A1(n2170), .A2(n2298), .ZN(n1958) );
  MUX2_X1 U2516 ( .A(n2098), .B(n1958), .S(n2230), .Z(n1976) );
  MUX2_X1 U2517 ( .A(n1960), .B(n1959), .S(n2290), .Z(n2189) );
  NAND2_X1 U2518 ( .A1(n2189), .A2(n2108), .ZN(n1975) );
  NAND2_X1 U2519 ( .A1(n1961), .A2(n1963), .ZN(n1962) );
  OAI21_X1 U2520 ( .B1(n1964), .B2(n1963), .A(n1962), .ZN(n2091) );
  INV_X1 U2521 ( .A(n1985), .ZN(n1967) );
  MUX2_X1 U2522 ( .A(n1967), .B(n1966), .S(n1965), .Z(n1968) );
  OAI22_X1 U2523 ( .A1(n1969), .A2(n1989), .B1(n1968), .B2(n1987), .ZN(n1970)
         );
  AOI21_X1 U2524 ( .B1(n2091), .B2(n2044), .A(n1970), .ZN(n1971) );
  OAI211_X1 U2525 ( .C1(n2149), .C2(n2333), .A(n1971), .B(n2219), .ZN(n1972)
         );
  INV_X1 U2526 ( .A(n1972), .ZN(n1974) );
  NAND2_X1 U2527 ( .A1(n2192), .A2(n4233), .ZN(n1973) );
  NAND4_X1 U2528 ( .A1(n1976), .A2(n1975), .A3(n1974), .A4(n1973), .ZN(n2412)
         );
  NAND2_X1 U2529 ( .A1(n2267), .A2(n4233), .ZN(n1998) );
  NAND2_X1 U2530 ( .A1(n4287), .A2(n2033), .ZN(n1997) );
  NAND2_X1 U2531 ( .A1(n1979), .A2(n1982), .ZN(n1980) );
  OAI21_X1 U2532 ( .B1(n1982), .B2(n1981), .A(n1980), .ZN(n2069) );
  INV_X1 U2533 ( .A(n2069), .ZN(n1992) );
  MUX2_X1 U2534 ( .A(n1985), .B(n1984), .S(n1983), .Z(n1986) );
  INV_X1 U2535 ( .A(n1986), .ZN(n1988) );
  OAI22_X1 U2536 ( .A1(n1990), .A2(n1989), .B1(n1988), .B2(n1987), .ZN(n1991)
         );
  AOI21_X1 U2537 ( .B1(n1992), .B2(n2044), .A(n1991), .ZN(n1993) );
  NAND2_X1 U2538 ( .A1(n2219), .A2(n1993), .ZN(n1994) );
  OAI21_X1 U2539 ( .B1(n2275), .B2(n2207), .A(n1999), .ZN(n2413) );
  OR2_X1 U2541 ( .A1(n2156), .A2(n2003), .ZN(n2008) );
  INV_X1 U2542 ( .A(n2194), .ZN(n2263) );
  OR2_X1 U2543 ( .A1(n2263), .A2(n2155), .ZN(n2007) );
  OR2_X1 U2544 ( .A1(n2159), .A2(n1647), .ZN(n2006) );
  OR2_X1 U2545 ( .A1(n2004), .A2(n2160), .ZN(n2005) );
  NAND4_X1 U2546 ( .A1(n2008), .A2(n2007), .A3(n2006), .A4(n2005), .ZN(n2235)
         );
  OAI22_X1 U2547 ( .A1(n4298), .A2(n2159), .B1(n2160), .B2(n2256), .ZN(n2011)
         );
  OAI22_X1 U2548 ( .A1(n2009), .A2(n2156), .B1(n2155), .B2(n2013), .ZN(n2010)
         );
  NOR2_X1 U2549 ( .A1(n2011), .A2(n2010), .ZN(n2073) );
  AOI22_X1 U2550 ( .A1(n2321), .A2(n2235), .B1(n2323), .B2(n2073), .ZN(n2020)
         );
  NAND2_X1 U2551 ( .A1(n2060), .A2(n4233), .ZN(n2019) );
  INV_X1 U2552 ( .A(n2239), .ZN(n2016) );
  NAND2_X1 U2553 ( .A1(n2155), .A2(n2012), .ZN(n2014) );
  NAND3_X1 U2554 ( .A1(n2014), .A2(n3387), .A3(n2013), .ZN(n2015) );
  OAI21_X1 U2555 ( .B1(n2017), .B2(n2016), .A(n2015), .ZN(n2081) );
  OAI21_X1 U2556 ( .B1(n426), .B2(n4231), .A(n2081), .ZN(n2018) );
  AND4_X1 U2557 ( .A1(n2019), .A2(n2020), .A3(n2021), .A4(n2018), .ZN(n2022)
         );
  NAND2_X1 U2558 ( .A1(n2024), .A2(n3363), .ZN(n2026) );
  AND2_X1 U2559 ( .A1(n2026), .A2(n2025), .ZN(n2032) );
  MUX2_X1 U2560 ( .A(n2028), .B(n2027), .S(n2115), .Z(n2114) );
  NAND2_X1 U2561 ( .A1(n2114), .A2(n2120), .ZN(n2029) );
  OAI21_X1 U2562 ( .B1(n180), .B2(n2155), .A(n2029), .ZN(n2031) );
  OAI21_X1 U2563 ( .B1(n2154), .B2(n2156), .A(n4231), .ZN(n2030) );
  OAI22_X1 U2564 ( .A1(n2162), .A2(n2032), .B1(n2031), .B2(n2030), .ZN(n2041)
         );
  AOI22_X1 U2565 ( .A1(n2329), .A2(n2033), .B1(n4287), .B2(n2267), .ZN(n2040)
         );
  AOI22_X1 U2566 ( .A1(n2146), .A2(n2268), .B1(n2035), .B2(n2034), .ZN(n2039)
         );
  NAND2_X1 U2567 ( .A1(n2221), .A2(n2104), .ZN(n2036) );
  OAI21_X1 U2568 ( .B1(n2214), .B2(n2305), .A(n2036), .ZN(n2037) );
  AOI21_X1 U2569 ( .B1(n2037), .B2(n92), .A(n1585), .ZN(n2255) );
  OR2_X1 U2570 ( .A1(n2255), .A2(n2207), .ZN(n2038) );
  AND4_X1 U2571 ( .A1(n2040), .A2(n2041), .A3(n2039), .A4(n2038), .ZN(n2042)
         );
  INV_X1 U2572 ( .A(n2043), .ZN(n2127) );
  NAND2_X1 U2573 ( .A1(n2127), .A2(n2044), .ZN(n2045) );
  AND2_X1 U2574 ( .A1(n2219), .A2(n2045), .ZN(n2135) );
  AND2_X1 U2575 ( .A1(n2135), .A2(n2068), .ZN(n2051) );
  OAI21_X1 U2576 ( .B1(n2174), .B2(n2127), .A(n2046), .ZN(n2279) );
  INV_X1 U2577 ( .A(n2047), .ZN(n2049) );
  AOI22_X1 U2578 ( .A1(n85), .A2(n2049), .B1(n2329), .B2(n2048), .ZN(n2050) );
  OAI22_X1 U2579 ( .A1(n2051), .A2(n2279), .B1(n2050), .B2(n1884), .ZN(n2054)
         );
  INV_X1 U2581 ( .A(n2052), .ZN(n2053) );
  OR2_X1 U2582 ( .A1(n2137), .A2(n2228), .ZN(n2057) );
  INV_X1 U2583 ( .A(n2129), .ZN(n2092) );
  OR2_X1 U2584 ( .A1(n2055), .A2(n2092), .ZN(n2056) );
  OAI211_X1 U2585 ( .C1(n2058), .C2(n2254), .A(n2057), .B(n2056), .ZN(n2059)
         );
  INV_X1 U2586 ( .A(n2059), .ZN(n2061) );
  NAND3_X1 U2587 ( .A1(n2062), .A2(n2061), .A3(n463), .ZN(n2406) );
  INV_X1 U2588 ( .A(n2288), .ZN(n2292) );
  NAND3_X1 U2589 ( .A1(n2170), .A2(n1635), .A3(n2064), .ZN(n2065) );
  OAI21_X1 U2590 ( .B1(n2137), .B2(n2270), .A(n2065), .ZN(n2071) );
  INV_X1 U2591 ( .A(n2066), .ZN(n2067) );
  OAI21_X1 U2592 ( .B1(n2068), .B2(n2067), .A(n2135), .ZN(n2097) );
  AOI22_X1 U2593 ( .A1(n2146), .A2(n2235), .B1(n2321), .B2(n2073), .ZN(n2074)
         );
  OAI22_X1 U2594 ( .A1(n2077), .A2(n2160), .B1(n2159), .B2(n2076), .ZN(n2079)
         );
  OAI22_X1 U2595 ( .A1(n2161), .A2(n2155), .B1(n2156), .B2(n2158), .ZN(n2078)
         );
  OR2_X1 U2596 ( .A1(n2079), .A2(n2078), .ZN(n2080) );
  AOI22_X1 U2597 ( .A1(n4288), .A2(n2234), .B1(n2162), .B2(n2080), .ZN(n2087)
         );
  AOI22_X1 U2598 ( .A1(n2082), .A2(n2329), .B1(n2103), .B2(n2081), .ZN(n2086)
         );
  AOI21_X1 U2599 ( .B1(n1820), .B2(n92), .A(n2105), .ZN(n2083) );
  AOI21_X1 U2600 ( .B1(n2084), .B2(n1884), .A(n2083), .ZN(n2248) );
  NAND2_X1 U2601 ( .A1(n2248), .A2(n2108), .ZN(n2085) );
  NAND4_X1 U2602 ( .A1(n2088), .A2(n2087), .A3(n2086), .A4(n2085), .ZN(n2402)
         );
  NOR2_X1 U2603 ( .A1(n2137), .A2(n2294), .ZN(n2096) );
  INV_X1 U2604 ( .A(n2090), .ZN(n2094) );
  INV_X1 U2605 ( .A(n2091), .ZN(n2093) );
  OAI22_X1 U2606 ( .A1(n2094), .A2(n2333), .B1(n2093), .B2(n2092), .ZN(n2095)
         );
  NOR3_X1 U2607 ( .A1(n2095), .A2(n2096), .A3(n2097), .ZN(n2099) );
  NAND2_X1 U2608 ( .A1(n2330), .A2(n4288), .ZN(n2113) );
  INV_X1 U2609 ( .A(n2100), .ZN(n2101) );
  AOI22_X1 U2610 ( .A1(n2103), .A2(n2102), .B1(n2329), .B2(n2101), .ZN(n2112)
         );
  AOI22_X1 U2611 ( .A1(n2132), .A2(n2105), .B1(n2184), .B2(n2104), .ZN(n2107)
         );
  OAI21_X1 U2612 ( .B1(n2107), .B2(n2106), .A(n2206), .ZN(n2311) );
  NAND2_X1 U2613 ( .A1(n2311), .A2(n2108), .ZN(n2111) );
  AOI22_X1 U2614 ( .A1(n2322), .A2(n2146), .B1(n2321), .B2(n2109), .ZN(n2110)
         );
  AND4_X1 U2615 ( .A1(n2112), .A2(n2113), .A3(n2111), .A4(n2110), .ZN(n2124)
         );
  NAND2_X1 U2616 ( .A1(n2162), .A2(n2114), .ZN(n2122) );
  MUX2_X1 U2617 ( .A(n2117), .B(n2116), .S(n2115), .Z(n2119) );
  AOI21_X1 U2618 ( .B1(n2162), .B2(n2119), .A(n2118), .ZN(n2121) );
  MUX2_X1 U2619 ( .A(n2122), .B(n2121), .S(n2120), .Z(n2123) );
  OAI211_X1 U2620 ( .C1(n2334), .C2(n2254), .A(n2124), .B(n2123), .ZN(n2403)
         );
  NAND2_X1 U2622 ( .A1(n4287), .A2(n2126), .ZN(n2136) );
  AOI22_X1 U2623 ( .A1(n2131), .A2(n2130), .B1(n2129), .B2(n2128), .ZN(n2134)
         );
  NAND3_X1 U2624 ( .A1(n2329), .A2(n2290), .A3(n2132), .ZN(n2133) );
  NAND4_X1 U2625 ( .A1(n2136), .A2(n2135), .A3(n2134), .A4(n2133), .ZN(n2139)
         );
  NOR2_X1 U2626 ( .A1(n2137), .A2(n2304), .ZN(n2138) );
  NOR2_X1 U2627 ( .A1(n2139), .A2(n2138), .ZN(n2140) );
  OAI22_X1 U2628 ( .A1(n2143), .A2(n2305), .B1(n106), .B2(n2142), .ZN(n2144)
         );
  AOI21_X1 U2629 ( .B1(n2144), .B2(n92), .A(n1585), .ZN(n2209) );
  AOI22_X1 U2630 ( .A1(n2190), .A2(n2146), .B1(n2321), .B2(n2145), .ZN(n2148)
         );
  NAND2_X1 U2631 ( .A1(n2192), .A2(n4288), .ZN(n2147) );
  NAND2_X1 U2634 ( .A1(n2189), .A2(n4233), .ZN(n2166) );
  OAI22_X1 U2635 ( .A1(n2157), .A2(n2156), .B1(n2155), .B2(n2154), .ZN(n2164)
         );
  OAI22_X1 U2636 ( .A1(n2161), .A2(n2160), .B1(n2159), .B2(n2158), .ZN(n2163)
         );
  OAI21_X1 U2637 ( .B1(n2164), .B2(n2163), .A(n2162), .ZN(n2165) );
  AOI22_X1 U2638 ( .A1(n2174), .A2(n3387), .B1(n2172), .B2(n2171), .ZN(n2278)
         );
  AND2_X1 U2639 ( .A1(n2174), .A2(n2173), .ZN(n2182) );
  NAND2_X1 U2640 ( .A1(n2296), .A2(n2175), .ZN(n2181) );
  INV_X1 U2641 ( .A(n2176), .ZN(n2177) );
  OR2_X1 U2642 ( .A1(n2280), .A2(n2177), .ZN(n2179) );
  MUX2_X1 U2643 ( .A(n2179), .B(n2219), .S(n2178), .Z(n2180) );
  OAI211_X1 U2644 ( .C1(n2278), .C2(n2182), .A(n2181), .B(n2180), .ZN(n2183)
         );
  AOI21_X1 U2645 ( .B1(n2299), .B2(n2184), .A(n2183), .ZN(n2187) );
  NAND2_X1 U2646 ( .A1(n2185), .A2(n2290), .ZN(n2186) );
  OAI211_X1 U2647 ( .C1(n2188), .C2(n2288), .A(n2187), .B(n2186), .ZN(n2415)
         );
  NAND2_X1 U2648 ( .A1(n2189), .A2(n4287), .ZN(n2213) );
  AOI22_X1 U2649 ( .A1(n2321), .A2(n2191), .B1(n2323), .B2(n2190), .ZN(n2204)
         );
  NAND2_X1 U2650 ( .A1(n2192), .A2(n2329), .ZN(n2203) );
  OR2_X1 U2651 ( .A1(n2199), .A2(n2193), .ZN(n2317) );
  INV_X1 U2652 ( .A(n2242), .ZN(n2195) );
  OAI22_X1 U2653 ( .A1(n2196), .A2(n2314), .B1(n2317), .B2(n2195), .ZN(n2197)
         );
  INV_X1 U2654 ( .A(n2197), .ZN(n2202) );
  OR2_X1 U2655 ( .A1(n2199), .A2(n2198), .ZN(n2313) );
  INV_X1 U2656 ( .A(n2313), .ZN(n2243) );
  MUX2_X1 U2657 ( .A(n2256), .B(n4298), .S(n2262), .Z(n2200) );
  NAND2_X1 U2658 ( .A1(n2243), .A2(n2200), .ZN(n2201) );
  AND4_X1 U2659 ( .A1(n2204), .A2(n2203), .A3(n2202), .A4(n2201), .ZN(n2212)
         );
  OAI22_X1 U2660 ( .A1(n2305), .A2(n2205), .B1(n106), .B2(n2294), .ZN(n2208)
         );
  OAI21_X1 U2661 ( .B1(n2207), .B2(n2206), .A(n4278), .ZN(n2307) );
  AOI21_X1 U2662 ( .B1(n2309), .B2(n2208), .A(n2307), .ZN(n2211) );
  OR2_X1 U2663 ( .A1(n2209), .A2(n2254), .ZN(n2210) );
  NAND4_X1 U2664 ( .A1(n2213), .A2(n2212), .A3(n2211), .A4(n2210), .ZN(n2396)
         );
  OAI22_X1 U2665 ( .A1(n2217), .A2(n2216), .B1(n2215), .B2(n2214), .ZN(n2225)
         );
  OAI22_X1 U2666 ( .A1(n2219), .A2(n2230), .B1(n3363), .B2(n2218), .ZN(n2295)
         );
  AOI21_X1 U2667 ( .B1(n2296), .B2(n2220), .A(n2295), .ZN(n2223) );
  NAND2_X1 U2668 ( .A1(n2299), .A2(n2221), .ZN(n2222) );
  NAND2_X1 U2669 ( .A1(n2223), .A2(n2222), .ZN(n2224) );
  AOI21_X1 U2670 ( .B1(n2230), .B2(n2225), .A(n2224), .ZN(n2226) );
  OAI21_X1 U2671 ( .B1(n2227), .B2(n2288), .A(n2226), .ZN(n2417) );
  INV_X1 U2672 ( .A(n2228), .ZN(n2276) );
  AND2_X1 U2673 ( .A1(n2309), .A2(n2276), .ZN(n2232) );
  OAI22_X1 U2674 ( .A1(n2232), .A2(n2231), .B1(n1635), .B2(n2229), .ZN(n2252)
         );
  AOI22_X1 U2675 ( .A1(n2329), .A2(n2234), .B1(n2233), .B2(n4287), .ZN(n2251)
         );
  NAND2_X1 U2676 ( .A1(n2323), .A2(n2235), .ZN(n2237) );
  OAI211_X1 U2677 ( .C1(n2317), .C2(n2238), .A(n2237), .B(n2236), .ZN(n2247)
         );
  NAND2_X1 U2678 ( .A1(n2321), .A2(n2239), .ZN(n2245) );
  INV_X1 U2679 ( .A(n2314), .ZN(n2241) );
  AOI22_X1 U2680 ( .A1(n2243), .A2(n2242), .B1(n2241), .B2(n2240), .ZN(n2244)
         );
  NAND2_X1 U2681 ( .A1(n2245), .A2(n2244), .ZN(n2246) );
  NOR2_X1 U2682 ( .A1(n2247), .A2(n2246), .ZN(n2250) );
  NAND2_X1 U2683 ( .A1(n2248), .A2(n4233), .ZN(n2249) );
  NAND4_X1 U2684 ( .A1(n2252), .A2(n2251), .A3(n2250), .A4(n2249), .ZN(n2394)
         );
  INV_X1 U2685 ( .A(n2307), .ZN(n2253) );
  OAI21_X1 U2686 ( .B1(n2255), .B2(n2254), .A(n2253), .ZN(n2274) );
  INV_X1 U2687 ( .A(n2256), .ZN(n2259) );
  MUX2_X1 U2688 ( .A(n2259), .B(n2258), .S(n2257), .Z(n2260) );
  INV_X1 U2689 ( .A(n4298), .ZN(n2264) );
  MUX2_X1 U2690 ( .A(n2264), .B(n2263), .S(n2262), .Z(n2312) );
  OAI22_X1 U2691 ( .A1(n2265), .A2(n2314), .B1(n2317), .B2(n2312), .ZN(n2266)
         );
  AOI22_X1 U2692 ( .A1(n2321), .A2(n2269), .B1(n2323), .B2(n2268), .ZN(n2273)
         );
  OAI22_X1 U2693 ( .A1(n2305), .A2(n164), .B1(n106), .B2(n2270), .ZN(n2271) );
  NAND2_X1 U2694 ( .A1(n2309), .A2(n2271), .ZN(n2272) );
  NAND2_X1 U2695 ( .A1(n2296), .A2(n2276), .ZN(n2283) );
  AOI21_X1 U2698 ( .B1(n2299), .B2(n1820), .A(n2284), .ZN(n2287) );
  NAND2_X1 U2699 ( .A1(n2285), .A2(n2290), .ZN(n2286) );
  NAND2_X1 U2700 ( .A1(n2291), .A2(n1635), .ZN(n2303) );
  NAND2_X1 U2701 ( .A1(n2293), .A2(n2292), .ZN(n2302) );
  INV_X1 U2702 ( .A(n2294), .ZN(n2297) );
  AOI21_X1 U2703 ( .B1(n2297), .B2(n2296), .A(n2295), .ZN(n2301) );
  NAND2_X1 U2704 ( .A1(n2299), .A2(n2298), .ZN(n2300) );
  NAND4_X1 U2705 ( .A1(n2303), .A2(n2302), .A3(n2301), .A4(n2300), .ZN(n2416)
         );
  OAI22_X1 U2706 ( .A1(n2306), .A2(n2305), .B1(n2304), .B2(n106), .ZN(n2308)
         );
  AOI21_X1 U2707 ( .B1(n2309), .B2(n2308), .A(n2307), .ZN(n2332) );
  NAND2_X1 U2708 ( .A1(n2311), .A2(n4233), .ZN(n2327) );
  OAI22_X1 U2709 ( .A1(n2315), .A2(n2314), .B1(n2313), .B2(n2312), .ZN(n2319)
         );
  NOR2_X1 U2710 ( .A1(n2317), .A2(n2316), .ZN(n2318) );
  NOR2_X1 U2711 ( .A1(n2319), .A2(n2318), .ZN(n2326) );
  NAND2_X1 U2712 ( .A1(n2321), .A2(n2320), .ZN(n2325) );
  NAND2_X1 U2713 ( .A1(n2323), .A2(n2322), .ZN(n2324) );
  NAND4_X1 U2714 ( .A1(n2327), .A2(n2326), .A3(n2325), .A4(n2324), .ZN(n2328)
         );
  AOI21_X1 U2715 ( .B1(n2330), .B2(n2329), .A(n2328), .ZN(n2331) );
  OAI211_X1 U2716 ( .C1(n4312), .C2(n2333), .A(n2332), .B(n2331), .ZN(n2395)
         );
  MUX2_X1 U2717 ( .A(n2420), .B(n2391), .S(n91), .Z(n3711) );
  INV_X1 U2718 ( .A(n3711), .ZN(n3965) );
  INV_X1 U2719 ( .A(bmask_a_i[0]), .ZN(n2335) );
  INV_X1 U2720 ( .A(n2725), .ZN(n2386) );
  INV_X1 U2721 ( .A(bmask_a_i[1]), .ZN(n2336) );
  OR2_X1 U2722 ( .A1(n2336), .A2(bmask_a_i[0]), .ZN(n2727) );
  INV_X1 U2723 ( .A(n2727), .ZN(n2367) );
  NAND2_X1 U2724 ( .A1(n4189), .A2(n2368), .ZN(n2337) );
  AOI21_X1 U2725 ( .B1(n3875), .B2(n2367), .A(n2338), .ZN(n2340) );
  MUX2_X1 U2726 ( .A(n2393), .B(n2418), .S(n2376), .Z(n3853) );
  NAND2_X1 U2727 ( .A1(n3853), .A2(n2372), .ZN(n2339) );
  MUX2_X1 U2728 ( .A(n2393), .B(n2418), .S(n91), .Z(n3852) );
  NAND2_X1 U2729 ( .A1(n3852), .A2(n2368), .ZN(n2343) );
  OAI211_X1 U2730 ( .C1(n4193), .C2(n2727), .A(n2344), .B(n2343), .ZN(n2383)
         );
  NOR2_X1 U2732 ( .A1(n2345), .A2(bmask_a_i[2]), .ZN(n2362) );
  NAND2_X1 U2733 ( .A1(n2362), .A2(n2369), .ZN(n2346) );
  NOR2_X1 U2735 ( .A1(n2348), .A2(bmask_a_i[3]), .ZN(n2370) );
  NAND2_X1 U2736 ( .A1(n2370), .A2(bmask_a_i[4]), .ZN(n2349) );
  NAND2_X1 U2737 ( .A1(n3595), .A2(n2367), .ZN(n2350) );
  INV_X1 U2738 ( .A(n3380), .ZN(n2649) );
  NAND2_X1 U2739 ( .A1(n2352), .A2(bmask_a_i[4]), .ZN(n2353) );
  MUX2_X1 U2740 ( .A(n4224), .B(n2403), .S(n2376), .Z(n3145) );
  NAND2_X1 U2741 ( .A1(n3145), .A2(n2367), .ZN(n2355) );
  NAND2_X1 U2742 ( .A1(n2967), .A2(n2725), .ZN(n2354) );
  NAND2_X1 U2743 ( .A1(n3788), .A2(n2367), .ZN(n2360) );
  NAND2_X1 U2745 ( .A1(n4015), .A2(n2725), .ZN(n2366) );
  MUX2_X1 U2746 ( .A(n2417), .B(n2394), .S(n2376), .Z(n3821) );
  NAND2_X1 U2747 ( .A1(n3821), .A2(n2372), .ZN(n2365) );
  NAND2_X1 U2748 ( .A1(n2362), .A2(bmask_a_i[4]), .ZN(n2363) );
  AOI21_X1 U2749 ( .B1(n3999), .B2(n2368), .A(n2363), .ZN(n2364) );
  AND3_X1 U2750 ( .A1(n2366), .A2(n2365), .A3(n2364), .ZN(n2380) );
  NAND2_X1 U2752 ( .A1(n3794), .A2(n2367), .ZN(n2379) );
  MUX2_X1 U2753 ( .A(n2415), .B(n2396), .S(n91), .Z(n4013) );
  NAND2_X1 U2754 ( .A1(n4013), .A2(n2367), .ZN(n2375) );
  MUX2_X1 U2755 ( .A(n2417), .B(n2394), .S(n91), .Z(n3820) );
  NAND2_X1 U2756 ( .A1(n3820), .A2(n2368), .ZN(n2374) );
  NAND2_X1 U2757 ( .A1(n2370), .A2(n2369), .ZN(n2371) );
  AOI21_X1 U2758 ( .B1(n4060), .B2(n2372), .A(n2371), .ZN(n2373) );
  AND3_X1 U2759 ( .A1(n2374), .A2(n2375), .A3(n2373), .ZN(n2378) );
  MUX2_X1 U2760 ( .A(n2395), .B(n2416), .S(n2376), .Z(n2846) );
  NAND2_X1 U2761 ( .A1(n2846), .A2(n2725), .ZN(n2377) );
  AOI22_X1 U2762 ( .A1(n2380), .A2(n2379), .B1(n2378), .B2(n2377), .ZN(n2381)
         );
  INV_X1 U2763 ( .A(operand_c_i[8]), .ZN(n2705) );
  NAND2_X1 U2764 ( .A1(n2385), .A2(n1014), .ZN(n2739) );
  OR2_X1 U2765 ( .A1(n2726), .A2(n2727), .ZN(n4184) );
  INV_X1 U2766 ( .A(n4184), .ZN(n3750) );
  AOI22_X1 U2767 ( .A1(n3750), .A2(n4015), .B1(n3595), .B2(n4059), .ZN(n2732)
         );
  OAI21_X1 U2768 ( .B1(n2408), .B2(n2388), .A(n2387), .ZN(n2422) );
  INV_X1 U2769 ( .A(n2422), .ZN(n2624) );
  NOR4_X1 U2770 ( .A1(n4225), .A2(n149), .A3(operand_a_i[9]), .A4(n167), .ZN(
        n2426) );
  NOR4_X1 U2771 ( .A1(operand_a_i[23]), .A2(operand_a_i[25]), .A3(
        operand_a_i[24]), .A4(operand_a_i[26]), .ZN(n2425) );
  NOR4_X1 U2772 ( .A1(operand_a_i[22]), .A2(operand_a_i[21]), .A3(
        operand_a_i[20]), .A4(operand_a_i[19]), .ZN(n2424) );
  NOR4_X1 U2773 ( .A1(n72), .A2(operand_a_i[17]), .A3(operand_a_i[15]), .A4(
        operand_a_i[16]), .ZN(n2423) );
  NAND4_X1 U2774 ( .A1(n2426), .A2(n2425), .A3(n2424), .A4(n2423), .ZN(n2427)
         );
  NOR3_X1 U2775 ( .A1(operand_a_i[28]), .A2(operand_a_i[11]), .A3(n2427), .ZN(
        n2431) );
  NOR2_X1 U2776 ( .A1(operand_a_i[27]), .A2(n4300), .ZN(n2430) );
  NOR2_X1 U2777 ( .A1(n163), .A2(operand_a_i[13]), .ZN(n2429) );
  NOR2_X1 U2778 ( .A1(n54), .A2(operand_a_i[30]), .ZN(n2428) );
  NAND4_X1 U2779 ( .A1(n2431), .A2(n2430), .A3(n2429), .A4(n2428), .ZN(n2461)
         );
  OAI22_X1 U2780 ( .A1(operand_b_i[19]), .A2(operand_a_i[19]), .B1(n4194), 
        .B2(n72), .ZN(n2435) );
  OAI22_X1 U2781 ( .A1(operand_a_i[5]), .A2(operand_b_i[5]), .B1(
        operand_a_i[13]), .B2(operand_b_i[13]), .ZN(n2434) );
  OAI22_X1 U2782 ( .A1(operand_b_i[2]), .A2(operand_a_i[2]), .B1(n4328), .B2(
        operand_a_i[17]), .ZN(n2433) );
  OAI22_X1 U2783 ( .A1(operand_a_i[30]), .A2(operand_b_i[30]), .B1(
        operand_a_i[20]), .B2(operand_b_i[20]), .ZN(n2432) );
  NOR4_X1 U2784 ( .A1(n2435), .A2(n2434), .A3(n2433), .A4(n2432), .ZN(n2459)
         );
  NOR2_X1 U2785 ( .A1(n163), .A2(operand_b_i[12]), .ZN(n2439) );
  NOR2_X1 U2786 ( .A1(operand_a_i[7]), .A2(operand_b_i[7]), .ZN(n2438) );
  OAI22_X1 U2787 ( .A1(n54), .A2(operand_b_i[29]), .B1(operand_a_i[23]), .B2(
        operand_b_i[23]), .ZN(n2437) );
  OAI22_X1 U2788 ( .A1(operand_b_i[4]), .A2(operand_a_i[4]), .B1(n4300), .B2(
        operand_b_i[14]), .ZN(n2436) );
  NOR4_X1 U2789 ( .A1(n2439), .A2(n2438), .A3(n2437), .A4(n2436), .ZN(n2458)
         );
  OAI22_X1 U2790 ( .A1(operand_b_i[3]), .A2(n48), .B1(operand_a_i[6]), .B2(
        operand_b_i[6]), .ZN(n2453) );
  NOR2_X1 U2791 ( .A1(operand_b_i[16]), .A2(operand_a_i[16]), .ZN(n2442) );
  NOR2_X1 U2792 ( .A1(n168), .A2(operand_b_i[10]), .ZN(n2441) );
  NOR2_X1 U2793 ( .A1(n110), .A2(operand_a_i[25]), .ZN(n2440) );
  NOR3_X1 U2794 ( .A1(n2442), .A2(n2441), .A3(n2440), .ZN(n2450) );
  NOR2_X1 U2795 ( .A1(operand_a_i[28]), .A2(operand_b_i[28]), .ZN(n2444) );
  NOR2_X1 U2796 ( .A1(n4304), .A2(operand_b_i[31]), .ZN(n2443) );
  NOR2_X1 U2797 ( .A1(n2444), .A2(n2443), .ZN(n2448) );
  NOR2_X1 U2798 ( .A1(n170), .A2(operand_a_i[26]), .ZN(n2446) );
  NOR2_X1 U2799 ( .A1(operand_a_i[21]), .A2(operand_b_i[21]), .ZN(n2445) );
  NOR2_X1 U2800 ( .A1(n2446), .A2(n2445), .ZN(n2447) );
  AND2_X1 U2801 ( .A1(n2448), .A2(n2447), .ZN(n2449) );
  OAI211_X1 U2802 ( .C1(operand_a_i[24]), .C2(n4340), .A(n2450), .B(n2449), 
        .ZN(n2452) );
  OAI22_X1 U2803 ( .A1(operand_a_i[22]), .A2(operand_b_i[22]), .B1(
        operand_a_i[27]), .B2(n64), .ZN(n2451) );
  OR3_X1 U2804 ( .A1(n2453), .A2(n2452), .A3(n2451), .ZN(n2456) );
  OAI22_X1 U2805 ( .A1(n149), .A2(n4196), .B1(operand_a_i[11]), .B2(n150), 
        .ZN(n2455) );
  OAI22_X1 U2806 ( .A1(operand_a_i[9]), .A2(n4195), .B1(operand_a_i[15]), .B2(
        operand_b_i[15]), .ZN(n2454) );
  NOR3_X1 U2807 ( .A1(n2456), .A2(n2455), .A3(n2454), .ZN(n2457) );
  NAND3_X1 U2808 ( .A1(n2459), .A2(n2458), .A3(n2457), .ZN(n2460) );
  MUX2_X1 U2809 ( .A(n2461), .B(n2460), .S(n3683), .Z(n2494) );
  NOR4_X1 U2810 ( .A1(operand_a_i[2]), .A2(n48), .A3(operand_a_i[4]), .A4(
        operand_a_i[5]), .ZN(n2462) );
  NAND4_X1 U2811 ( .A1(n4127), .A2(n2543), .A3(n4071), .A4(n2462), .ZN(n2466)
         );
  OR2_X1 U2812 ( .A1(n2463), .A2(operand_b_i[0]), .ZN(n2545) );
  OAI21_X1 U2813 ( .B1(operand_a_i[0]), .B2(n2661), .A(n2545), .ZN(n4145) );
  XNOR2_X1 U2814 ( .A(n2464), .B(operand_a_i[1]), .ZN(n3689) );
  NAND2_X1 U2815 ( .A1(n4145), .A2(n3689), .ZN(n2465) );
  MUX2_X1 U2816 ( .A(n2466), .B(n2465), .S(n3683), .Z(n2467) );
  INV_X1 U2817 ( .A(n2467), .ZN(n2492) );
  AOI22_X1 U2818 ( .A1(operand_a_i[20]), .A2(operand_b_i[20]), .B1(
        operand_a_i[13]), .B2(operand_b_i[13]), .ZN(n2471) );
  AOI22_X1 U2819 ( .A1(operand_b_i[3]), .A2(n48), .B1(operand_a_i[23]), .B2(
        operand_b_i[23]), .ZN(n2470) );
  AOI22_X1 U2820 ( .A1(operand_b_i[4]), .A2(operand_a_i[4]), .B1(n4194), .B2(
        n72), .ZN(n2469) );
  AOI22_X1 U2821 ( .A1(operand_b_i[19]), .A2(operand_a_i[19]), .B1(
        operand_a_i[22]), .B2(operand_b_i[22]), .ZN(n2468) );
  NAND4_X1 U2822 ( .A1(n2471), .A2(n2470), .A3(n2469), .A4(n2468), .ZN(n2490)
         );
  AOI22_X1 U2823 ( .A1(operand_a_i[9]), .A2(n4195), .B1(operand_a_i[2]), .B2(
        operand_b_i[2]), .ZN(n2483) );
  AOI22_X1 U2824 ( .A1(operand_a_i[5]), .A2(operand_b_i[5]), .B1(
        operand_a_i[6]), .B2(operand_b_i[6]), .ZN(n2475) );
  AOI22_X1 U2825 ( .A1(n4328), .A2(operand_a_i[17]), .B1(operand_a_i[30]), 
        .B2(operand_b_i[30]), .ZN(n2474) );
  NAND2_X1 U2826 ( .A1(operand_a_i[21]), .A2(operand_b_i[21]), .ZN(n2473) );
  NAND2_X1 U2827 ( .A1(operand_a_i[7]), .A2(operand_b_i[7]), .ZN(n2472) );
  NAND4_X1 U2828 ( .A1(n2475), .A2(n2474), .A3(n2473), .A4(n2472), .ZN(n2481)
         );
  NAND2_X1 U2829 ( .A1(n163), .A2(operand_b_i[12]), .ZN(n2479) );
  NAND2_X1 U2830 ( .A1(operand_a_i[28]), .A2(operand_b_i[28]), .ZN(n2478) );
  NAND2_X1 U2831 ( .A1(n168), .A2(operand_b_i[10]), .ZN(n2477) );
  NAND2_X1 U2832 ( .A1(n110), .A2(operand_a_i[25]), .ZN(n2476) );
  NAND4_X1 U2833 ( .A1(n2479), .A2(n2478), .A3(n2477), .A4(n2476), .ZN(n2480)
         );
  AOI211_X1 U2834 ( .C1(operand_a_i[27]), .C2(n64), .A(n2481), .B(n2480), .ZN(
        n2482) );
  NAND2_X1 U2835 ( .A1(operand_a_i[31]), .A2(operand_b_i[31]), .ZN(n3949) );
  NAND3_X1 U2836 ( .A1(n2483), .A2(n2482), .A3(n148), .ZN(n2489) );
  AOI22_X1 U2837 ( .A1(n4340), .A2(operand_a_i[24]), .B1(n4300), .B2(
        operand_b_i[14]), .ZN(n2487) );
  AOI22_X1 U2838 ( .A1(operand_a_i[26]), .A2(n170), .B1(n54), .B2(
        operand_b_i[29]), .ZN(n2486) );
  AOI22_X1 U2839 ( .A1(operand_b_i[16]), .A2(operand_a_i[16]), .B1(
        operand_a_i[11]), .B2(n150), .ZN(n2485) );
  AOI22_X1 U2840 ( .A1(n149), .A2(n4196), .B1(operand_a_i[15]), .B2(
        operand_b_i[15]), .ZN(n2484) );
  NAND4_X1 U2841 ( .A1(n2487), .A2(n2486), .A3(n2485), .A4(n2484), .ZN(n2488)
         );
  NOR3_X1 U2842 ( .A1(n2490), .A2(n2489), .A3(n2488), .ZN(n2491) );
  NAND2_X1 U2843 ( .A1(n2492), .A2(n2491), .ZN(n2493) );
  OR2_X1 U2844 ( .A1(n2494), .A2(n2493), .ZN(n2626) );
  INV_X1 U2845 ( .A(n2497), .ZN(n2498) );
  NAND2_X1 U2846 ( .A1(n2498), .A2(n4131), .ZN(n2499) );
  OR2_X1 U2847 ( .A1(n2662), .A2(n2500), .ZN(n2667) );
  INV_X1 U2848 ( .A(n4038), .ZN(n4146) );
  OR2_X1 U2849 ( .A1(n2667), .A2(n52), .ZN(n2944) );
  INV_X1 U2850 ( .A(n2944), .ZN(n2501) );
  NAND2_X1 U2851 ( .A1(n2501), .A2(n4337), .ZN(n3443) );
  INV_X1 U2852 ( .A(n3443), .ZN(n2892) );
  INV_X1 U2853 ( .A(operand_b_i[23]), .ZN(n2945) );
  OR2_X1 U2854 ( .A1(n2945), .A2(operand_a_i[23]), .ZN(n2517) );
  BUF_X1 U2855 ( .A(n2517), .Z(n2504) );
  NAND2_X1 U2856 ( .A1(operand_a_i[23]), .A2(n2505), .ZN(n2518) );
  OAI21_X1 U2857 ( .B1(n2621), .B2(n2507), .A(n2506), .ZN(n2520) );
  NOR2_X1 U2858 ( .A1(n2508), .A2(operand_a_i[17]), .ZN(n2587) );
  NAND2_X1 U2859 ( .A1(n3765), .A2(operand_a_i[16]), .ZN(n2510) );
  NAND2_X1 U2860 ( .A1(n2508), .A2(operand_a_i[17]), .ZN(n2589) );
  INV_X1 U2861 ( .A(operand_b_i[18]), .ZN(n3163) );
  NAND2_X1 U2862 ( .A1(n3163), .A2(operand_a_i[18]), .ZN(n2509) );
  OAI211_X1 U2863 ( .C1(n2587), .C2(n2510), .A(n2589), .B(n2509), .ZN(n2512)
         );
  AOI22_X1 U2864 ( .A1(operand_b_i[19]), .A2(n4105), .B1(n71), .B2(
        operand_b_i[18]), .ZN(n2511) );
  INV_X1 U2865 ( .A(operand_b_i[19]), .ZN(n3025) );
  INV_X1 U2866 ( .A(operand_b_i[20]), .ZN(n3918) );
  AOI22_X1 U2867 ( .A1(operand_a_i[19]), .A2(n3025), .B1(n3918), .B2(
        operand_a_i[20]), .ZN(n2513) );
  AOI22_X1 U2868 ( .A1(operand_b_i[20]), .A2(n4067), .B1(n4075), .B2(
        operand_b_i[21]), .ZN(n2516) );
  OR2_X1 U2869 ( .A1(n2514), .A2(operand_b_i[22]), .ZN(n3120) );
  OAI21_X1 U2870 ( .B1(operand_b_i[21]), .B2(n4075), .A(n3120), .ZN(n2515) );
  AND2_X1 U2871 ( .A1(n2517), .A2(n2518), .ZN(n2918) );
  INV_X1 U2872 ( .A(operand_b_i[22]), .ZN(n3130) );
  OR2_X1 U2873 ( .A1(n3130), .A2(operand_a_i[22]), .ZN(n3119) );
  INV_X1 U2874 ( .A(operand_b_i[27]), .ZN(n2848) );
  OR2_X1 U2875 ( .A1(n2848), .A2(operand_a_i[27]), .ZN(n2532) );
  AND2_X1 U2876 ( .A1(n2528), .A2(n2532), .ZN(n2852) );
  INV_X1 U2877 ( .A(n2531), .ZN(n2523) );
  INV_X1 U2878 ( .A(operand_b_i[28]), .ZN(n3854) );
  OR2_X1 U2879 ( .A1(n3854), .A2(operand_a_i[28]), .ZN(n2534) );
  AND2_X1 U2880 ( .A1(n2523), .A2(n2534), .ZN(n3860) );
  NAND2_X1 U2881 ( .A1(n3949), .A2(n2524), .ZN(n3950) );
  XNOR2_X1 U2882 ( .A(operand_a_i[24]), .B(operand_b_i[24]), .ZN(n3533) );
  XNOR2_X1 U2883 ( .A(operand_a_i[26]), .B(operand_b_i[26]), .ZN(n3190) );
  XNOR2_X1 U2884 ( .A(operand_a_i[25]), .B(operand_b_i[25]), .ZN(n4037) );
  XNOR2_X1 U2885 ( .A(operand_a_i[29]), .B(operand_b_i[29]), .ZN(n2821) );
  XNOR2_X1 U2886 ( .A(operand_a_i[30]), .B(operand_b_i[30]), .ZN(n3295) );
  INV_X1 U2887 ( .A(n2565), .ZN(n2584) );
  NAND2_X1 U2888 ( .A1(n4115), .A2(operand_b_i[31]), .ZN(n2542) );
  OR2_X1 U2889 ( .A1(n4115), .A2(operand_b_i[31]), .ZN(n2536) );
  NAND2_X1 U2890 ( .A1(n4112), .A2(operand_b_i[30]), .ZN(n2525) );
  NAND2_X1 U2891 ( .A1(n3950), .A2(n2525), .ZN(n2526) );
  OAI21_X1 U2892 ( .B1(n4302), .B2(n2536), .A(n2526), .ZN(n2541) );
  INV_X1 U2893 ( .A(operand_b_i[24]), .ZN(n3530) );
  INV_X1 U2894 ( .A(operand_b_i[25]), .ZN(n4020) );
  AOI22_X1 U2895 ( .A1(operand_a_i[24]), .A2(n3530), .B1(n4020), .B2(
        operand_a_i[25]), .ZN(n2530) );
  OAI22_X1 U2896 ( .A1(operand_a_i[25]), .A2(n4020), .B1(n3186), .B2(
        operand_a_i[26]), .ZN(n2529) );
  NAND2_X1 U2897 ( .A1(n3186), .A2(operand_a_i[26]), .ZN(n2527) );
  OAI211_X1 U2898 ( .C1(n2530), .C2(n2529), .A(n2528), .B(n2527), .ZN(n2533)
         );
  AOI21_X1 U2899 ( .B1(n2533), .B2(n2532), .A(n2531), .ZN(n2539) );
  INV_X1 U2900 ( .A(operand_b_i[29]), .ZN(n2775) );
  OAI21_X1 U2901 ( .B1(operand_a_i[29]), .B2(n2775), .A(n2534), .ZN(n2538) );
  INV_X1 U2902 ( .A(operand_b_i[30]), .ZN(n2535) );
  AOI22_X1 U2903 ( .A1(operand_a_i[29]), .A2(n2775), .B1(n2535), .B2(
        operand_a_i[30]), .ZN(n2537) );
  INV_X1 U2904 ( .A(n2554), .ZN(n2544) );
  OR2_X1 U2905 ( .A1(n588), .A2(operand_a_i[7]), .ZN(n2558) );
  NAND2_X1 U2906 ( .A1(n2554), .A2(n2558), .ZN(n3976) );
  NOR2_X1 U2907 ( .A1(n3663), .A2(operand_a_i[6]), .ZN(n3652) );
  AOI21_X1 U2908 ( .B1(n2621), .B2(n2544), .A(n2602), .ZN(n2560) );
  AOI22_X1 U2909 ( .A1(operand_b_i[1]), .A2(n2546), .B1(n2547), .B2(
        operand_b_i[2]), .ZN(n2550) );
  OAI21_X1 U2910 ( .B1(operand_b_i[1]), .B2(n2546), .A(n2545), .ZN(n2549) );
  INV_X1 U2911 ( .A(operand_a_i[3]), .ZN(n3011) );
  OAI22_X1 U2912 ( .A1(operand_b_i[3]), .A2(n3011), .B1(n2547), .B2(
        operand_b_i[2]), .ZN(n2548) );
  AOI21_X1 U2913 ( .B1(n2550), .B2(n2549), .A(n2548), .ZN(n2552) );
  OAI22_X1 U2914 ( .A1(operand_a_i[4]), .A2(n3812), .B1(n3479), .B2(
        operand_a_i[3]), .ZN(n2551) );
  OAI22_X1 U2915 ( .A1(n2552), .A2(n2551), .B1(operand_b_i[4]), .B2(n4108), 
        .ZN(n2557) );
  NAND2_X1 U2916 ( .A1(n4079), .A2(operand_b_i[5]), .ZN(n2556) );
  OR2_X1 U2917 ( .A1(n2553), .A2(operand_b_i[6]), .ZN(n2599) );
  OAI211_X1 U2918 ( .C1(operand_b_i[5]), .C2(n4079), .A(n2554), .B(n2599), 
        .ZN(n2555) );
  AOI21_X1 U2919 ( .B1(n2557), .B2(n2556), .A(n2555), .ZN(n2559) );
  OAI22_X1 U2920 ( .A1(n2559), .A2(n2560), .B1(n158), .B2(n2558), .ZN(n3355)
         );
  OR2_X1 U2921 ( .A1(n162), .A2(operand_b_i[12]), .ZN(n2575) );
  OR2_X1 U2922 ( .A1(n3240), .A2(operand_a_i[12]), .ZN(n2580) );
  AND2_X1 U2923 ( .A1(n2575), .A2(n2580), .ZN(n3229) );
  OR2_X1 U2924 ( .A1(n3578), .A2(operand_a_i[13]), .ZN(n2579) );
  AND2_X1 U2925 ( .A1(n2581), .A2(n2579), .ZN(n3564) );
  INV_X1 U2926 ( .A(operand_b_i[11]), .ZN(n2562) );
  OR2_X1 U2927 ( .A1(n2562), .A2(operand_a_i[11]), .ZN(n2573) );
  NAND2_X1 U2928 ( .A1(operand_a_i[11]), .A2(n2562), .ZN(n2576) );
  AND2_X1 U2929 ( .A1(n2573), .A2(n2576), .ZN(n3607) );
  XNOR2_X1 U2930 ( .A(n167), .B(operand_b_i[10]), .ZN(n3324) );
  NAND4_X1 U2931 ( .A1(n3229), .A2(n3564), .A3(n3607), .A4(n3324), .ZN(n2564)
         );
  XNOR2_X1 U2932 ( .A(operand_a_i[15]), .B(operand_b_i[15]), .ZN(n3042) );
  OR2_X1 U2933 ( .A1(n3092), .A2(operand_a_i[14]), .ZN(n3078) );
  AND2_X1 U2934 ( .A1(n3042), .A2(n3078), .ZN(n2582) );
  OR2_X1 U2935 ( .A1(n4098), .A2(operand_b_i[14]), .ZN(n3079) );
  XNOR2_X1 U2936 ( .A(operand_a_i[9]), .B(n4195), .ZN(n3499) );
  XNOR2_X1 U2937 ( .A(operand_a_i[8]), .B(operand_b_i[8]), .ZN(n2563) );
  NOR2_X1 U2938 ( .A1(n4095), .A2(operand_b_i[15]), .ZN(n2583) );
  OAI211_X1 U2939 ( .C1(n2567), .C2(operand_a_i[9]), .A(operand_a_i[8]), .B(
        n2566), .ZN(n2569) );
  NAND2_X1 U2940 ( .A1(n2567), .A2(operand_a_i[9]), .ZN(n2568) );
  OAI211_X1 U2941 ( .C1(operand_b_i[10]), .C2(n2570), .A(n2569), .B(n2568), 
        .ZN(n2574) );
  OR2_X1 U2942 ( .A1(n2571), .A2(n168), .ZN(n2572) );
  NAND3_X1 U2943 ( .A1(n4095), .A2(vector_mode_i[1]), .A3(operand_b_i[15]), 
        .ZN(n2620) );
  AOI21_X1 U2945 ( .B1(n2639), .B2(n3355), .A(n2586), .ZN(n2616) );
  INV_X1 U2946 ( .A(n2587), .ZN(n2588) );
  XNOR2_X1 U2947 ( .A(operand_a_i[16]), .B(operand_b_i[16]), .ZN(n2590) );
  XNOR2_X1 U2948 ( .A(operand_a_i[18]), .B(operand_b_i[18]), .ZN(n3152) );
  NAND3_X1 U2949 ( .A1(n3120), .A2(n2590), .A3(n3152), .ZN(n2592) );
  XNOR2_X1 U2950 ( .A(operand_a_i[19]), .B(operand_b_i[19]), .ZN(n3012) );
  XNOR2_X1 U2951 ( .A(operand_a_i[21]), .B(operand_b_i[21]), .ZN(n3261) );
  NAND2_X1 U2952 ( .A1(n3012), .A2(n3261), .ZN(n2591) );
  NOR2_X1 U2953 ( .A1(n2592), .A2(n2591), .ZN(n2593) );
  XNOR2_X1 U2954 ( .A(operand_a_i[20]), .B(operand_b_i[20]), .ZN(n3902) );
  INV_X1 U2956 ( .A(n2598), .ZN(n2752) );
  INV_X1 U2957 ( .A(n2599), .ZN(n3653) );
  XNOR2_X1 U2958 ( .A(operand_a_i[3]), .B(operand_b_i[3]), .ZN(n3467) );
  XNOR2_X1 U2959 ( .A(operand_a_i[4]), .B(operand_b_i[4]), .ZN(n3798) );
  AND2_X1 U2960 ( .A1(n3467), .A2(n3798), .ZN(n2601) );
  XNOR2_X1 U2961 ( .A(operand_a_i[2]), .B(operand_b_i[2]), .ZN(n3416) );
  XNOR2_X1 U2962 ( .A(operand_a_i[5]), .B(operand_b_i[5]), .ZN(n3727) );
  AND2_X1 U2963 ( .A1(n3416), .A2(n3727), .ZN(n2600) );
  XNOR2_X1 U2964 ( .A(n2770), .B(n154), .ZN(n2743) );
  INV_X1 U2966 ( .A(n2606), .ZN(n2607) );
  XNOR2_X1 U2967 ( .A(n2607), .B(n3683), .ZN(n2610) );
  OR2_X1 U2968 ( .A1(n4163), .A2(n3834), .ZN(n2628) );
  INV_X1 U2969 ( .A(n2628), .ZN(n2609) );
  NAND2_X1 U2970 ( .A1(n2610), .A2(n2609), .ZN(n2769) );
  NAND3_X1 U2972 ( .A1(n66), .A2(n4159), .A3(n2651), .ZN(n2627) );
  INV_X1 U2973 ( .A(n2627), .ZN(n2612) );
  NAND2_X1 U2974 ( .A1(n2612), .A2(n3834), .ZN(n2613) );
  AND2_X1 U2975 ( .A1(n2497), .A2(n2613), .ZN(n2767) );
  NAND2_X1 U2976 ( .A1(n2767), .A2(n2628), .ZN(n2768) );
  OR2_X1 U2977 ( .A1(n2616), .A2(n2668), .ZN(n2617) );
  OAI22_X1 U2978 ( .A1(n2619), .A2(n3363), .B1(n158), .B2(n2620), .ZN(n2622)
         );
  OR2_X1 U2979 ( .A1(n3357), .A2(n2622), .ZN(n2644) );
  MUX2_X1 U2980 ( .A(n2767), .B(n2768), .S(n2644), .Z(n2623) );
  AND2_X1 U2981 ( .A1(n2769), .A2(n2623), .ZN(n2717) );
  NAND2_X1 U2982 ( .A1(n2624), .A2(n4131), .ZN(n2631) );
  NOR2_X1 U2983 ( .A1(n2497), .A2(int_div_div_op_a_signed), .ZN(n2625) );
  AND2_X1 U2984 ( .A1(n2626), .A2(n2625), .ZN(n2630) );
  OAI211_X1 U2985 ( .C1(n169), .C2(is_clpx_i), .A(n2628), .B(n2627), .ZN(n2629) );
  AOI21_X1 U2986 ( .B1(n2631), .B2(n2630), .A(n2629), .ZN(n3437) );
  INV_X1 U2987 ( .A(n2949), .ZN(n2633) );
  OAI21_X1 U2988 ( .B1(n3437), .B2(n2633), .A(n3443), .ZN(n3446) );
  OAI21_X1 U2989 ( .B1(n2892), .B2(n2717), .A(n3446), .ZN(n3596) );
  OAI21_X1 U2990 ( .B1(n149), .B2(n4038), .A(n3596), .ZN(n2634) );
  MUX2_X1 U2991 ( .A(n4017), .B(n2634), .S(n4196), .Z(n2724) );
  OR2_X1 U2992 ( .A1(n3437), .A2(n169), .ZN(n3360) );
  INV_X1 U2993 ( .A(n2717), .ZN(n2635) );
  NOR2_X1 U2994 ( .A1(n3360), .A2(n2635), .ZN(n3628) );
  NAND2_X1 U2995 ( .A1(n3628), .A2(n4315), .ZN(n2722) );
  NAND2_X1 U2996 ( .A1(n2639), .A2(vector_mode_i[1]), .ZN(n3362) );
  AOI22_X1 U2997 ( .A1(n2638), .A2(n3362), .B1(n2641), .B2(n2640), .ZN(n2655)
         );
  INV_X1 U2998 ( .A(n2642), .ZN(n2643) );
  INV_X1 U2999 ( .A(n3361), .ZN(n4162) );
  AOI21_X1 U3000 ( .B1(n2655), .B2(n498), .A(n4162), .ZN(n2645) );
  NAND3_X1 U3001 ( .A1(n2660), .A2(n4160), .A3(n498), .ZN(n2902) );
  INV_X1 U3002 ( .A(n2902), .ZN(n3372) );
  MUX2_X1 U3003 ( .A(n2645), .B(n3372), .S(n2644), .Z(n2659) );
  NOR2_X1 U3004 ( .A1(n2662), .A2(n2646), .ZN(n3373) );
  AND2_X1 U3006 ( .A1(n4160), .A2(n3831), .ZN(n2656) );
  BUF_X1 U3007 ( .A(n2647), .Z(n2652) );
  NAND3_X1 U3008 ( .A1(n2649), .A2(n487), .A3(n2648), .ZN(n2650) );
  OAI21_X1 U3009 ( .B1(n2652), .B2(n2651), .A(n2650), .ZN(n2653) );
  INV_X1 U3010 ( .A(n2653), .ZN(n2654) );
  OAI211_X1 U3011 ( .C1(n2902), .C2(n3834), .A(n2656), .B(n2654), .ZN(n2893)
         );
  MUX2_X1 U3012 ( .A(n3373), .B(n2893), .S(n2655), .Z(n2658) );
  NAND2_X1 U3013 ( .A1(n2656), .A2(n2660), .ZN(n2657) );
  OAI21_X1 U3014 ( .B1(n4162), .B2(n4337), .A(n2657), .ZN(n2903) );
  OAI21_X1 U3015 ( .B1(n2659), .B2(n2658), .A(n2903), .ZN(n3576) );
  INV_X1 U3016 ( .A(n3576), .ZN(n3623) );
  NAND2_X1 U3017 ( .A1(result_div[8]), .A2(n3988), .ZN(n2714) );
  NAND3_X1 U3018 ( .A1(n2660), .A2(n398), .A3(n498), .ZN(n2684) );
  OR2_X1 U3019 ( .A1(n2684), .A2(n4337), .ZN(n2674) );
  NOR2_X1 U3020 ( .A1(n2674), .A2(n4131), .ZN(n2786) );
  OR2_X1 U3021 ( .A1(n2684), .A2(n3834), .ZN(n2794) );
  NOR2_X1 U3022 ( .A1(n2794), .A2(n2661), .ZN(n3389) );
  OAI21_X1 U3023 ( .B1(n2786), .B2(n3389), .A(n2784), .ZN(n2664) );
  OR3_X1 U3024 ( .A1(n2662), .A2(n3834), .A3(n3350), .ZN(n3386) );
  INV_X1 U3025 ( .A(n3386), .ZN(n2671) );
  NAND2_X1 U3026 ( .A1(n390), .A2(imm_vec_ext_i[0]), .ZN(n2666) );
  NAND2_X1 U3027 ( .A1(n3387), .A2(imm_vec_ext_i[1]), .ZN(n2663) );
  OAI21_X1 U3028 ( .B1(vector_mode_i[0]), .B2(n2666), .A(n2663), .ZN(n2672) );
  NAND2_X1 U3029 ( .A1(n2671), .A2(n2672), .ZN(n2787) );
  NAND2_X1 U3030 ( .A1(n2664), .A2(n2787), .ZN(n3384) );
  NOR2_X1 U3031 ( .A1(n2794), .A2(n3363), .ZN(n3382) );
  AND2_X1 U3032 ( .A1(n3382), .A2(n4195), .ZN(n2665) );
  OR2_X1 U3033 ( .A1(n3384), .A2(n2665), .ZN(n2691) );
  INV_X1 U3034 ( .A(n2666), .ZN(n3395) );
  OAI21_X1 U3035 ( .B1(n2784), .B2(n3395), .A(n2671), .ZN(n2910) );
  INV_X1 U3036 ( .A(n2740), .ZN(n3351) );
  NOR2_X1 U3037 ( .A1(n2667), .A2(n3351), .ZN(n3396) );
  INV_X1 U3038 ( .A(n3396), .ZN(n2788) );
  NAND3_X1 U3039 ( .A1(n2910), .A2(n2668), .A3(n2788), .ZN(n2796) );
  NAND2_X1 U3040 ( .A1(vector_mode_i[1]), .A2(n4196), .ZN(n2669) );
  NOR2_X1 U3041 ( .A1(n2794), .A2(n2669), .ZN(n2670) );
  OR2_X1 U3042 ( .A1(n2796), .A2(n2670), .ZN(n2690) );
  AND2_X1 U3043 ( .A1(n2691), .A2(n2690), .ZN(n2697) );
  INV_X1 U3044 ( .A(n2697), .ZN(n2679) );
  NAND2_X1 U3045 ( .A1(n3396), .A2(n3387), .ZN(n3393) );
  INV_X1 U3046 ( .A(n3393), .ZN(n2683) );
  INV_X1 U3047 ( .A(imm_vec_ext_i[0]), .ZN(n3385) );
  AND2_X1 U3048 ( .A1(n2683), .A2(n3385), .ZN(n2782) );
  AOI22_X1 U3049 ( .A1(n3396), .A2(n2672), .B1(n3387), .B2(n2671), .ZN(n2676)
         );
  INV_X1 U3050 ( .A(n3683), .ZN(n4161) );
  NAND2_X1 U3051 ( .A1(n2784), .A2(n4161), .ZN(n2673) );
  OR2_X1 U3052 ( .A1(n2684), .A2(n2673), .ZN(n2777) );
  INV_X1 U3053 ( .A(n2777), .ZN(n2675) );
  INV_X2 U3054 ( .A(n2674), .ZN(n3394) );
  AOI22_X1 U3055 ( .A1(n2675), .A2(n2464), .B1(n3394), .B2(n3363), .ZN(n3398)
         );
  NAND2_X1 U3056 ( .A1(n2676), .A2(n3398), .ZN(n2678) );
  NAND2_X1 U3057 ( .A1(n3382), .A2(n52), .ZN(n3391) );
  NOR2_X1 U3058 ( .A1(n3391), .A2(operand_b_i[10]), .ZN(n2677) );
  OR3_X1 U3059 ( .A1(n2782), .A2(n2678), .A3(n2677), .ZN(n2687) );
  INV_X1 U3060 ( .A(n2687), .ZN(n2701) );
  NOR2_X1 U3061 ( .A1(n2679), .A2(n2701), .ZN(n3606) );
  NOR2_X1 U3062 ( .A1(n3386), .A2(n52), .ZN(n2703) );
  INV_X1 U3063 ( .A(operand_c_i[24]), .ZN(n3534) );
  NAND2_X1 U3064 ( .A1(n2703), .A2(n4304), .ZN(n3219) );
  NAND2_X1 U3065 ( .A1(n3394), .A2(n4340), .ZN(n2680) );
  OAI211_X1 U3066 ( .C1(n3228), .C2(n3534), .A(n3219), .B(n2680), .ZN(n4135)
         );
  INV_X1 U3067 ( .A(n2690), .ZN(n2688) );
  AND2_X1 U3068 ( .A1(n2691), .A2(n2688), .ZN(n2699) );
  INV_X1 U3069 ( .A(n2699), .ZN(n2681) );
  NOR2_X1 U3070 ( .A1(n2681), .A2(n2701), .ZN(n3617) );
  INV_X1 U3071 ( .A(operand_c_i[16]), .ZN(n3768) );
  NAND2_X1 U3072 ( .A1(n2703), .A2(operand_a_i[23]), .ZN(n3221) );
  NAND2_X1 U3073 ( .A1(n3394), .A2(operand_b_i[16]), .ZN(n2682) );
  OAI211_X1 U3074 ( .C1(n3228), .C2(n3768), .A(n3221), .B(n2682), .ZN(n4153)
         );
  AOI22_X1 U3075 ( .A1(n3606), .A2(n4135), .B1(n3617), .B2(n4153), .ZN(n2713)
         );
  MUX2_X1 U3076 ( .A(n4106), .B(n4127), .S(n2683), .Z(n3771) );
  INV_X1 U3077 ( .A(n3771), .ZN(n4140) );
  NAND3_X1 U3078 ( .A1(n2788), .A2(n2684), .A3(n3386), .ZN(n3407) );
  AND2_X1 U3079 ( .A1(n3387), .A2(n52), .ZN(n2685) );
  NAND2_X1 U3080 ( .A1(n3394), .A2(n2685), .ZN(n3979) );
  NAND2_X1 U3081 ( .A1(n3407), .A2(n3979), .ZN(n2686) );
  NOR2_X1 U3082 ( .A1(n2687), .A2(n2686), .ZN(n2700) );
  INV_X1 U3083 ( .A(n2700), .ZN(n2689) );
  OR2_X1 U3084 ( .A1(n2691), .A2(n2688), .ZN(n2702) );
  NOR2_X1 U3085 ( .A1(n2689), .A2(n2702), .ZN(n3601) );
  NOR2_X1 U3086 ( .A1(n2691), .A2(n2690), .ZN(n2698) );
  INV_X1 U3087 ( .A(n2698), .ZN(n2692) );
  NOR2_X1 U3088 ( .A1(n2692), .A2(n2701), .ZN(n3598) );
  INV_X1 U3089 ( .A(operand_c_i[0]), .ZN(n2694) );
  NAND2_X1 U3090 ( .A1(n2703), .A2(operand_a_i[7]), .ZN(n3223) );
  NAND2_X1 U3091 ( .A1(n3394), .A2(operand_b_i[0]), .ZN(n2693) );
  OAI211_X1 U3092 ( .C1(n3228), .C2(n2694), .A(n3223), .B(n2693), .ZN(n4141)
         );
  AOI22_X1 U3093 ( .A1(n4140), .A2(n3601), .B1(n3598), .B2(n4141), .ZN(n2712)
         );
  INV_X1 U3094 ( .A(n3076), .ZN(n3225) );
  NAND2_X1 U3095 ( .A1(n3225), .A2(n3844), .ZN(n2696) );
  OAI21_X1 U3096 ( .B1(n4140), .B2(n3225), .A(n2696), .ZN(n4132) );
  NAND2_X1 U3097 ( .A1(n2700), .A2(n2697), .ZN(n3562) );
  NAND2_X1 U3098 ( .A1(n2700), .A2(n2698), .ZN(n3612) );
  OAI22_X1 U3099 ( .A1(n4132), .A2(n3562), .B1(n3612), .B2(n4127), .ZN(n2710)
         );
  NAND2_X1 U3100 ( .A1(n2700), .A2(n2699), .ZN(n3570) );
  MUX2_X1 U3101 ( .A(operand_a_i[16]), .B(n4198), .S(n3076), .Z(n4143) );
  INV_X1 U3102 ( .A(n4143), .ZN(n2708) );
  NOR2_X1 U3103 ( .A1(n2702), .A2(n2701), .ZN(n3615) );
  NAND2_X1 U3104 ( .A1(n2703), .A2(operand_a_i[15]), .ZN(n3227) );
  NAND2_X1 U3105 ( .A1(n3394), .A2(n4196), .ZN(n2704) );
  OAI211_X1 U3106 ( .C1(n3228), .C2(n2705), .A(n3227), .B(n2704), .ZN(n4137)
         );
  NAND2_X1 U3107 ( .A1(n3615), .A2(n4137), .ZN(n2707) );
  OR2_X1 U3108 ( .A1(n3979), .A2(n2705), .ZN(n2706) );
  OAI211_X1 U3109 ( .C1(n3570), .C2(n2708), .A(n2707), .B(n2706), .ZN(n2709)
         );
  NOR2_X1 U3110 ( .A1(n2710), .A2(n2709), .ZN(n2711) );
  NAND4_X1 U3111 ( .A1(n2714), .A2(n2713), .A3(n2712), .A4(n2711), .ZN(n2715)
         );
  NOR2_X1 U3112 ( .A1(n3623), .A2(n2715), .ZN(n2721) );
  INV_X1 U3113 ( .A(is_clpx_i), .ZN(n2950) );
  OAI21_X1 U3114 ( .B1(n2950), .B2(n2949), .A(n2944), .ZN(n3432) );
  INV_X1 U3115 ( .A(n3432), .ZN(n2716) );
  OAI21_X1 U3116 ( .B1(n3437), .B2(n2717), .A(n2716), .ZN(n3626) );
  OR2_X1 U3117 ( .A1(n2733), .A2(n3683), .ZN(n3990) );
  OR3_X1 U3118 ( .A1(n2495), .A2(n2745), .A3(n3351), .ZN(n4021) );
  MUX2_X1 U3119 ( .A(n4038), .B(n4021), .S(n4196), .Z(n2718) );
  OAI21_X1 U3120 ( .B1(n2735), .B2(n3990), .A(n2718), .ZN(n2719) );
  OAI21_X1 U3121 ( .B1(n3626), .B2(n2719), .A(n149), .ZN(n2720) );
  NAND3_X1 U3122 ( .A1(n2722), .A2(n2721), .A3(n2720), .ZN(n2723) );
  NOR2_X1 U3123 ( .A1(n2724), .A2(n2723), .ZN(n2731) );
  NOR2_X1 U3124 ( .A1(n2726), .A2(n2725), .ZN(n4012) );
  NAND2_X1 U3125 ( .A1(n4012), .A2(n2727), .ZN(n4182) );
  INV_X1 U3126 ( .A(n4182), .ZN(n3944) );
  NAND2_X1 U3127 ( .A1(n4365), .A2(n3944), .ZN(n2730) );
  INV_X1 U3128 ( .A(n2728), .ZN(n4121) );
  INV_X1 U3129 ( .A(n4121), .ZN(n4014) );
  NAND2_X1 U3130 ( .A1(n3280), .A2(n4014), .ZN(n2729) );
  NOR2_X2 U3131 ( .A1(n2733), .A2(n4161), .ZN(n4007) );
  NAND2_X1 U3132 ( .A1(n222), .A2(n4007), .ZN(n2734) );
  NAND2_X1 U3133 ( .A1(n2734), .A2(n4151), .ZN(n2736) );
  NAND2_X1 U3134 ( .A1(n2736), .A2(n2735), .ZN(n2737) );
  NAND2_X1 U3135 ( .A1(n2739), .A2(n2738), .ZN(result_o[8]) );
  INV_X1 U3136 ( .A(n4163), .ZN(n2741) );
  INV_X1 U3138 ( .A(n4160), .ZN(n2744) );
  OR2_X1 U3139 ( .A1(n2745), .A2(n2744), .ZN(n3370) );
  MUX2_X1 U3140 ( .A(n3370), .B(n2902), .S(n2770), .Z(n2762) );
  NAND2_X1 U3141 ( .A1(n2747), .A2(n2753), .ZN(n2746) );
  OAI21_X1 U3142 ( .B1(n2748), .B2(n2747), .A(n2746), .ZN(n2758) );
  BUF_X1 U3143 ( .A(n61), .Z(n2750) );
  INV_X1 U3144 ( .A(n2750), .ZN(n2755) );
  INV_X1 U3145 ( .A(n2753), .ZN(n2754) );
  AOI21_X1 U3146 ( .B1(n2758), .B2(n2757), .A(n2756), .ZN(n2761) );
  NAND2_X1 U3148 ( .A1(n3463), .A2(n4007), .ZN(n2764) );
  NAND2_X1 U3149 ( .A1(n2764), .A2(n4151), .ZN(n2766) );
  INV_X1 U3150 ( .A(operand_c_i[29]), .ZN(n2822) );
  INV_X1 U3152 ( .A(n3853), .ZN(n3490) );
  INV_X1 U3153 ( .A(n4059), .ZN(n4192) );
  INV_X1 U3154 ( .A(n3820), .ZN(n3793) );
  AOI22_X1 U3155 ( .A1(n3944), .A2(n3875), .B1(n3463), .B2(n4014), .ZN(n2841)
         );
  NAND2_X1 U3156 ( .A1(n2769), .A2(n2767), .ZN(n3358) );
  NAND2_X1 U3157 ( .A1(n2769), .A2(n2768), .ZN(n3359) );
  MUX2_X1 U3158 ( .A(n3358), .B(n3359), .S(n161), .Z(n2833) );
  NAND2_X1 U3159 ( .A1(n2833), .A2(n3443), .ZN(n2771) );
  AND2_X1 U3160 ( .A1(n3446), .A2(n2771), .ZN(n4016) );
  MUX2_X1 U3161 ( .A(n4017), .B(n4016), .S(operand_b_i[29]), .Z(n2839) );
  INV_X1 U3162 ( .A(n2833), .ZN(n2772) );
  OAI21_X1 U3163 ( .B1(n3437), .B2(n2772), .A(n2944), .ZN(n4023) );
  INV_X1 U3164 ( .A(n3990), .ZN(n4126) );
  NAND2_X1 U3165 ( .A1(n2773), .A2(n4126), .ZN(n2774) );
  OAI21_X1 U3166 ( .B1(n4021), .B2(n2775), .A(n2774), .ZN(n2776) );
  OAI21_X1 U3167 ( .B1(n4023), .B2(n2776), .A(n54), .ZN(n2837) );
  AND2_X1 U3168 ( .A1(n2784), .A2(n3385), .ZN(n2779) );
  OAI21_X1 U3169 ( .B1(n2777), .B2(n4328), .A(n3386), .ZN(n2778) );
  AOI21_X1 U3170 ( .B1(n3396), .B2(n2779), .A(n2778), .ZN(n2780) );
  OAI21_X1 U3171 ( .B1(n3393), .B2(imm_vec_ext_i[1]), .A(n2780), .ZN(n2908) );
  NOR2_X1 U3172 ( .A1(n3391), .A2(n170), .ZN(n2781) );
  OR3_X1 U3173 ( .A1(n2782), .A2(n2908), .A3(n2781), .ZN(n2816) );
  AND2_X1 U3174 ( .A1(n3387), .A2(n4131), .ZN(n2783) );
  NAND2_X1 U3175 ( .A1(n3394), .A2(n2783), .ZN(n4040) );
  NAND2_X1 U3176 ( .A1(n3407), .A2(n4040), .ZN(n2909) );
  OR2_X1 U3177 ( .A1(n2816), .A2(n2909), .ZN(n2825) );
  INV_X1 U3178 ( .A(n2825), .ZN(n2799) );
  NOR2_X1 U3179 ( .A1(n2794), .A2(n3765), .ZN(n2785) );
  OAI21_X1 U3180 ( .B1(n2786), .B2(n2785), .A(n2784), .ZN(n2789) );
  NAND3_X1 U3181 ( .A1(n2789), .A2(n2788), .A3(n2787), .ZN(n2914) );
  INV_X1 U3182 ( .A(n3382), .ZN(n2790) );
  NOR2_X1 U3183 ( .A1(n2790), .A2(n4020), .ZN(n2791) );
  OR2_X1 U3184 ( .A1(n2914), .A2(n2791), .ZN(n2815) );
  INV_X1 U3185 ( .A(n2815), .ZN(n2792) );
  NAND2_X1 U3186 ( .A1(n2799), .A2(n2792), .ZN(n2812) );
  NAND2_X1 U3187 ( .A1(vector_mode_i[1]), .A2(n4340), .ZN(n2793) );
  NOR2_X1 U3188 ( .A1(n2794), .A2(n2793), .ZN(n2795) );
  NOR2_X1 U3189 ( .A1(n2796), .A2(n2795), .ZN(n2814) );
  OR2_X1 U3190 ( .A1(n2812), .A2(n2814), .ZN(n4034) );
  NAND3_X1 U3191 ( .A1(n3076), .A2(vector_mode_i[0]), .A3(n4079), .ZN(n2798)
         );
  NAND2_X1 U3192 ( .A1(n3393), .A2(n4101), .ZN(n2797) );
  NAND2_X1 U3193 ( .A1(n2798), .A2(n2797), .ZN(n3561) );
  INV_X1 U3194 ( .A(n2814), .ZN(n2801) );
  AND2_X1 U3195 ( .A1(n2815), .A2(n2801), .ZN(n2804) );
  NAND2_X1 U3196 ( .A1(n2799), .A2(n2804), .ZN(n3537) );
  INV_X1 U3197 ( .A(n3537), .ZN(n4027) );
  OR2_X1 U3198 ( .A1(n3076), .A2(n53), .ZN(n2800) );
  OAI21_X1 U3199 ( .B1(n3561), .B2(n3225), .A(n2800), .ZN(n3732) );
  NOR2_X1 U3200 ( .A1(n2815), .A2(n2801), .ZN(n2802) );
  AND2_X1 U3201 ( .A1(n2802), .A2(n2816), .ZN(n4025) );
  INV_X1 U3202 ( .A(operand_c_i[5]), .ZN(n3728) );
  NAND2_X1 U3203 ( .A1(n3394), .A2(operand_b_i[5]), .ZN(n2803) );
  OAI211_X1 U3204 ( .C1(n3228), .C2(n3728), .A(n3223), .B(n2803), .ZN(n3726)
         );
  AOI22_X1 U3205 ( .A1(n4027), .A2(n3732), .B1(n4025), .B2(n3726), .ZN(n2811)
         );
  AND2_X1 U3206 ( .A1(n2804), .A2(n2816), .ZN(n4031) );
  NOR2_X1 U3207 ( .A1(n3228), .A2(n2822), .ZN(n2807) );
  NAND2_X1 U3208 ( .A1(n3394), .A2(operand_b_i[29]), .ZN(n2805) );
  NAND2_X1 U3209 ( .A1(n3219), .A2(n2805), .ZN(n2806) );
  NOR2_X1 U3210 ( .A1(n2807), .A2(n2806), .ZN(n3723) );
  INV_X1 U3211 ( .A(n3723), .ZN(n3560) );
  NOR2_X1 U3212 ( .A1(n2815), .A2(n2814), .ZN(n2808) );
  AND2_X1 U3213 ( .A1(n2808), .A2(n2816), .ZN(n4029) );
  INV_X1 U3214 ( .A(operand_c_i[13]), .ZN(n3565) );
  NAND2_X1 U3215 ( .A1(n3394), .A2(operand_b_i[13]), .ZN(n2809) );
  OAI211_X1 U3216 ( .C1(n3228), .C2(n3565), .A(n3227), .B(n2809), .ZN(n3725)
         );
  AOI22_X1 U3217 ( .A1(n4031), .A2(n3560), .B1(n4029), .B2(n3725), .ZN(n2810)
         );
  OAI211_X1 U3218 ( .C1(n4034), .C2(n3561), .A(n2811), .B(n2810), .ZN(n2831)
         );
  INV_X1 U3219 ( .A(n2812), .ZN(n2813) );
  AND2_X1 U3220 ( .A1(n2813), .A2(n2814), .ZN(n4036) );
  NAND2_X1 U3221 ( .A1(n4036), .A2(operand_a_i[5]), .ZN(n2829) );
  NAND2_X1 U3222 ( .A1(n2815), .A2(n2814), .ZN(n2824) );
  INV_X1 U3223 ( .A(n2824), .ZN(n2817) );
  AND2_X1 U3224 ( .A1(n2817), .A2(n2816), .ZN(n4043) );
  INV_X1 U3225 ( .A(operand_c_i[21]), .ZN(n3262) );
  NOR2_X1 U3226 ( .A1(n3228), .A2(n3262), .ZN(n2820) );
  NAND2_X1 U3227 ( .A1(n3394), .A2(operand_b_i[21]), .ZN(n2818) );
  NAND2_X1 U3228 ( .A1(n3221), .A2(n2818), .ZN(n2819) );
  NOR2_X1 U3229 ( .A1(n2820), .A2(n2819), .ZN(n3720) );
  INV_X1 U3230 ( .A(n3720), .ZN(n3559) );
  OAI22_X1 U3231 ( .A1(n4040), .A2(n2822), .B1(n4038), .B2(n2821), .ZN(n2823)
         );
  AOI21_X1 U3232 ( .B1(n4043), .B2(n3559), .A(n2823), .ZN(n2828) );
  NOR2_X1 U3233 ( .A1(n2825), .A2(n2824), .ZN(n4045) );
  NAND2_X1 U3234 ( .A1(n3076), .A2(operand_a_i[5]), .ZN(n2826) );
  OAI21_X1 U3235 ( .B1(n3076), .B2(n4075), .A(n2826), .ZN(n3731) );
  NAND2_X1 U3236 ( .A1(n4045), .A2(n3731), .ZN(n2827) );
  NAND3_X1 U3237 ( .A1(n2829), .A2(n2828), .A3(n2827), .ZN(n2830) );
  NOR2_X1 U3238 ( .A1(n2831), .A2(n2830), .ZN(n2836) );
  NAND2_X1 U3239 ( .A1(n2832), .A2(n2903), .ZN(n4054) );
  AOI21_X1 U3240 ( .B1(n2833), .B2(n2950), .A(n2949), .ZN(n4052) );
  NAND2_X1 U3241 ( .A1(n4052), .A2(n2834), .ZN(n2835) );
  NAND4_X1 U3242 ( .A1(n2837), .A2(n2836), .A3(n4054), .A4(n2835), .ZN(n2838)
         );
  AOI211_X1 U3243 ( .C1(result_div[29]), .C2(n3988), .A(n2839), .B(n2838), 
        .ZN(n2840) );
  OAI211_X1 U3244 ( .C1(n3793), .C2(n4184), .A(n2841), .B(n2840), .ZN(n2842)
         );
  INV_X1 U3245 ( .A(n2842), .ZN(n2843) );
  INV_X1 U3246 ( .A(operand_c_i[27]), .ZN(n2858) );
  INV_X1 U3250 ( .A(n2846), .ZN(n3753) );
  MUX2_X1 U3251 ( .A(n4017), .B(n4016), .S(n64), .Z(n2869) );
  NAND2_X1 U3252 ( .A1(n2875), .A2(n4126), .ZN(n2847) );
  OAI21_X1 U3253 ( .B1(n4021), .B2(n2848), .A(n2847), .ZN(n2849) );
  OAI21_X1 U3254 ( .B1(n4023), .B2(n2849), .A(operand_a_i[27]), .ZN(n2867) );
  MUX2_X1 U3255 ( .A(n48), .B(operand_a_i[11]), .S(n3393), .Z(n3602) );
  NOR2_X1 U3256 ( .A1(n3076), .A2(n2521), .ZN(n2850) );
  AOI21_X1 U3257 ( .B1(n3602), .B2(n3076), .A(n2850), .ZN(n3472) );
  NAND2_X1 U3258 ( .A1(n4036), .A2(n48), .ZN(n2855) );
  INV_X1 U3259 ( .A(operand_c_i[19]), .ZN(n3013) );
  NAND2_X1 U3260 ( .A1(n3394), .A2(operand_b_i[19]), .ZN(n2851) );
  OAI211_X1 U3261 ( .C1(n3228), .C2(n3013), .A(n3221), .B(n2851), .ZN(n3616)
         );
  OAI22_X1 U3262 ( .A1(n4040), .A2(n2858), .B1(n4038), .B2(n2852), .ZN(n2853)
         );
  AOI21_X1 U3263 ( .B1(n4043), .B2(n3616), .A(n2853), .ZN(n2854) );
  OAI211_X1 U3264 ( .C1(n3472), .C2(n3537), .A(n2855), .B(n2854), .ZN(n2863)
         );
  INV_X1 U3265 ( .A(n3602), .ZN(n3017) );
  MUX2_X1 U3266 ( .A(operand_a_i[19]), .B(n48), .S(n3076), .Z(n3603) );
  INV_X1 U3267 ( .A(operand_c_i[11]), .ZN(n3608) );
  NAND2_X1 U3268 ( .A1(n3394), .A2(n150), .ZN(n2856) );
  OAI211_X1 U3269 ( .C1(n3228), .C2(n3608), .A(n3227), .B(n2856), .ZN(n3614)
         );
  AOI22_X1 U3270 ( .A1(n4045), .A2(n3603), .B1(n4029), .B2(n3614), .ZN(n2861)
         );
  NAND2_X1 U3271 ( .A1(n3394), .A2(n64), .ZN(n2857) );
  OAI211_X1 U3272 ( .C1(n3228), .C2(n2858), .A(n3219), .B(n2857), .ZN(n3605)
         );
  INV_X1 U3273 ( .A(operand_c_i[3]), .ZN(n3468) );
  NAND2_X1 U3274 ( .A1(n3394), .A2(operand_b_i[3]), .ZN(n2859) );
  OAI211_X1 U3275 ( .C1(n3228), .C2(n3468), .A(n3223), .B(n2859), .ZN(n3597)
         );
  AOI22_X1 U3276 ( .A1(n4031), .A2(n3605), .B1(n4025), .B2(n3597), .ZN(n2860)
         );
  OAI211_X1 U3277 ( .C1(n4034), .C2(n3017), .A(n2861), .B(n2860), .ZN(n2862)
         );
  NOR2_X1 U3278 ( .A1(n2863), .A2(n2862), .ZN(n2866) );
  NAND2_X1 U3279 ( .A1(n4052), .A2(n2864), .ZN(n2865) );
  NAND4_X1 U3280 ( .A1(n2867), .A2(n2866), .A3(n4054), .A4(n2865), .ZN(n2868)
         );
  AOI211_X1 U3281 ( .C1(result_div[27]), .C2(n3988), .A(n2869), .B(n2868), 
        .ZN(n2870) );
  INV_X1 U3282 ( .A(n2870), .ZN(n2871) );
  AOI21_X1 U3283 ( .B1(n3821), .B2(n4014), .A(n2871), .ZN(n2873) );
  AOI22_X1 U3284 ( .A1(n3875), .A2(n3750), .B1(n3944), .B2(n3820), .ZN(n2872)
         );
  OAI211_X1 U3285 ( .C1(n3753), .C2(n4192), .A(n2873), .B(n2872), .ZN(n2879)
         );
  AOI21_X1 U3286 ( .B1(n3821), .B2(n4007), .A(n4006), .ZN(n2874) );
  INV_X1 U3287 ( .A(n2874), .ZN(n2877) );
  INV_X1 U3289 ( .A(operand_c_i[23]), .ZN(n2921) );
  NAND2_X1 U3292 ( .A1(n4365), .A2(n4007), .ZN(n2883) );
  NAND2_X1 U3293 ( .A1(n2883), .A2(n4151), .ZN(n2884) );
  AOI22_X1 U3294 ( .A1(n125), .A2(n3750), .B1(n3521), .B2(n4059), .ZN(n2961)
         );
  NAND2_X1 U3295 ( .A1(n2888), .A2(n3387), .ZN(n2889) );
  AND2_X1 U3296 ( .A1(n2890), .A2(n2889), .ZN(n2894) );
  INV_X1 U3297 ( .A(n2894), .ZN(n2901) );
  OR2_X1 U3298 ( .A1(n3358), .A2(n2901), .ZN(n2891) );
  OAI21_X1 U3299 ( .B1(n3359), .B2(n2894), .A(n2891), .ZN(n2948) );
  OAI21_X1 U3300 ( .B1(n2892), .B2(n2948), .A(n3446), .ZN(n3890) );
  MUX2_X1 U3301 ( .A(n4179), .B(n3890), .S(operand_b_i[23]), .Z(n2956) );
  INV_X1 U3302 ( .A(n2893), .ZN(n3368) );
  AOI21_X1 U3303 ( .B1(n2894), .B2(n3361), .A(n3373), .ZN(n2900) );
  NOR2_X1 U3304 ( .A1(n2896), .A2(n3363), .ZN(n2897) );
  NOR2_X1 U3305 ( .A1(n2898), .A2(n2897), .ZN(n2899) );
  MUX2_X1 U3306 ( .A(n3368), .B(n2900), .S(n2899), .Z(n2905) );
  MUX2_X1 U3307 ( .A(n3370), .B(n2902), .S(n2901), .Z(n2904) );
  INV_X1 U3308 ( .A(n2903), .ZN(n3374) );
  AOI21_X1 U3309 ( .B1(n2905), .B2(n2904), .A(n3374), .ZN(n3917) );
  NOR2_X1 U3310 ( .A1(n3391), .A2(n4194), .ZN(n2907) );
  OAI21_X1 U3311 ( .B1(n3393), .B2(n3385), .A(n3979), .ZN(n2906) );
  OR3_X1 U3312 ( .A1(n2908), .A2(n2907), .A3(n2906), .ZN(n2931) );
  NOR2_X1 U3313 ( .A1(n2931), .A2(n2909), .ZN(n2937) );
  INV_X1 U3314 ( .A(n2937), .ZN(n2912) );
  NAND2_X1 U3315 ( .A1(n3382), .A2(operand_b_i[16]), .ZN(n2911) );
  AND2_X1 U3316 ( .A1(n2911), .A2(n2910), .ZN(n2929) );
  INV_X1 U3317 ( .A(n2929), .ZN(n2926) );
  NOR2_X1 U3318 ( .A1(n2912), .A2(n2926), .ZN(n2934) );
  INV_X1 U3319 ( .A(n2934), .ZN(n2915) );
  AND2_X1 U3320 ( .A1(n3382), .A2(n4328), .ZN(n2913) );
  OR2_X1 U3321 ( .A1(n2914), .A2(n2913), .ZN(n2933) );
  OR2_X1 U3322 ( .A1(n2915), .A2(n2933), .ZN(n3901) );
  NOR2_X1 U3323 ( .A1(n3901), .A2(n2543), .ZN(n2925) );
  MUX2_X1 U3324 ( .A(operand_a_i[7]), .B(operand_a_i[15]), .S(n3393), .Z(n3970) );
  INV_X1 U3325 ( .A(n3970), .ZN(n3948) );
  NOR2_X1 U3326 ( .A1(n2933), .A2(n2929), .ZN(n2916) );
  NAND2_X1 U3327 ( .A1(n2937), .A2(n2916), .ZN(n3911) );
  AND2_X1 U3328 ( .A1(n2916), .A2(n2931), .ZN(n3906) );
  INV_X1 U3329 ( .A(operand_c_i[15]), .ZN(n3044) );
  NAND2_X1 U3330 ( .A1(n3394), .A2(operand_b_i[15]), .ZN(n2917) );
  OAI211_X1 U3331 ( .C1(n3228), .C2(n3044), .A(n3227), .B(n2917), .ZN(n3981)
         );
  OAI22_X1 U3332 ( .A1(n4040), .A2(n2921), .B1(n4038), .B2(n2918), .ZN(n2919)
         );
  AOI21_X1 U3333 ( .B1(n3906), .B2(n3981), .A(n2919), .ZN(n2923) );
  AND3_X1 U3334 ( .A1(n2931), .A2(n2929), .A3(n2933), .ZN(n3908) );
  NAND2_X1 U3335 ( .A1(n3394), .A2(operand_b_i[23]), .ZN(n2920) );
  OAI211_X1 U3336 ( .C1(n3228), .C2(n2921), .A(n3221), .B(n2920), .ZN(n3971)
         );
  NAND2_X1 U3337 ( .A1(n3908), .A2(n3971), .ZN(n2922) );
  OAI211_X1 U3338 ( .C1(n3948), .C2(n3911), .A(n2923), .B(n2922), .ZN(n2924)
         );
  NOR2_X1 U3339 ( .A1(n2925), .A2(n2924), .ZN(n2942) );
  NAND2_X1 U3340 ( .A1(n2933), .A2(n2926), .ZN(n2935) );
  INV_X1 U3341 ( .A(n2931), .ZN(n2927) );
  OR2_X1 U3342 ( .A1(n2935), .A2(n2927), .ZN(n3770) );
  INV_X1 U3343 ( .A(n3770), .ZN(n3896) );
  INV_X1 U3344 ( .A(operand_c_i[31]), .ZN(n3937) );
  NAND2_X1 U3345 ( .A1(n3394), .A2(operand_b_i[31]), .ZN(n2928) );
  OAI211_X1 U3346 ( .C1(n3228), .C2(n3937), .A(n3219), .B(n2928), .ZN(n3975)
         );
  INV_X1 U3347 ( .A(n2933), .ZN(n2930) );
  AND3_X1 U3348 ( .A1(n2931), .A2(n2930), .A3(n2929), .ZN(n3894) );
  INV_X1 U3349 ( .A(operand_c_i[7]), .ZN(n3978) );
  NAND2_X1 U3350 ( .A1(n3394), .A2(operand_b_i[7]), .ZN(n2932) );
  OAI211_X1 U3351 ( .C1(n3228), .C2(n3978), .A(n3223), .B(n2932), .ZN(n3974)
         );
  AOI22_X1 U3352 ( .A1(n3896), .A2(n3975), .B1(n3894), .B2(n3974), .ZN(n2941)
         );
  AND2_X1 U3353 ( .A1(n2934), .A2(n2933), .ZN(n3892) );
  MUX2_X1 U3354 ( .A(n585), .B(n2543), .S(n3076), .Z(n3048) );
  INV_X1 U3355 ( .A(n3048), .ZN(n3972) );
  NAND2_X1 U3356 ( .A1(n3892), .A2(n3972), .ZN(n2940) );
  INV_X1 U3357 ( .A(n2935), .ZN(n2936) );
  NAND2_X1 U3358 ( .A1(n2937), .A2(n2936), .ZN(n3899) );
  NOR2_X1 U3359 ( .A1(n3076), .A2(n4115), .ZN(n2938) );
  AOI21_X1 U3360 ( .B1(n3970), .B2(n3076), .A(n2938), .ZN(n3945) );
  OR2_X1 U3361 ( .A1(n3899), .A2(n3945), .ZN(n2939) );
  NAND4_X1 U3362 ( .A1(n2942), .A2(n2941), .A3(n2940), .A4(n2939), .ZN(n2943)
         );
  NOR2_X1 U3363 ( .A1(n3917), .A2(n2943), .ZN(n2955) );
  OAI21_X1 U3364 ( .B1(n3437), .B2(n2948), .A(n2944), .ZN(n3921) );
  OAI22_X1 U3365 ( .A1(n2946), .A2(n3990), .B1(n2505), .B2(n4021), .ZN(n2947)
         );
  OAI21_X1 U3366 ( .B1(n3921), .B2(n2947), .A(operand_a_i[23]), .ZN(n2954) );
  INV_X1 U3367 ( .A(n2948), .ZN(n2951) );
  AOI21_X1 U3368 ( .B1(n2951), .B2(n2950), .A(n169), .ZN(n3923) );
  NAND2_X1 U3369 ( .A1(n3923), .A2(n2952), .ZN(n2953) );
  NAND4_X1 U3370 ( .A1(n2956), .A2(n2955), .A3(n2954), .A4(n2953), .ZN(n2957)
         );
  AOI21_X1 U3371 ( .B1(result_div[23]), .B2(n3988), .A(n2957), .ZN(n2960) );
  NAND2_X1 U3372 ( .A1(n222), .A2(n3944), .ZN(n2959) );
  NAND2_X1 U3373 ( .A1(n4365), .A2(n4014), .ZN(n2958) );
  NAND4_X1 U3374 ( .A1(n2961), .A2(n2960), .A3(n2959), .A4(n2958), .ZN(n2962)
         );
  INV_X1 U3376 ( .A(operand_c_i[17]), .ZN(n2980) );
  INV_X1 U3379 ( .A(n3788), .ZN(n3104) );
  INV_X1 U3380 ( .A(n2968), .ZN(n3759) );
  INV_X1 U3381 ( .A(n3921), .ZN(n2970) );
  INV_X1 U3382 ( .A(n4021), .ZN(n4125) );
  AOI22_X1 U3383 ( .A1(n3000), .A2(n4126), .B1(n4328), .B2(n4125), .ZN(n2969)
         );
  AOI21_X1 U3384 ( .B1(n2970), .B2(n2969), .A(n538), .ZN(n2993) );
  MUX2_X1 U3385 ( .A(n4179), .B(n3890), .S(n4328), .Z(n2991) );
  MUX2_X1 U3386 ( .A(n4225), .B(operand_a_i[9]), .S(n3393), .Z(n3687) );
  OR2_X1 U3387 ( .A1(n3076), .A2(operand_a_i[25]), .ZN(n2971) );
  OAI21_X1 U3388 ( .B1(n3687), .B2(n3225), .A(n2971), .ZN(n3688) );
  MUX2_X1 U3389 ( .A(operand_a_i[17]), .B(n4225), .S(n3076), .Z(n4044) );
  NAND2_X1 U3390 ( .A1(n3892), .A2(n4044), .ZN(n2975) );
  INV_X1 U3391 ( .A(operand_c_i[25]), .ZN(n4039) );
  NAND2_X1 U3392 ( .A1(n3394), .A2(n110), .ZN(n2972) );
  OAI211_X1 U3393 ( .C1(n3228), .C2(n4039), .A(n3219), .B(n2972), .ZN(n4030)
         );
  INV_X1 U3394 ( .A(operand_c_i[1]), .ZN(n3682) );
  NAND2_X1 U3395 ( .A1(n3394), .A2(operand_b_i[1]), .ZN(n2973) );
  OAI211_X1 U3396 ( .C1(n3228), .C2(n3682), .A(n3223), .B(n2973), .ZN(n4024)
         );
  AOI22_X1 U3397 ( .A1(n3896), .A2(n4030), .B1(n3894), .B2(n4024), .ZN(n2974)
         );
  OAI211_X1 U3398 ( .C1(n3688), .C2(n3899), .A(n2975), .B(n2974), .ZN(n2986)
         );
  NOR2_X1 U3399 ( .A1(n3901), .A2(n2546), .ZN(n2984) );
  INV_X1 U3400 ( .A(n3687), .ZN(n4035) );
  INV_X1 U3401 ( .A(operand_c_i[9]), .ZN(n3500) );
  NAND2_X1 U3402 ( .A1(n3394), .A2(n4195), .ZN(n2976) );
  OAI211_X1 U3403 ( .C1(n3228), .C2(n3500), .A(n3227), .B(n2976), .ZN(n4028)
         );
  OAI22_X1 U3404 ( .A1(n4040), .A2(n2980), .B1(n4038), .B2(n2977), .ZN(n2978)
         );
  AOI21_X1 U3405 ( .B1(n3906), .B2(n4028), .A(n2978), .ZN(n2982) );
  NAND2_X1 U3406 ( .A1(n3394), .A2(n4328), .ZN(n2979) );
  OAI211_X1 U3407 ( .C1(n3228), .C2(n2980), .A(n3221), .B(n2979), .ZN(n4042)
         );
  NAND2_X1 U3408 ( .A1(n3908), .A2(n4042), .ZN(n2981) );
  OAI211_X1 U3409 ( .C1(n3911), .C2(n4035), .A(n2982), .B(n2981), .ZN(n2983)
         );
  OR2_X1 U3410 ( .A1(n2984), .A2(n2983), .ZN(n2985) );
  NOR2_X1 U3411 ( .A1(n2986), .A2(n2985), .ZN(n2990) );
  NAND2_X1 U3412 ( .A1(n3923), .A2(n2987), .ZN(n2989) );
  INV_X1 U3413 ( .A(n3917), .ZN(n2988) );
  NAND4_X1 U3414 ( .A1(n2991), .A2(n2990), .A3(n2989), .A4(n2988), .ZN(n2992)
         );
  AOI211_X1 U3415 ( .C1(result_div[17]), .C2(n3988), .A(n2993), .B(n2992), 
        .ZN(n2996) );
  NAND2_X1 U3416 ( .A1(n3763), .A2(n4059), .ZN(n2995) );
  OAI211_X1 U3417 ( .C1(n3759), .C2(n4184), .A(n2996), .B(n2995), .ZN(n2997)
         );
  AOI21_X1 U3418 ( .B1(n4014), .B2(n3216), .A(n2997), .ZN(n2998) );
  OAI21_X1 U3419 ( .B1(n3104), .B2(n4182), .A(n2998), .ZN(n3004) );
  AOI21_X1 U3420 ( .B1(n3216), .B2(n4007), .A(n4006), .ZN(n2999) );
  INV_X1 U3421 ( .A(n2999), .ZN(n3002) );
  NAND2_X1 U3422 ( .A1(n3006), .A2(n3005), .ZN(result_o[17]) );
  INV_X1 U3425 ( .A(n3217), .ZN(n3008) );
  INV_X1 U3426 ( .A(n4007), .ZN(n4122) );
  OAI21_X1 U3427 ( .B1(n3008), .B2(n4122), .A(n4151), .ZN(n3009) );
  MUX2_X1 U3428 ( .A(n4179), .B(n3890), .S(operand_b_i[19]), .Z(n3031) );
  NOR2_X1 U3429 ( .A1(n3901), .A2(n3011), .ZN(n3019) );
  OAI22_X1 U3430 ( .A1(n4040), .A2(n3013), .B1(n4038), .B2(n3012), .ZN(n3014)
         );
  AOI21_X1 U3431 ( .B1(n3906), .B2(n3614), .A(n3014), .ZN(n3016) );
  NAND2_X1 U3432 ( .A1(n3908), .A2(n3616), .ZN(n3015) );
  OAI211_X1 U3433 ( .C1(n3017), .C2(n3911), .A(n3016), .B(n3015), .ZN(n3018)
         );
  NOR2_X1 U3434 ( .A1(n3019), .A2(n3018), .ZN(n3023) );
  AOI22_X1 U3435 ( .A1(n3896), .A2(n3605), .B1(n3894), .B2(n3597), .ZN(n3022)
         );
  NAND2_X1 U3436 ( .A1(n3892), .A2(n3603), .ZN(n3021) );
  OR2_X1 U3437 ( .A1(n3899), .A2(n3472), .ZN(n3020) );
  NAND4_X1 U3438 ( .A1(n3023), .A2(n3022), .A3(n3021), .A4(n3020), .ZN(n3024)
         );
  NOR2_X1 U3439 ( .A1(n3917), .A2(n3024), .ZN(n3030) );
  INV_X1 U3440 ( .A(n4125), .ZN(n3989) );
  OAI22_X1 U3441 ( .A1(n3026), .A2(n3990), .B1(n3025), .B2(n3989), .ZN(n3027)
         );
  OAI21_X1 U3442 ( .B1(n3921), .B2(n3027), .A(operand_a_i[19]), .ZN(n3029) );
  NAND4_X1 U3443 ( .A1(n3031), .A2(n3030), .A3(n3029), .A4(n3028), .ZN(n3032)
         );
  AOI21_X1 U3444 ( .B1(result_div[19]), .B2(n3988), .A(n3032), .ZN(n3033) );
  INV_X1 U3445 ( .A(n3033), .ZN(n3034) );
  AOI21_X1 U3446 ( .B1(n3590), .B2(n4059), .A(n3034), .ZN(n3036) );
  NAND2_X1 U3447 ( .A1(n4309), .A2(n4012), .ZN(n3035) );
  OAI211_X1 U3448 ( .C1(n4121), .C2(n3008), .A(n3036), .B(n3035), .ZN(n3037)
         );
  NAND2_X1 U3452 ( .A1(result_div[15]), .A2(n3988), .ZN(n3060) );
  AOI22_X1 U3453 ( .A1(n3606), .A2(n3975), .B1(n3617), .B2(n3971), .ZN(n3053)
         );
  AOI22_X1 U3454 ( .A1(n3970), .A2(n3601), .B1(n3598), .B2(n3974), .ZN(n3052)
         );
  OAI22_X1 U3455 ( .A1(n3945), .A2(n3562), .B1(n3612), .B2(n2543), .ZN(n3050)
         );
  NAND2_X1 U3456 ( .A1(n3615), .A2(n3981), .ZN(n3047) );
  OAI22_X1 U3457 ( .A1(n3979), .A2(n3044), .B1(n4038), .B2(n3042), .ZN(n3045)
         );
  INV_X1 U3458 ( .A(n3045), .ZN(n3046) );
  OAI211_X1 U3459 ( .C1(n3570), .C2(n3048), .A(n3047), .B(n3046), .ZN(n3049)
         );
  NOR2_X1 U3460 ( .A1(n3050), .A2(n3049), .ZN(n3051) );
  NAND4_X1 U3461 ( .A1(n3576), .A2(n3053), .A3(n3052), .A4(n3051), .ZN(n3054)
         );
  MUX2_X1 U3462 ( .A(n4179), .B(n3596), .S(operand_b_i[15]), .Z(n3058) );
  OAI22_X1 U3463 ( .A1(n3067), .A2(n3990), .B1(n3055), .B2(n3989), .ZN(n3056)
         );
  OAI21_X1 U3464 ( .B1(n3626), .B2(n3056), .A(operand_a_i[15]), .ZN(n3057) );
  NAND4_X1 U3465 ( .A1(n3060), .A2(n3059), .A3(n3058), .A4(n3057), .ZN(n3061)
         );
  AOI21_X1 U3466 ( .B1(n3763), .B2(n4014), .A(n3061), .ZN(n3062) );
  OAI21_X1 U3467 ( .B1(n3759), .B2(n4182), .A(n3062), .ZN(n3063) );
  AOI21_X1 U3468 ( .B1(n4059), .B2(n3216), .A(n3063), .ZN(n3064) );
  OAI21_X1 U3469 ( .B1(n3104), .B2(n4184), .A(n3064), .ZN(n3070) );
  NAND2_X1 U3470 ( .A1(n3763), .A2(n4007), .ZN(n3065) );
  NAND2_X1 U3471 ( .A1(n3065), .A2(n4151), .ZN(n3068) );
  AND2_X1 U3472 ( .A1(n3068), .A2(n3067), .ZN(n3069) );
  NAND2_X1 U3473 ( .A1(n3072), .A2(n3071), .ZN(result_o[15]) );
  INV_X1 U3474 ( .A(operand_c_i[14]), .ZN(n3086) );
  MUX2_X1 U3477 ( .A(n4179), .B(n3596), .S(operand_b_i[14]), .Z(n3099) );
  INV_X1 U3478 ( .A(n3562), .ZN(n3600) );
  MUX2_X1 U3479 ( .A(n4071), .B(n4098), .S(n3393), .Z(n3294) );
  OR2_X1 U3480 ( .A1(n3076), .A2(n4112), .ZN(n3074) );
  OAI21_X1 U3481 ( .B1(n3294), .B2(n3225), .A(n3074), .ZN(n3645) );
  INV_X1 U3482 ( .A(operand_c_i[6]), .ZN(n3655) );
  NAND2_X1 U3483 ( .A1(n3394), .A2(operand_b_i[6]), .ZN(n3075) );
  OAI211_X1 U3484 ( .C1(n3228), .C2(n3655), .A(n3223), .B(n3075), .ZN(n3647)
         );
  AOI22_X1 U3485 ( .A1(n3600), .A2(n3645), .B1(n3598), .B2(n3647), .ZN(n3090)
         );
  INV_X1 U3486 ( .A(n3570), .ZN(n3604) );
  MUX2_X1 U3487 ( .A(n4072), .B(n4071), .S(n3076), .Z(n3300) );
  INV_X1 U3488 ( .A(n3300), .ZN(n3657) );
  INV_X1 U3489 ( .A(n3294), .ZN(n3644) );
  AOI22_X1 U3490 ( .A1(n3604), .A2(n3657), .B1(n3644), .B2(n3601), .ZN(n3089)
         );
  INV_X1 U3491 ( .A(operand_c_i[30]), .ZN(n3296) );
  NAND2_X1 U3492 ( .A1(n3394), .A2(operand_b_i[30]), .ZN(n3077) );
  OAI211_X1 U3493 ( .C1(n3228), .C2(n3296), .A(n3219), .B(n3077), .ZN(n3291)
         );
  NAND2_X1 U3494 ( .A1(n3606), .A2(n3291), .ZN(n3082) );
  INV_X1 U3495 ( .A(n3979), .ZN(n4147) );
  NAND2_X1 U3496 ( .A1(n3079), .A2(n3078), .ZN(n3080) );
  AOI22_X1 U3497 ( .A1(n4147), .A2(operand_c_i[14]), .B1(n4146), .B2(n3080), 
        .ZN(n3081) );
  OAI211_X1 U3498 ( .C1(n3612), .C2(n4071), .A(n3082), .B(n3081), .ZN(n3083)
         );
  INV_X1 U3499 ( .A(n3083), .ZN(n3088) );
  INV_X1 U3500 ( .A(operand_c_i[22]), .ZN(n3111) );
  NAND2_X1 U3501 ( .A1(n3394), .A2(operand_b_i[22]), .ZN(n3084) );
  OAI211_X1 U3502 ( .C1(n3228), .C2(n3111), .A(n3221), .B(n3084), .ZN(n3648)
         );
  NAND2_X1 U3503 ( .A1(n3394), .A2(operand_b_i[14]), .ZN(n3085) );
  OAI211_X1 U3504 ( .C1(n3228), .C2(n3086), .A(n3227), .B(n3085), .ZN(n3646)
         );
  AOI22_X1 U3505 ( .A1(n3617), .A2(n3648), .B1(n3615), .B2(n3646), .ZN(n3087)
         );
  NAND4_X1 U3506 ( .A1(n3090), .A2(n3089), .A3(n3088), .A4(n3087), .ZN(n3091)
         );
  AOI211_X1 U3507 ( .C1(result_div[14]), .C2(n3988), .A(n3623), .B(n3091), 
        .ZN(n3098) );
  INV_X1 U3508 ( .A(n3105), .ZN(n3093) );
  OAI22_X1 U3509 ( .A1(n3093), .A2(n3990), .B1(n3092), .B2(n3989), .ZN(n3094)
         );
  OAI21_X1 U3510 ( .B1(n3626), .B2(n3094), .A(n4300), .ZN(n3097) );
  NAND2_X1 U3511 ( .A1(n3628), .A2(n3095), .ZN(n3096) );
  NAND4_X1 U3512 ( .A1(n3099), .A2(n3098), .A3(n3097), .A4(n3096), .ZN(n3100)
         );
  AOI21_X1 U3513 ( .B1(n2968), .B2(n4059), .A(n3100), .ZN(n3102) );
  AOI22_X1 U3514 ( .A1(n3750), .A2(n3217), .B1(n3216), .B2(n3944), .ZN(n3101)
         );
  OAI211_X1 U3515 ( .C1(n4121), .C2(n3104), .A(n3102), .B(n3101), .ZN(n3103)
         );
  OAI21_X1 U3516 ( .B1(n3104), .B2(n4122), .A(n4151), .ZN(n3106) );
  NAND2_X1 U3517 ( .A1(n3106), .A2(n3093), .ZN(n3107) );
  NAND2_X1 U3518 ( .A1(n3110), .A2(n3109), .ZN(result_o[14]) );
  AOI21_X1 U3521 ( .B1(n3595), .B2(n4007), .A(n4006), .ZN(n3113) );
  INV_X1 U3522 ( .A(n3113), .ZN(n3114) );
  NAND2_X1 U3523 ( .A1(n3114), .A2(n3131), .ZN(n3115) );
  INV_X1 U3524 ( .A(n3595), .ZN(n3141) );
  MUX2_X1 U3525 ( .A(n4179), .B(n3890), .S(operand_b_i[22]), .Z(n3137) );
  NAND2_X1 U3526 ( .A1(n3892), .A2(n3657), .ZN(n3118) );
  AOI22_X1 U3527 ( .A1(n3906), .A2(n3646), .B1(n3894), .B2(n3647), .ZN(n3117)
         );
  OAI211_X1 U3528 ( .C1(n3294), .C2(n3911), .A(n3118), .B(n3117), .ZN(n3129)
         );
  INV_X1 U3529 ( .A(n3291), .ZN(n3650) );
  NAND2_X1 U3530 ( .A1(n3908), .A2(n3648), .ZN(n3123) );
  INV_X1 U3531 ( .A(n4040), .ZN(n3952) );
  NAND2_X1 U3532 ( .A1(n60), .A2(n3119), .ZN(n3121) );
  AOI22_X1 U3533 ( .A1(n3952), .A2(operand_c_i[22]), .B1(n4146), .B2(n3121), 
        .ZN(n3122) );
  OAI211_X1 U3534 ( .C1(n3650), .C2(n3770), .A(n3123), .B(n3122), .ZN(n3124)
         );
  INV_X1 U3535 ( .A(n3124), .ZN(n3127) );
  INV_X1 U3536 ( .A(n3645), .ZN(n3125) );
  OR2_X1 U3537 ( .A1(n3125), .A2(n3899), .ZN(n3126) );
  OAI211_X1 U3538 ( .C1(n3901), .C2(n4071), .A(n3127), .B(n3126), .ZN(n3128)
         );
  NOR3_X1 U3539 ( .A1(n3917), .A2(n3129), .A3(n3128), .ZN(n3136) );
  OAI22_X1 U3540 ( .A1(n3131), .A2(n3990), .B1(n3130), .B2(n3989), .ZN(n3132)
         );
  OAI21_X1 U3541 ( .B1(n3921), .B2(n3132), .A(operand_a_i[22]), .ZN(n3135) );
  NAND2_X1 U3542 ( .A1(n3923), .A2(n3133), .ZN(n3134) );
  NAND4_X1 U3543 ( .A1(n3137), .A2(n3136), .A3(n3135), .A4(n3134), .ZN(n3138)
         );
  AOI21_X1 U3544 ( .B1(result_div[22]), .B2(n3988), .A(n3138), .ZN(n3140) );
  NAND2_X1 U3545 ( .A1(n222), .A2(n4059), .ZN(n3139) );
  OAI211_X1 U3546 ( .C1(n3141), .C2(n4121), .A(n3140), .B(n3139), .ZN(n3142)
         );
  INV_X1 U3547 ( .A(operand_c_i[18]), .ZN(n3155) );
  AOI22_X1 U3550 ( .A1(n4014), .A2(n3558), .B1(n3590), .B2(n3944), .ZN(n3171)
         );
  MUX2_X1 U3551 ( .A(n4179), .B(n3890), .S(n4194), .Z(n3168) );
  MUX2_X1 U3552 ( .A(n4087), .B(n2570), .S(n3393), .Z(n3322) );
  NOR2_X1 U3553 ( .A1(n3076), .A2(operand_a_i[26]), .ZN(n3146) );
  AOI21_X1 U3554 ( .B1(n3322), .B2(n3076), .A(n3146), .ZN(n3402) );
  INV_X1 U3555 ( .A(n3402), .ZN(n3323) );
  MUX2_X1 U3556 ( .A(n71), .B(n4087), .S(n3076), .Z(n3329) );
  INV_X1 U3557 ( .A(n3329), .ZN(n3405) );
  NAND2_X1 U3558 ( .A1(n3892), .A2(n3405), .ZN(n3150) );
  INV_X1 U3559 ( .A(operand_c_i[26]), .ZN(n3191) );
  NAND2_X1 U3560 ( .A1(n3394), .A2(n170), .ZN(n3147) );
  OAI211_X1 U3561 ( .C1(n3228), .C2(n3191), .A(n3219), .B(n3147), .ZN(n3403)
         );
  INV_X1 U3562 ( .A(operand_c_i[2]), .ZN(n3417) );
  NAND2_X1 U3563 ( .A1(n3394), .A2(operand_b_i[2]), .ZN(n3148) );
  OAI211_X1 U3564 ( .C1(n3228), .C2(n3417), .A(n3223), .B(n3148), .ZN(n3414)
         );
  AOI22_X1 U3565 ( .A1(n3896), .A2(n3403), .B1(n3894), .B2(n3414), .ZN(n3149)
         );
  OAI211_X1 U3566 ( .C1(n3323), .C2(n3899), .A(n3150), .B(n3149), .ZN(n3161)
         );
  NOR2_X1 U3567 ( .A1(n3901), .A2(n4087), .ZN(n3159) );
  INV_X1 U3568 ( .A(operand_c_i[10]), .ZN(n3325) );
  NAND2_X1 U3569 ( .A1(n3394), .A2(operand_b_i[10]), .ZN(n3151) );
  OAI211_X1 U3570 ( .C1(n3228), .C2(n3325), .A(n3227), .B(n3151), .ZN(n3413)
         );
  OAI22_X1 U3571 ( .A1(n4040), .A2(n3155), .B1(n4038), .B2(n3152), .ZN(n3153)
         );
  AOI21_X1 U3572 ( .B1(n3906), .B2(n3413), .A(n3153), .ZN(n3157) );
  NAND2_X1 U3573 ( .A1(n3394), .A2(n4194), .ZN(n3154) );
  OAI211_X1 U3574 ( .C1(n3228), .C2(n3155), .A(n3221), .B(n3154), .ZN(n3406)
         );
  NAND2_X1 U3575 ( .A1(n3908), .A2(n3406), .ZN(n3156) );
  OAI211_X1 U3576 ( .C1(n3322), .C2(n3911), .A(n3157), .B(n3156), .ZN(n3158)
         );
  OR2_X1 U3577 ( .A1(n3159), .A2(n3158), .ZN(n3160) );
  NOR3_X1 U3578 ( .A1(n3917), .A2(n3161), .A3(n3160), .ZN(n3167) );
  NAND2_X1 U3579 ( .A1(n3174), .A2(n4126), .ZN(n3162) );
  OAI21_X1 U3580 ( .B1(n4021), .B2(n3163), .A(n3162), .ZN(n3164) );
  OAI21_X1 U3581 ( .B1(n3921), .B2(n3164), .A(n72), .ZN(n3166) );
  NAND2_X1 U3582 ( .A1(n3923), .A2(n1043), .ZN(n3165) );
  NAND4_X1 U3583 ( .A1(n3168), .A2(n3167), .A3(n3166), .A4(n3165), .ZN(n3169)
         );
  AOI21_X1 U3584 ( .B1(result_div[18]), .B2(n3988), .A(n3169), .ZN(n3170) );
  OAI211_X1 U3585 ( .C1(n3144), .C2(n4184), .A(n3170), .B(n3171), .ZN(n3172)
         );
  INV_X1 U3586 ( .A(n3172), .ZN(n3181) );
  INV_X1 U3587 ( .A(n3558), .ZN(n3173) );
  OAI21_X1 U3588 ( .B1(n3173), .B2(n4122), .A(n4151), .ZN(n3176) );
  INV_X1 U3589 ( .A(n3174), .ZN(n3175) );
  NAND2_X1 U3590 ( .A1(n3176), .A2(n3175), .ZN(n3179) );
  INV_X1 U3591 ( .A(n4309), .ZN(n3178) );
  INV_X1 U3595 ( .A(n3206), .ZN(n3212) );
  MUX2_X1 U3596 ( .A(n4017), .B(n4016), .S(n170), .Z(n3202) );
  NAND2_X1 U3597 ( .A1(n3206), .A2(n4126), .ZN(n3185) );
  OAI21_X1 U3598 ( .B1(n4021), .B2(n3186), .A(n3185), .ZN(n3187) );
  OAI21_X1 U3599 ( .B1(n4023), .B2(n3187), .A(operand_a_i[26]), .ZN(n3200) );
  AOI22_X1 U3600 ( .A1(n4027), .A2(n3402), .B1(n4025), .B2(n3414), .ZN(n3189)
         );
  AOI22_X1 U3601 ( .A1(n4031), .A2(n3403), .B1(n4029), .B2(n3413), .ZN(n3188)
         );
  OAI211_X1 U3602 ( .C1(n3322), .C2(n4034), .A(n3189), .B(n3188), .ZN(n3196)
         );
  INV_X1 U3603 ( .A(n4045), .ZN(n3866) );
  NAND2_X1 U3604 ( .A1(n4036), .A2(operand_a_i[2]), .ZN(n3194) );
  OAI22_X1 U3605 ( .A1(n4040), .A2(n3191), .B1(n4038), .B2(n3190), .ZN(n3192)
         );
  AOI21_X1 U3606 ( .B1(n4043), .B2(n3406), .A(n3192), .ZN(n3193) );
  OAI211_X1 U3607 ( .C1(n3329), .C2(n3866), .A(n3194), .B(n3193), .ZN(n3195)
         );
  NOR2_X1 U3608 ( .A1(n3196), .A2(n3195), .ZN(n3199) );
  NAND2_X1 U3609 ( .A1(n4052), .A2(n3197), .ZN(n3198) );
  NAND4_X1 U3610 ( .A1(n3200), .A2(n3199), .A3(n3198), .A4(n4054), .ZN(n3201)
         );
  AOI211_X1 U3611 ( .C1(result_div[26]), .C2(n3988), .A(n3202), .B(n3201), 
        .ZN(n3204) );
  NAND2_X1 U3612 ( .A1(n4305), .A2(n3750), .ZN(n3203) );
  OAI211_X1 U3613 ( .C1(n3793), .C2(n4192), .A(n3204), .B(n3203), .ZN(n3205)
         );
  AOI21_X1 U3614 ( .B1(n4014), .B2(n3794), .A(n3205), .ZN(n3210) );
  AOI21_X1 U3615 ( .B1(n3794), .B2(n4007), .A(n4006), .ZN(n3207) );
  INV_X1 U3616 ( .A(operand_c_i[12]), .ZN(n3230) );
  INV_X1 U3618 ( .A(n3251), .ZN(n3214) );
  INV_X1 U3620 ( .A(n3216), .ZN(n3250) );
  AOI22_X1 U3621 ( .A1(n3944), .A2(n3217), .B1(n4309), .B2(n4014), .ZN(n3249)
         );
  MUX2_X1 U3622 ( .A(n4179), .B(n3596), .S(operand_b_i[12]), .Z(n3246) );
  INV_X1 U3623 ( .A(operand_c_i[28]), .ZN(n3861) );
  NAND2_X1 U3624 ( .A1(n3394), .A2(operand_b_i[28]), .ZN(n3218) );
  OAI211_X1 U3625 ( .C1(n3228), .C2(n3861), .A(n3219), .B(n3218), .ZN(n3895)
         );
  INV_X1 U3626 ( .A(operand_c_i[20]), .ZN(n3903) );
  NAND2_X1 U3627 ( .A1(n3394), .A2(operand_b_i[20]), .ZN(n3220) );
  OAI211_X1 U3628 ( .C1(n3228), .C2(n3903), .A(n3221), .B(n3220), .ZN(n3907)
         );
  AOI22_X1 U3629 ( .A1(n3606), .A2(n3895), .B1(n3617), .B2(n3907), .ZN(n3238)
         );
  MUX2_X1 U3630 ( .A(n4108), .B(n2561), .S(n3393), .Z(n3912) );
  INV_X1 U3631 ( .A(n3912), .ZN(n3803) );
  INV_X1 U3632 ( .A(operand_c_i[4]), .ZN(n3799) );
  NAND2_X1 U3633 ( .A1(n3394), .A2(operand_b_i[4]), .ZN(n3222) );
  OAI211_X1 U3634 ( .C1(n3228), .C2(n3799), .A(n3223), .B(n3222), .ZN(n3893)
         );
  AOI22_X1 U3635 ( .A1(n3803), .A2(n3601), .B1(n3598), .B2(n3893), .ZN(n3237)
         );
  OR2_X1 U3636 ( .A1(n3076), .A2(n2522), .ZN(n3224) );
  OAI21_X1 U3637 ( .B1(n3912), .B2(n3225), .A(n3224), .ZN(n3857) );
  INV_X1 U3638 ( .A(n3857), .ZN(n3900) );
  OAI22_X1 U3639 ( .A1(n3900), .A2(n3562), .B1(n3612), .B2(n4108), .ZN(n3235)
         );
  MUX2_X1 U3640 ( .A(n4067), .B(n4108), .S(n3076), .Z(n3865) );
  NAND2_X1 U3641 ( .A1(n3394), .A2(operand_b_i[12]), .ZN(n3226) );
  OAI211_X1 U3642 ( .C1(n3228), .C2(n3230), .A(n3227), .B(n3226), .ZN(n3905)
         );
  NAND2_X1 U3643 ( .A1(n3615), .A2(n3905), .ZN(n3233) );
  OAI22_X1 U3644 ( .A1(n3979), .A2(n3230), .B1(n4038), .B2(n3229), .ZN(n3231)
         );
  INV_X1 U3645 ( .A(n3231), .ZN(n3232) );
  OAI211_X1 U3646 ( .C1(n3570), .C2(n3865), .A(n3233), .B(n3232), .ZN(n3234)
         );
  NOR2_X1 U3647 ( .A1(n3235), .A2(n3234), .ZN(n3236) );
  NAND4_X1 U3648 ( .A1(n3576), .A2(n3238), .A3(n3237), .A4(n3236), .ZN(n3239)
         );
  AOI21_X1 U3649 ( .B1(result_div[12]), .B2(n3988), .A(n3239), .ZN(n3245) );
  OAI22_X1 U3650 ( .A1(n3251), .A2(n3990), .B1(n3240), .B2(n4021), .ZN(n3241)
         );
  OAI21_X1 U3651 ( .B1(n3626), .B2(n3241), .A(n163), .ZN(n3244) );
  NAND2_X1 U3652 ( .A1(n3628), .A2(n3242), .ZN(n3243) );
  NAND4_X1 U3653 ( .A1(n3246), .A2(n3245), .A3(n3244), .A4(n3243), .ZN(n3247)
         );
  AOI21_X1 U3654 ( .B1(n3558), .B2(n4059), .A(n3247), .ZN(n3248) );
  OAI211_X1 U3655 ( .C1(n3250), .C2(n4184), .A(n3249), .B(n3248), .ZN(n3254)
         );
  OAI21_X1 U3656 ( .B1(n3178), .B2(n4122), .A(n4151), .ZN(n3252) );
  NAND2_X1 U3657 ( .A1(n3256), .A2(n3255), .ZN(result_o[12]) );
  INV_X1 U3658 ( .A(n3320), .ZN(n3636) );
  OAI21_X1 U3659 ( .B1(n3636), .B2(n4122), .A(n4151), .ZN(n3258) );
  MUX2_X1 U3661 ( .A(n4179), .B(n3890), .S(operand_b_i[21]), .Z(n3278) );
  INV_X1 U3662 ( .A(n3732), .ZN(n3563) );
  NAND2_X1 U3663 ( .A1(n3892), .A2(n3731), .ZN(n3260) );
  AOI22_X1 U3664 ( .A1(n3896), .A2(n3560), .B1(n3894), .B2(n3726), .ZN(n3259)
         );
  OAI211_X1 U3665 ( .C1(n3563), .C2(n3899), .A(n3260), .B(n3259), .ZN(n3269)
         );
  NOR2_X1 U3666 ( .A1(n3901), .A2(n4079), .ZN(n3267) );
  OAI22_X1 U3667 ( .A1(n4040), .A2(n3262), .B1(n4038), .B2(n3261), .ZN(n3263)
         );
  AOI21_X1 U3668 ( .B1(n3906), .B2(n3725), .A(n3263), .ZN(n3265) );
  NAND2_X1 U3669 ( .A1(n3908), .A2(n3559), .ZN(n3264) );
  OAI211_X1 U3670 ( .C1(n3561), .C2(n3911), .A(n3265), .B(n3264), .ZN(n3266)
         );
  OR2_X1 U3671 ( .A1(n3267), .A2(n3266), .ZN(n3268) );
  NOR3_X1 U3672 ( .A1(n3917), .A2(n3269), .A3(n3268), .ZN(n3277) );
  NAND2_X1 U3673 ( .A1(n3270), .A2(n4126), .ZN(n3272) );
  NAND2_X1 U3674 ( .A1(n4125), .A2(operand_b_i[21]), .ZN(n3271) );
  NAND2_X1 U3675 ( .A1(n3272), .A2(n3271), .ZN(n3273) );
  OAI21_X1 U3676 ( .B1(n3921), .B2(n3273), .A(operand_a_i[21]), .ZN(n3276) );
  NAND2_X1 U3677 ( .A1(n3923), .A2(n3274), .ZN(n3275) );
  NAND4_X1 U3678 ( .A1(n3278), .A2(n3277), .A3(n3276), .A4(n3275), .ZN(n3279)
         );
  AOI21_X1 U3679 ( .B1(result_div[21]), .B2(n3988), .A(n3279), .ZN(n3282) );
  NAND2_X1 U3680 ( .A1(n222), .A2(n3750), .ZN(n3281) );
  OAI211_X1 U3681 ( .C1(n3144), .C2(n4192), .A(n3282), .B(n3281), .ZN(n3283)
         );
  INV_X1 U3682 ( .A(n3283), .ZN(n3286) );
  INV_X1 U3683 ( .A(n125), .ZN(n3346) );
  OAI22_X1 U3684 ( .A1(n3346), .A2(n4182), .B1(n3636), .B2(n4121), .ZN(n3284)
         );
  INV_X1 U3685 ( .A(n3284), .ZN(n3285) );
  AND2_X1 U3688 ( .A1(n4316), .A2(n4059), .ZN(n3309) );
  MUX2_X1 U3689 ( .A(n4017), .B(n4016), .S(operand_b_i[30]), .Z(n3307) );
  INV_X1 U3690 ( .A(n4023), .ZN(n3289) );
  AOI22_X1 U3691 ( .A1(n3313), .A2(n4126), .B1(operand_b_i[30]), .B2(n4125), 
        .ZN(n3288) );
  AOI21_X1 U3692 ( .B1(n3289), .B2(n3288), .A(n4112), .ZN(n3306) );
  NAND2_X1 U3693 ( .A1(n4052), .A2(n3290), .ZN(n3304) );
  AOI22_X1 U3694 ( .A1(n4027), .A2(n3645), .B1(n4025), .B2(n3647), .ZN(n3293)
         );
  AOI22_X1 U3695 ( .A1(n4031), .A2(n3291), .B1(n4029), .B2(n3646), .ZN(n3292)
         );
  OAI211_X1 U3696 ( .C1(n4034), .C2(n3294), .A(n3293), .B(n3292), .ZN(n3302)
         );
  NAND2_X1 U3697 ( .A1(n4036), .A2(operand_a_i[6]), .ZN(n3299) );
  OAI22_X1 U3698 ( .A1(n4040), .A2(n3296), .B1(n4038), .B2(n3295), .ZN(n3297)
         );
  AOI21_X1 U3699 ( .B1(n4043), .B2(n3648), .A(n3297), .ZN(n3298) );
  OAI211_X1 U3700 ( .C1(n3866), .C2(n3300), .A(n3299), .B(n3298), .ZN(n3301)
         );
  NOR2_X1 U3701 ( .A1(n3302), .A2(n3301), .ZN(n3303) );
  NAND3_X1 U3702 ( .A1(n3304), .A2(n3303), .A3(n4054), .ZN(n3305) );
  OR3_X1 U3703 ( .A1(n3307), .A2(n3306), .A3(n3305), .ZN(n3308) );
  AOI211_X1 U3704 ( .C1(result_div[30]), .C2(n3988), .A(n3309), .B(n3308), 
        .ZN(n3311) );
  NAND2_X1 U3705 ( .A1(n3711), .A2(n3944), .ZN(n3310) );
  OAI211_X1 U3706 ( .C1(n4121), .C2(n4193), .A(n3311), .B(n3310), .ZN(n3312)
         );
  OAI21_X1 U3707 ( .B1(n4193), .B2(n4122), .A(n4151), .ZN(n3315) );
  NAND2_X1 U3708 ( .A1(n3315), .A2(n3314), .ZN(n3316) );
  AOI22_X1 U3711 ( .A1(n4012), .A2(n4311), .B1(n125), .B2(n4014), .ZN(n3345)
         );
  MUX2_X1 U3712 ( .A(n4179), .B(n3596), .S(operand_b_i[10]), .Z(n3342) );
  NAND2_X1 U3713 ( .A1(result_div[10]), .A2(n3988), .ZN(n3335) );
  AOI22_X1 U3714 ( .A1(n3606), .A2(n3403), .B1(n3617), .B2(n3406), .ZN(n3334)
         );
  INV_X1 U3715 ( .A(n3322), .ZN(n3422) );
  AOI22_X1 U3716 ( .A1(n3422), .A2(n3601), .B1(n3598), .B2(n3414), .ZN(n3333)
         );
  OAI22_X1 U3717 ( .A1(n3323), .A2(n3562), .B1(n3612), .B2(n4087), .ZN(n3331)
         );
  NAND2_X1 U3718 ( .A1(n3615), .A2(n3413), .ZN(n3328) );
  OAI22_X1 U3719 ( .A1(n3979), .A2(n3325), .B1(n4038), .B2(n3324), .ZN(n3326)
         );
  INV_X1 U3720 ( .A(n3326), .ZN(n3327) );
  OAI211_X1 U3721 ( .C1(n3570), .C2(n3329), .A(n3328), .B(n3327), .ZN(n3330)
         );
  NOR2_X1 U3722 ( .A1(n3331), .A2(n3330), .ZN(n3332) );
  NAND4_X1 U3723 ( .A1(n3335), .A2(n3334), .A3(n3333), .A4(n3332), .ZN(n3336)
         );
  AOI211_X1 U3724 ( .C1(n3628), .C2(n3337), .A(n3623), .B(n3336), .ZN(n3341)
         );
  INV_X1 U3725 ( .A(n3347), .ZN(n3338) );
  OAI22_X1 U3726 ( .A1(n3338), .A2(n3990), .B1(n2571), .B2(n3989), .ZN(n3339)
         );
  OAI21_X1 U3727 ( .B1(n3626), .B2(n3339), .A(n167), .ZN(n3340) );
  NAND3_X1 U3728 ( .A1(n3342), .A2(n3341), .A3(n3340), .ZN(n3343) );
  AOI21_X1 U3729 ( .B1(n3321), .B2(n4059), .A(n3343), .ZN(n3344) );
  OAI21_X1 U3730 ( .B1(n3346), .B2(n4122), .A(n4151), .ZN(n3348) );
  NAND2_X1 U3731 ( .A1(n3348), .A2(n3338), .ZN(n3349) );
  INV_X1 U3732 ( .A(n3852), .ZN(n3849) );
  NAND2_X1 U3733 ( .A1(n4123), .A2(n3750), .ZN(n3450) );
  INV_X1 U3734 ( .A(n3740), .ZN(n3354) );
  NOR2_X1 U3735 ( .A1(n3354), .A2(n3351), .ZN(n3796) );
  MUX2_X1 U3736 ( .A(n4161), .B(n3882), .S(ff1_result[2]), .Z(n3352) );
  AOI21_X1 U3737 ( .B1(n3353), .B2(n3796), .A(n3352), .ZN(n3442) );
  NOR2_X1 U3738 ( .A1(ff_no_one), .A2(n3354), .ZN(n3700) );
  INV_X1 U3739 ( .A(n3700), .ZN(n4172) );
  AND2_X1 U3740 ( .A1(n3355), .A2(n3387), .ZN(n3356) );
  NOR2_X1 U3741 ( .A1(n3357), .A2(n3356), .ZN(n3371) );
  MUX2_X1 U3742 ( .A(n3359), .B(n3358), .S(n3371), .Z(n3444) );
  NOR2_X1 U3743 ( .A1(n3360), .A2(n3444), .ZN(n4177) );
  AND2_X1 U3744 ( .A1(n3796), .A2(n4304), .ZN(n3379) );
  NOR2_X1 U3745 ( .A1(n3373), .A2(n3361), .ZN(n3367) );
  NAND3_X1 U3746 ( .A1(n2638), .A2(n3363), .A3(n3362), .ZN(n3365) );
  NAND2_X1 U3747 ( .A1(n3365), .A2(n3364), .ZN(n3366) );
  MUX2_X1 U3748 ( .A(n3368), .B(n3367), .S(n3366), .Z(n3369) );
  NAND3_X1 U3749 ( .A1(n3371), .A2(n3370), .A3(n3369), .ZN(n3378) );
  INV_X1 U3750 ( .A(n3371), .ZN(n3376) );
  NOR2_X1 U3751 ( .A1(n3373), .A2(n3372), .ZN(n3375) );
  AOI21_X1 U3752 ( .B1(n3376), .B2(n3375), .A(n3374), .ZN(n3377) );
  AND2_X1 U3753 ( .A1(n3378), .A2(n3377), .ZN(n3986) );
  AOI21_X1 U3754 ( .B1(ff_no_one), .B2(n3379), .A(n3986), .ZN(n4171) );
  NOR2_X1 U3755 ( .A1(n498), .A2(n3380), .ZN(n3381) );
  AND2_X1 U3756 ( .A1(n3835), .A2(n3381), .ZN(n4169) );
  AND2_X1 U3757 ( .A1(n3382), .A2(operand_b_i[1]), .ZN(n3383) );
  OR2_X1 U3758 ( .A1(n3384), .A2(n3383), .ZN(n3411) );
  NOR2_X1 U3759 ( .A1(n3386), .A2(n3385), .ZN(n3388) );
  OAI21_X1 U3760 ( .B1(n3389), .B2(n3388), .A(n3387), .ZN(n3410) );
  INV_X1 U3761 ( .A(n3410), .ZN(n3390) );
  NAND2_X1 U3762 ( .A1(n3411), .A2(n3390), .ZN(n3401) );
  OR2_X1 U3763 ( .A1(n3391), .A2(operand_b_i[2]), .ZN(n3400) );
  INV_X1 U3764 ( .A(imm_vec_ext_i[1]), .ZN(n3392) );
  OR2_X1 U3765 ( .A1(n3393), .A2(n3392), .ZN(n3399) );
  AOI22_X1 U3766 ( .A1(n3396), .A2(n3395), .B1(n3394), .B2(n4131), .ZN(n3397)
         );
  NAND4_X1 U3767 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3431)
         );
  INV_X1 U3768 ( .A(n3431), .ZN(n3412) );
  OR2_X1 U3769 ( .A1(n3401), .A2(n3412), .ZN(n3722) );
  INV_X1 U3770 ( .A(n3722), .ZN(n4136) );
  NOR2_X1 U3771 ( .A1(n3401), .A2(n3431), .ZN(n4133) );
  AOI22_X1 U3772 ( .A1(n4136), .A2(n3403), .B1(n4133), .B2(n3402), .ZN(n3426)
         );
  NAND2_X1 U3773 ( .A1(n3411), .A2(n3410), .ZN(n3404) );
  OR2_X1 U3774 ( .A1(n3404), .A2(n3412), .ZN(n3721) );
  INV_X1 U3775 ( .A(n3721), .ZN(n4154) );
  NOR2_X1 U3776 ( .A1(n3404), .A2(n3431), .ZN(n4144) );
  AOI22_X1 U3777 ( .A1(n4154), .A2(n3406), .B1(n4144), .B2(n3405), .ZN(n3425)
         );
  NAND2_X1 U3778 ( .A1(n3410), .A2(n3407), .ZN(n3408) );
  NOR2_X1 U3779 ( .A1(n3411), .A2(n3408), .ZN(n3434) );
  INV_X1 U3780 ( .A(n3434), .ZN(n3409) );
  NOR2_X1 U3781 ( .A1(n3409), .A2(n3412), .ZN(n4142) );
  OR2_X1 U3782 ( .A1(n3411), .A2(n3410), .ZN(n3415) );
  NOR2_X1 U3783 ( .A1(n3415), .A2(n3412), .ZN(n4138) );
  AOI22_X1 U3784 ( .A1(n4142), .A2(n3414), .B1(n4138), .B2(n3413), .ZN(n3424)
         );
  NOR2_X1 U3785 ( .A1(n3415), .A2(n3431), .ZN(n4139) );
  NAND2_X1 U3786 ( .A1(result_div[2]), .A2(n3988), .ZN(n3420) );
  OAI22_X1 U3787 ( .A1(n3979), .A2(n3417), .B1(n4038), .B2(n3416), .ZN(n3418)
         );
  INV_X1 U3788 ( .A(n3418), .ZN(n3419) );
  NAND2_X1 U3789 ( .A1(n3420), .A2(n3419), .ZN(n3421) );
  AOI21_X1 U3790 ( .B1(n4139), .B2(n3422), .A(n3421), .ZN(n3423) );
  NAND4_X1 U3791 ( .A1(n3426), .A2(n3425), .A3(n3424), .A4(n3423), .ZN(n3427)
         );
  AOI21_X1 U3792 ( .B1(cnt_result[2]), .B2(n4169), .A(n3427), .ZN(n3428) );
  NAND2_X1 U3793 ( .A1(n4171), .A2(n3428), .ZN(n3429) );
  AOI21_X1 U3794 ( .B1(n4177), .B2(n3430), .A(n3429), .ZN(n3441) );
  INV_X1 U3795 ( .A(n3444), .ZN(n3436) );
  NOR2_X1 U3796 ( .A1(n3431), .A2(n4147), .ZN(n3433) );
  AOI21_X1 U3797 ( .B1(n3434), .B2(n3433), .A(n3432), .ZN(n3435) );
  OAI21_X1 U3798 ( .B1(n3437), .B2(n3436), .A(n3435), .ZN(n4124) );
  OAI22_X1 U3799 ( .A1(n3456), .A2(n3990), .B1(n3438), .B2(n3989), .ZN(n3439)
         );
  OAI21_X1 U3800 ( .B1(n4124), .B2(n3439), .A(operand_a_i[2]), .ZN(n3440) );
  OAI211_X1 U3801 ( .C1(n3442), .C2(n4172), .A(n3441), .B(n3440), .ZN(n3448)
         );
  NAND2_X1 U3802 ( .A1(n3444), .A2(n3443), .ZN(n3445) );
  AND2_X1 U3803 ( .A1(n3446), .A2(n3445), .ZN(n3718) );
  MUX2_X1 U3804 ( .A(n4017), .B(n3718), .S(operand_b_i[2]), .Z(n3447) );
  NOR2_X1 U3805 ( .A1(n3448), .A2(n3447), .ZN(n3449) );
  NAND2_X1 U3806 ( .A1(n3450), .A2(n3449), .ZN(n3451) );
  AOI21_X1 U3807 ( .B1(n3875), .B2(n4014), .A(n3451), .ZN(n3453) );
  NAND2_X1 U3808 ( .A1(n3463), .A2(n3944), .ZN(n3452) );
  OAI211_X1 U3809 ( .C1(n3849), .C2(n4192), .A(n3453), .B(n3452), .ZN(n3454)
         );
  NAND2_X1 U3810 ( .A1(n3875), .A2(n4007), .ZN(n3455) );
  NAND2_X1 U3811 ( .A1(n3455), .A2(n4151), .ZN(n3457) );
  NAND2_X1 U3812 ( .A1(n3457), .A2(n3456), .ZN(n3458) );
  INV_X1 U3813 ( .A(n3463), .ZN(n4185) );
  INV_X1 U3814 ( .A(n3796), .ZN(n3685) );
  MUX2_X1 U3816 ( .A(n3683), .B(n4116), .S(ff1_result[3]), .Z(n3465) );
  OAI21_X1 U3817 ( .B1(n3464), .B2(n3685), .A(n3465), .ZN(n3487) );
  MUX2_X1 U3818 ( .A(n4017), .B(n3718), .S(operand_b_i[3]), .Z(n3486) );
  INV_X1 U3819 ( .A(n4177), .ZN(n3484) );
  INV_X1 U3820 ( .A(n3466), .ZN(n3483) );
  OAI22_X1 U3821 ( .A1(n3979), .A2(n3468), .B1(n4038), .B2(n3467), .ZN(n3471)
         );
  INV_X1 U3822 ( .A(n3605), .ZN(n3469) );
  NOR2_X1 U3823 ( .A1(n3722), .A2(n3469), .ZN(n3470) );
  AOI211_X1 U3824 ( .C1(n3988), .C2(result_div[3]), .A(n3471), .B(n3470), .ZN(
        n3476) );
  AOI22_X1 U3825 ( .A1(n3602), .A2(n4139), .B1(n4138), .B2(n3614), .ZN(n3475)
         );
  INV_X1 U3826 ( .A(n3472), .ZN(n3599) );
  AOI22_X1 U3827 ( .A1(n4133), .A2(n3599), .B1(n4144), .B2(n3603), .ZN(n3474)
         );
  AOI22_X1 U3828 ( .A1(n4154), .A2(n3616), .B1(n4142), .B2(n3597), .ZN(n3473)
         );
  NAND4_X1 U3829 ( .A1(n3476), .A2(n3475), .A3(n3474), .A4(n3473), .ZN(n3478)
         );
  INV_X1 U3830 ( .A(n4171), .ZN(n3477) );
  AOI211_X1 U3831 ( .C1(cnt_result[3]), .C2(n4169), .A(n3478), .B(n3477), .ZN(
        n3482) );
  OAI22_X1 U3832 ( .A1(n3491), .A2(n3990), .B1(n3479), .B2(n3989), .ZN(n3480)
         );
  OAI21_X1 U3833 ( .B1(n4124), .B2(n3480), .A(n48), .ZN(n3481) );
  OAI211_X1 U3834 ( .C1(n3484), .C2(n3483), .A(n3482), .B(n3481), .ZN(n3485)
         );
  AOI211_X1 U3835 ( .C1(n3487), .C2(n3700), .A(n3486), .B(n3485), .ZN(n3488)
         );
  OAI21_X1 U3836 ( .B1(n4185), .B2(n4192), .A(n3488), .ZN(n3489) );
  AOI21_X1 U3837 ( .B1(n4014), .B2(n3853), .A(n3489), .ZN(n3494) );
  OAI21_X1 U3838 ( .B1(n3490), .B2(n4122), .A(n4151), .ZN(n3492) );
  AOI22_X1 U3839 ( .A1(n3492), .A2(n3491), .B1(n3750), .B2(n3794), .ZN(n3493)
         );
  OAI211_X1 U3840 ( .C1(n3849), .C2(n4182), .A(n3494), .B(n3493), .ZN(n3495)
         );
  NAND2_X1 U3841 ( .A1(n3497), .A2(n3496), .ZN(result_o[3]) );
  NAND2_X1 U3842 ( .A1(n3498), .A2(n1007), .ZN(n3528) );
  AOI22_X1 U3843 ( .A1(n3750), .A2(n3321), .B1(n3595), .B2(n3944), .ZN(n3520)
         );
  MUX2_X1 U3844 ( .A(n4179), .B(n3596), .S(n4195), .Z(n3516) );
  NAND2_X1 U3845 ( .A1(result_div[9]), .A2(n3988), .ZN(n3510) );
  AOI22_X1 U3846 ( .A1(n3617), .A2(n4042), .B1(n3606), .B2(n4030), .ZN(n3509)
         );
  AOI22_X1 U3847 ( .A1(n3687), .A2(n3601), .B1(n3598), .B2(n4024), .ZN(n3508)
         );
  OAI22_X1 U3848 ( .A1(n3688), .A2(n3562), .B1(n3612), .B2(n2546), .ZN(n3506)
         );
  INV_X1 U3849 ( .A(n4044), .ZN(n3504) );
  NAND2_X1 U3850 ( .A1(n3615), .A2(n4028), .ZN(n3503) );
  OAI22_X1 U3851 ( .A1(n3979), .A2(n3500), .B1(n4038), .B2(n3499), .ZN(n3501)
         );
  INV_X1 U3852 ( .A(n3501), .ZN(n3502) );
  OAI211_X1 U3853 ( .C1(n3570), .C2(n3504), .A(n3503), .B(n3502), .ZN(n3505)
         );
  NOR2_X1 U3854 ( .A1(n3506), .A2(n3505), .ZN(n3507) );
  NAND4_X1 U3855 ( .A1(n3510), .A2(n3509), .A3(n3508), .A4(n3507), .ZN(n3511)
         );
  AOI211_X1 U3856 ( .C1(n3628), .C2(n3512), .A(n3623), .B(n3511), .ZN(n3515)
         );
  OAI22_X1 U3857 ( .A1(n3523), .A2(n3990), .B1(n2567), .B2(n3989), .ZN(n3513)
         );
  OAI21_X1 U3858 ( .B1(n3626), .B2(n3513), .A(operand_a_i[9]), .ZN(n3514) );
  NAND3_X1 U3859 ( .A1(n3516), .A2(n3515), .A3(n3514), .ZN(n3517) );
  AOI21_X1 U3860 ( .B1(n4365), .B2(n4059), .A(n3517), .ZN(n3519) );
  NAND2_X1 U3861 ( .A1(n3521), .A2(n4014), .ZN(n3518) );
  NAND3_X1 U3862 ( .A1(n3520), .A2(n3519), .A3(n3518), .ZN(n3526) );
  AOI21_X1 U3863 ( .B1(n3521), .B2(n4007), .A(n4006), .ZN(n3522) );
  INV_X1 U3864 ( .A(n3522), .ZN(n3524) );
  NAND2_X1 U3865 ( .A1(n3528), .A2(n3527), .ZN(result_o[9]) );
  INV_X1 U3867 ( .A(n4305), .ZN(n4000) );
  MUX2_X1 U3868 ( .A(n4017), .B(n4016), .S(n4340), .Z(n3547) );
  INV_X1 U3869 ( .A(n3552), .ZN(n3531) );
  OAI22_X1 U3870 ( .A1(n3531), .A2(n3990), .B1(n3530), .B2(n3989), .ZN(n3532)
         );
  OAI21_X1 U3871 ( .B1(n4023), .B2(n3532), .A(operand_a_i[24]), .ZN(n3545) );
  OAI22_X1 U3872 ( .A1(n4040), .A2(n3534), .B1(n4038), .B2(n3533), .ZN(n3535)
         );
  AOI21_X1 U3873 ( .B1(n4043), .B2(n4153), .A(n3535), .ZN(n3536) );
  OAI21_X1 U3874 ( .B1(n3537), .B2(n4132), .A(n3536), .ZN(n3541) );
  AOI22_X1 U3875 ( .A1(n4045), .A2(n4143), .B1(n4029), .B2(n4137), .ZN(n3539)
         );
  AOI22_X1 U3876 ( .A1(n4031), .A2(n4135), .B1(n4025), .B2(n4141), .ZN(n3538)
         );
  OAI211_X1 U3877 ( .C1(n4034), .C2(n3771), .A(n3539), .B(n3538), .ZN(n3540)
         );
  AOI211_X1 U3878 ( .C1(n4198), .C2(n4036), .A(n3541), .B(n3540), .ZN(n3544)
         );
  NAND2_X1 U3879 ( .A1(n4052), .A2(n3542), .ZN(n3543) );
  NAND4_X1 U3880 ( .A1(n3545), .A2(n3544), .A3(n4054), .A4(n3543), .ZN(n3546)
         );
  AOI211_X1 U3881 ( .C1(result_div[24]), .C2(n3988), .A(n3547), .B(n3546), 
        .ZN(n3549) );
  NAND2_X1 U3882 ( .A1(n3999), .A2(n4014), .ZN(n3548) );
  OAI211_X1 U3883 ( .C1(n4000), .C2(n4182), .A(n3549), .B(n3548), .ZN(n3550)
         );
  AOI21_X1 U3884 ( .B1(n4059), .B2(n4279), .A(n3550), .ZN(n3555) );
  AOI21_X1 U3885 ( .B1(n3999), .B2(n4007), .A(n4006), .ZN(n3551) );
  NAND2_X1 U3886 ( .A1(n3558), .A2(n4012), .ZN(n3588) );
  MUX2_X1 U3887 ( .A(n4179), .B(n3596), .S(operand_b_i[13]), .Z(n3585) );
  AOI22_X1 U3888 ( .A1(n3606), .A2(n3560), .B1(n3617), .B2(n3559), .ZN(n3575)
         );
  INV_X1 U3889 ( .A(n3561), .ZN(n3730) );
  AOI22_X1 U3890 ( .A1(n3730), .A2(n3601), .B1(n3598), .B2(n3726), .ZN(n3574)
         );
  OAI22_X1 U3891 ( .A1(n3563), .A2(n3562), .B1(n3612), .B2(n4079), .ZN(n3572)
         );
  INV_X1 U3892 ( .A(n3731), .ZN(n3569) );
  NAND2_X1 U3893 ( .A1(n3615), .A2(n3725), .ZN(n3568) );
  OAI22_X1 U3894 ( .A1(n3979), .A2(n3565), .B1(n4038), .B2(n3564), .ZN(n3566)
         );
  INV_X1 U3895 ( .A(n3566), .ZN(n3567) );
  OAI211_X1 U3896 ( .C1(n3570), .C2(n3569), .A(n3568), .B(n3567), .ZN(n3571)
         );
  NOR2_X1 U3897 ( .A1(n3572), .A2(n3571), .ZN(n3573) );
  NAND4_X1 U3898 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3577)
         );
  AOI21_X1 U3899 ( .B1(result_div[13]), .B2(n3988), .A(n3577), .ZN(n3584) );
  INV_X1 U3900 ( .A(n3591), .ZN(n3579) );
  OAI22_X1 U3901 ( .A1(n3579), .A2(n3990), .B1(n3578), .B2(n4021), .ZN(n3580)
         );
  OAI21_X1 U3902 ( .B1(n3626), .B2(n3580), .A(operand_a_i[13]), .ZN(n3583) );
  NAND2_X1 U3903 ( .A1(n3628), .A2(n3581), .ZN(n3582) );
  NAND4_X1 U3904 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3586)
         );
  AOI21_X1 U3905 ( .B1(n3590), .B2(n4014), .A(n3586), .ZN(n3587) );
  OAI211_X1 U3906 ( .C1(n3008), .C2(n4192), .A(n3588), .B(n3587), .ZN(n3589)
         );
  INV_X1 U3907 ( .A(n3590), .ZN(n3934) );
  OAI21_X1 U3908 ( .B1(n3934), .B2(n4122), .A(n4151), .ZN(n3592) );
  NAND2_X1 U3909 ( .A1(n3592), .A2(n3579), .ZN(n3593) );
  AOI22_X1 U3910 ( .A1(n3944), .A2(n3321), .B1(n3595), .B2(n3750), .ZN(n3635)
         );
  MUX2_X1 U3911 ( .A(n4179), .B(n3596), .S(n150), .Z(n3632) );
  AOI22_X1 U3912 ( .A1(n3600), .A2(n3599), .B1(n3598), .B2(n3597), .ZN(n3621)
         );
  AOI22_X1 U3913 ( .A1(n3604), .A2(n3603), .B1(n3602), .B2(n3601), .ZN(n3620)
         );
  NAND2_X1 U3914 ( .A1(n3606), .A2(n3605), .ZN(n3611) );
  OAI22_X1 U3915 ( .A1(n3979), .A2(n3608), .B1(n4038), .B2(n3607), .ZN(n3609)
         );
  INV_X1 U3916 ( .A(n3609), .ZN(n3610) );
  OAI211_X1 U3917 ( .C1(n3612), .C2(n3011), .A(n3611), .B(n3610), .ZN(n3613)
         );
  INV_X1 U3918 ( .A(n3613), .ZN(n3619) );
  AOI22_X1 U3919 ( .A1(n3617), .A2(n3616), .B1(n3615), .B2(n3614), .ZN(n3618)
         );
  NAND4_X1 U3920 ( .A1(n3621), .A2(n3620), .A3(n3619), .A4(n3618), .ZN(n3622)
         );
  AOI211_X1 U3921 ( .C1(result_div[11]), .C2(n3988), .A(n3623), .B(n3622), 
        .ZN(n3631) );
  INV_X1 U3922 ( .A(n3637), .ZN(n3624) );
  OAI22_X1 U3923 ( .A1(n3624), .A2(n3990), .B1(n2562), .B2(n4021), .ZN(n3625)
         );
  OAI21_X1 U3924 ( .B1(n3626), .B2(n3625), .A(operand_a_i[11]), .ZN(n3630) );
  NAND2_X1 U3925 ( .A1(n3628), .A2(n3627), .ZN(n3629) );
  NAND4_X1 U3926 ( .A1(n3632), .A2(n3631), .A3(n3630), .A4(n3629), .ZN(n3633)
         );
  AOI21_X1 U3927 ( .B1(n3889), .B2(n4014), .A(n3633), .ZN(n3634) );
  OAI211_X1 U3928 ( .C1(n3636), .C2(n4192), .A(n3635), .B(n3634), .ZN(n3640)
         );
  OAI21_X1 U3929 ( .B1(n3144), .B2(n4122), .A(n4151), .ZN(n3638) );
  AOI22_X1 U3930 ( .A1(n3944), .A2(n4015), .B1(n4013), .B2(n4014), .ZN(n3676)
         );
  MUX2_X1 U3931 ( .A(n4017), .B(n3718), .S(operand_b_i[6]), .Z(n3671) );
  NAND2_X1 U3932 ( .A1(n4177), .A2(n3643), .ZN(n3669) );
  AOI22_X1 U3933 ( .A1(n4133), .A2(n3645), .B1(n4139), .B2(n3644), .ZN(n3661)
         );
  AOI22_X1 U3934 ( .A1(n4142), .A2(n3647), .B1(n4138), .B2(n3646), .ZN(n3660)
         );
  INV_X1 U3935 ( .A(n3648), .ZN(n3649) );
  OAI22_X1 U3936 ( .A1(n3650), .A2(n3722), .B1(n3721), .B2(n3649), .ZN(n3651)
         );
  INV_X1 U3937 ( .A(n3651), .ZN(n3659) );
  NOR2_X1 U3938 ( .A1(n3653), .A2(n3652), .ZN(n3654) );
  OAI22_X1 U3939 ( .A1(n3979), .A2(n3655), .B1(n4038), .B2(n3654), .ZN(n3656)
         );
  AOI21_X1 U3940 ( .B1(n4144), .B2(n3657), .A(n3656), .ZN(n3658) );
  NAND4_X1 U3941 ( .A1(n3661), .A2(n3660), .A3(n3659), .A4(n3658), .ZN(n3662)
         );
  AOI21_X1 U3942 ( .B1(n3988), .B2(result_div[6]), .A(n3662), .ZN(n3668) );
  INV_X1 U3943 ( .A(n3986), .ZN(n3667) );
  OAI22_X1 U3944 ( .A1(n3664), .A2(n3990), .B1(n3663), .B2(n4021), .ZN(n3665)
         );
  OAI21_X1 U3945 ( .B1(n4124), .B2(n3665), .A(operand_a_i[6]), .ZN(n3666) );
  NAND4_X1 U3946 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3670)
         );
  NOR2_X1 U3947 ( .A1(n3671), .A2(n3670), .ZN(n3675) );
  NAND2_X1 U3948 ( .A1(n3999), .A2(n4059), .ZN(n3674) );
  NAND2_X1 U3949 ( .A1(n4365), .A2(n3750), .ZN(n3673) );
  NAND4_X1 U3950 ( .A1(n3676), .A2(n3675), .A3(n3674), .A4(n3673), .ZN(n3680)
         );
  NAND2_X1 U3951 ( .A1(n4013), .A2(n4007), .ZN(n3678) );
  AOI21_X1 U3952 ( .B1(n3678), .B2(n4151), .A(n3677), .ZN(n3679) );
  OAI21_X1 U3953 ( .B1(n3965), .B2(n4122), .A(n4151), .ZN(n3714) );
  INV_X1 U3954 ( .A(n4012), .ZN(n3786) );
  AND2_X1 U3955 ( .A1(n4123), .A2(n4059), .ZN(n3710) );
  MUX2_X1 U3956 ( .A(n3683), .B(n4226), .S(ff1_result[1]), .Z(n3684) );
  OAI21_X1 U3957 ( .B1(n3686), .B2(n3685), .A(n3684), .ZN(n3701) );
  AOI22_X1 U3958 ( .A1(n4136), .A2(n4030), .B1(n4139), .B2(n3687), .ZN(n3696)
         );
  INV_X1 U3959 ( .A(n3688), .ZN(n4026) );
  AOI22_X1 U3960 ( .A1(n4026), .A2(n4133), .B1(n4138), .B2(n4028), .ZN(n3695)
         );
  AOI22_X1 U3961 ( .A1(n4154), .A2(n4042), .B1(n4142), .B2(n4024), .ZN(n3694)
         );
  NAND2_X1 U3962 ( .A1(result_div[1]), .A2(n3988), .ZN(n3691) );
  AOI22_X1 U3963 ( .A1(n4147), .A2(operand_c_i[1]), .B1(n4146), .B2(n3689), 
        .ZN(n3690) );
  NAND2_X1 U3964 ( .A1(n3691), .A2(n3690), .ZN(n3692) );
  AOI21_X1 U3965 ( .B1(n4144), .B2(n4044), .A(n3692), .ZN(n3693) );
  NAND4_X1 U3966 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3693), .ZN(n3697)
         );
  AOI21_X1 U3967 ( .B1(cnt_result[1]), .B2(n4169), .A(n3697), .ZN(n3698) );
  NAND2_X1 U3968 ( .A1(n4171), .A2(n3698), .ZN(n3699) );
  AOI21_X1 U3969 ( .B1(n3701), .B2(n3700), .A(n3699), .ZN(n3708) );
  INV_X1 U3970 ( .A(n3718), .ZN(n4178) );
  MUX2_X1 U3971 ( .A(n4179), .B(n4178), .S(operand_b_i[1]), .Z(n3707) );
  OAI22_X1 U3972 ( .A1(n3715), .A2(n3990), .B1(n2464), .B2(n3989), .ZN(n3703)
         );
  OAI21_X1 U3973 ( .B1(n4124), .B2(n3703), .A(n4225), .ZN(n3706) );
  NAND2_X1 U3974 ( .A1(n4177), .A2(n3704), .ZN(n3705) );
  NAND4_X1 U3975 ( .A1(n3708), .A2(n3707), .A3(n3706), .A4(n3705), .ZN(n3709)
         );
  AOI211_X1 U3976 ( .C1(n3711), .C2(n4014), .A(n3710), .B(n3709), .ZN(n3712)
         );
  OAI21_X1 U3977 ( .B1(n4193), .B2(n3786), .A(n3712), .ZN(n3713) );
  NAND2_X1 U3978 ( .A1(n3821), .A2(n4059), .ZN(n3748) );
  NOR2_X1 U3979 ( .A1(n3717), .A2(ff_no_one), .ZN(n4092) );
  MUX2_X1 U3980 ( .A(n4017), .B(n3718), .S(operand_b_i[5]), .Z(n3746) );
  NAND2_X1 U3981 ( .A1(n4177), .A2(n3719), .ZN(n3744) );
  OAI22_X1 U3982 ( .A1(n3723), .A2(n3722), .B1(n3721), .B2(n3720), .ZN(n3724)
         );
  AOI21_X1 U3983 ( .B1(n3988), .B2(result_div[5]), .A(n3724), .ZN(n3736) );
  AOI22_X1 U3984 ( .A1(n4142), .A2(n3726), .B1(n4138), .B2(n3725), .ZN(n3735)
         );
  OAI22_X1 U3985 ( .A1(n3979), .A2(n3728), .B1(n4038), .B2(n3727), .ZN(n3729)
         );
  AOI21_X1 U3986 ( .B1(n4139), .B2(n3730), .A(n3729), .ZN(n3734) );
  AOI22_X1 U3987 ( .A1(n4133), .A2(n3732), .B1(n4144), .B2(n3731), .ZN(n3733)
         );
  NAND4_X1 U3988 ( .A1(n3736), .A2(n3735), .A3(n3734), .A4(n3733), .ZN(n3737)
         );
  AOI211_X1 U3989 ( .C1(cnt_result[5]), .C2(n4169), .A(n3986), .B(n3737), .ZN(
        n3743) );
  OAI22_X1 U3990 ( .A1(n3755), .A2(n3990), .B1(n3738), .B2(n3989), .ZN(n3739)
         );
  OAI21_X1 U3991 ( .B1(n4124), .B2(n3739), .A(operand_a_i[5]), .ZN(n3742) );
  NAND3_X1 U3992 ( .A1(ff_no_one), .A2(n4337), .A3(n3740), .ZN(n3741) );
  NAND4_X1 U3993 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3745)
         );
  AOI211_X1 U3994 ( .C1(n4092), .C2(n3796), .A(n3746), .B(n3745), .ZN(n3747)
         );
  NAND2_X1 U3995 ( .A1(n3748), .A2(n3747), .ZN(n3749) );
  AOI21_X1 U3996 ( .B1(n3750), .B2(n3852), .A(n3749), .ZN(n3752) );
  NAND2_X1 U3997 ( .A1(n3794), .A2(n3944), .ZN(n3751) );
  OAI211_X1 U3998 ( .C1(n4121), .C2(n3753), .A(n3752), .B(n3751), .ZN(n3757)
         );
  OAI21_X1 U3999 ( .B1(n3753), .B2(n4122), .A(n4151), .ZN(n3756) );
  INV_X1 U4000 ( .A(n3767), .ZN(n3762) );
  OAI21_X1 U4001 ( .B1(n3759), .B2(n4122), .A(n4151), .ZN(n3760) );
  INV_X1 U4002 ( .A(n3763), .ZN(n3787) );
  OAI21_X1 U4003 ( .B1(operand_a_i[16]), .B2(n4038), .A(n3890), .ZN(n3764) );
  MUX2_X1 U4004 ( .A(n4017), .B(n3764), .S(operand_b_i[16]), .Z(n3784) );
  MUX2_X1 U4005 ( .A(n4125), .B(n4146), .S(n3765), .Z(n3766) );
  AOI211_X1 U4006 ( .C1(n4126), .C2(n3767), .A(n3766), .B(n3921), .ZN(n3782)
         );
  INV_X1 U4007 ( .A(n4135), .ZN(n3769) );
  OAI22_X1 U4008 ( .A1(n3770), .A2(n3769), .B1(n4040), .B2(n3768), .ZN(n3773)
         );
  NOR2_X1 U4009 ( .A1(n3911), .A2(n3771), .ZN(n3772) );
  AOI211_X1 U4010 ( .C1(n3908), .C2(n4153), .A(n3773), .B(n3772), .ZN(n3777)
         );
  AOI22_X1 U4011 ( .A1(n3906), .A2(n4137), .B1(n3894), .B2(n4141), .ZN(n3774)
         );
  OAI21_X1 U4012 ( .B1(n3899), .B2(n4132), .A(n3774), .ZN(n3775) );
  AOI21_X1 U4013 ( .B1(n3892), .B2(n4143), .A(n3775), .ZN(n3776) );
  OAI211_X1 U4014 ( .C1(n4127), .C2(n3901), .A(n3777), .B(n3776), .ZN(n3778)
         );
  AOI211_X1 U4015 ( .C1(result_div[16]), .C2(n3988), .A(n3917), .B(n3778), 
        .ZN(n3781) );
  NAND2_X1 U4016 ( .A1(n3923), .A2(n3779), .ZN(n3780) );
  OAI211_X1 U4017 ( .C1(n3782), .C2(n4097), .A(n3781), .B(n3780), .ZN(n3783)
         );
  AOI211_X1 U4018 ( .C1(n2968), .C2(n4014), .A(n3784), .B(n3783), .ZN(n3785)
         );
  OAI21_X1 U4019 ( .B1(n3787), .B2(n3786), .A(n3785), .ZN(n3790) );
  NAND2_X1 U4020 ( .A1(n3792), .A2(n941), .ZN(n3829) );
  OAI21_X1 U4021 ( .B1(n3793), .B2(n4122), .A(n4151), .ZN(n3826) );
  INV_X1 U4022 ( .A(n3794), .ZN(n3824) );
  MUX2_X1 U4023 ( .A(n4161), .B(n3882), .S(ff1_result[4]), .Z(n3795) );
  AOI21_X1 U4024 ( .B1(n3797), .B2(n3796), .A(n3795), .ZN(n3818) );
  NAND2_X1 U4025 ( .A1(cnt_result[4]), .A2(n4169), .ZN(n3809) );
  OAI22_X1 U4026 ( .A1(n3979), .A2(n3799), .B1(n4038), .B2(n3798), .ZN(n3800)
         );
  AOI21_X1 U4027 ( .B1(result_div[4]), .B2(n3988), .A(n3800), .ZN(n3802) );
  NAND2_X1 U4028 ( .A1(n4142), .A2(n3893), .ZN(n3801) );
  AND2_X1 U4029 ( .A1(n3802), .A2(n3801), .ZN(n3807) );
  INV_X1 U4030 ( .A(n3865), .ZN(n3891) );
  AOI22_X1 U4031 ( .A1(n3891), .A2(n4144), .B1(n4139), .B2(n3803), .ZN(n3806)
         );
  AOI22_X1 U4032 ( .A1(n4136), .A2(n3895), .B1(n4138), .B2(n3905), .ZN(n3805)
         );
  AOI22_X1 U4033 ( .A1(n4154), .A2(n3907), .B1(n4133), .B2(n3857), .ZN(n3804)
         );
  AND4_X1 U4034 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3808)
         );
  NAND3_X1 U4035 ( .A1(n3809), .A2(n4171), .A3(n3808), .ZN(n3810) );
  AOI21_X1 U4036 ( .B1(n4177), .B2(n3811), .A(n3810), .ZN(n3815) );
  OAI22_X1 U4037 ( .A1(n3827), .A2(n3990), .B1(n3812), .B2(n4021), .ZN(n3813)
         );
  OAI21_X1 U4038 ( .B1(n4124), .B2(n3813), .A(operand_a_i[4]), .ZN(n3814) );
  AND2_X1 U4039 ( .A1(n3815), .A2(n3814), .ZN(n3817) );
  MUX2_X1 U4040 ( .A(n4179), .B(n4178), .S(operand_b_i[4]), .Z(n3816) );
  OAI211_X1 U4041 ( .C1(n3818), .C2(n4172), .A(n3817), .B(n3816), .ZN(n3819)
         );
  AOI21_X1 U4042 ( .B1(n3820), .B2(n4014), .A(n3819), .ZN(n3823) );
  NAND2_X1 U4043 ( .A1(n3821), .A2(n4012), .ZN(n3822) );
  OAI211_X1 U4044 ( .C1(n3824), .C2(n4192), .A(n3823), .B(n3822), .ZN(n3825)
         );
  NAND2_X1 U4045 ( .A1(n3829), .A2(n3828), .ZN(result_o[4]) );
  OR4_X1 U4046 ( .A1(cnt_result[0]), .A2(cnt_result[3]), .A3(cnt_result[4]), 
        .A4(cnt_result[5]), .ZN(n3830) );
  NOR3_X1 U4047 ( .A1(cnt_result[1]), .A2(cnt_result[2]), .A3(n3830), .ZN(
        n2389) );
  AND2_X1 U4048 ( .A1(n4289), .A2(n3834), .ZN(n3836) );
  OAI21_X1 U4049 ( .B1(n3837), .B2(n3836), .A(int_div_div_op_a_signed), .ZN(
        n3840) );
  MUX2_X1 U4050 ( .A(n4228), .B(n4113), .S(n4087), .Z(n3838) );
  OAI21_X1 U4051 ( .B1(n4088), .B2(n53), .A(n3838), .ZN(ff_input[29]) );
  MUX2_X1 U4052 ( .A(n4085), .B(n4099), .S(operand_a_i[17]), .Z(n3839) );
  OAI21_X1 U4053 ( .B1(n4227), .B2(n4098), .A(n3839), .ZN(ff_input[14]) );
  MUX2_X1 U4054 ( .A(n4099), .B(n4085), .S(n71), .Z(n3841) );
  OAI21_X1 U4055 ( .B1(n4116), .B2(n4101), .A(n3841), .ZN(ff_input[13]) );
  MUX2_X1 U4056 ( .A(n4099), .B(n4085), .S(n4105), .Z(n3842) );
  OAI21_X1 U4057 ( .B1(n4227), .B2(n2561), .A(n3842), .ZN(ff_input[12]) );
  MUX2_X1 U4058 ( .A(n4229), .B(n4113), .S(n2543), .Z(n3843) );
  OAI21_X1 U4059 ( .B1(n4088), .B2(n3844), .A(n3843), .ZN(ff_input[24]) );
  OAI21_X1 U4060 ( .B1(n4226), .B2(n3846), .A(n3845), .ZN(ff_input[25]) );
  MUX2_X1 U4061 ( .A(n4228), .B(n4085), .S(n4079), .Z(n3847) );
  OAI21_X1 U4062 ( .B1(n4226), .B2(n3848), .A(n3847), .ZN(ff_input[26]) );
  OAI21_X1 U4064 ( .B1(n3849), .B2(n4122), .A(n4151), .ZN(n3850) );
  NAND2_X1 U4065 ( .A1(n3852), .A2(n4014), .ZN(n3879) );
  NAND2_X1 U4066 ( .A1(n3853), .A2(n4012), .ZN(n3878) );
  MUX2_X1 U4067 ( .A(n4017), .B(n4016), .S(operand_b_i[28]), .Z(n3874) );
  OAI22_X1 U4068 ( .A1(n3855), .A2(n3990), .B1(n3854), .B2(n4021), .ZN(n3856)
         );
  OAI21_X1 U4069 ( .B1(n4023), .B2(n3856), .A(operand_a_i[28]), .ZN(n3872) );
  AOI22_X1 U4070 ( .A1(n4027), .A2(n3857), .B1(n4025), .B2(n3893), .ZN(n3859)
         );
  AOI22_X1 U4071 ( .A1(n4031), .A2(n3895), .B1(n4029), .B2(n3905), .ZN(n3858)
         );
  OAI211_X1 U4072 ( .C1(n4034), .C2(n3912), .A(n3859), .B(n3858), .ZN(n3868)
         );
  NAND2_X1 U4073 ( .A1(n4036), .A2(operand_a_i[4]), .ZN(n3864) );
  OAI22_X1 U4074 ( .A1(n4040), .A2(n3861), .B1(n4038), .B2(n3860), .ZN(n3862)
         );
  AOI21_X1 U4075 ( .B1(n4043), .B2(n3907), .A(n3862), .ZN(n3863) );
  OAI211_X1 U4076 ( .C1(n3866), .C2(n3865), .A(n3864), .B(n3863), .ZN(n3867)
         );
  NOR2_X1 U4077 ( .A1(n3868), .A2(n3867), .ZN(n3871) );
  NAND2_X1 U4078 ( .A1(n4052), .A2(n3869), .ZN(n3870) );
  NAND4_X1 U4079 ( .A1(n3872), .A2(n3871), .A3(n4054), .A4(n3870), .ZN(n3873)
         );
  AOI211_X1 U4080 ( .C1(result_div[28]), .C2(n3988), .A(n3874), .B(n3873), 
        .ZN(n3877) );
  NAND2_X1 U4081 ( .A1(n3875), .A2(n4059), .ZN(n3876) );
  NAND4_X1 U4082 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3880)
         );
  OAI21_X1 U4083 ( .B1(n4116), .B2(n4075), .A(n3881), .ZN(ff_input[21]) );
  MUX2_X1 U4084 ( .A(n4085), .B(n4229), .S(operand_a_i[9]), .Z(n3883) );
  OAI21_X1 U4085 ( .B1(n4226), .B2(n4072), .A(n3883), .ZN(ff_input[22]) );
  OAI21_X1 U4086 ( .B1(n4088), .B2(n4067), .A(n3884), .ZN(ff_input[20]) );
  AOI21_X1 U4088 ( .B1(n3321), .B2(n4007), .A(n4006), .ZN(n3886) );
  INV_X1 U4089 ( .A(n3886), .ZN(n3887) );
  AOI22_X1 U4090 ( .A1(n125), .A2(n4059), .B1(n3889), .B2(n3944), .ZN(n3933)
         );
  MUX2_X1 U4091 ( .A(n4179), .B(n3890), .S(operand_b_i[20]), .Z(n3927) );
  NAND2_X1 U4092 ( .A1(n3892), .A2(n3891), .ZN(n3898) );
  AOI22_X1 U4093 ( .A1(n3896), .A2(n3895), .B1(n3894), .B2(n3893), .ZN(n3897)
         );
  OAI211_X1 U4094 ( .C1(n3900), .C2(n3899), .A(n3898), .B(n3897), .ZN(n3916)
         );
  NOR2_X1 U4095 ( .A1(n3901), .A2(n4108), .ZN(n3914) );
  OAI22_X1 U4096 ( .A1(n4040), .A2(n3903), .B1(n4038), .B2(n3902), .ZN(n3904)
         );
  AOI21_X1 U4097 ( .B1(n3906), .B2(n3905), .A(n3904), .ZN(n3910) );
  NAND2_X1 U4098 ( .A1(n3908), .A2(n3907), .ZN(n3909) );
  OAI211_X1 U4099 ( .C1(n3912), .C2(n3911), .A(n3910), .B(n3909), .ZN(n3913)
         );
  OR2_X1 U4100 ( .A1(n3914), .A2(n3913), .ZN(n3915) );
  NOR3_X1 U4101 ( .A1(n3917), .A2(n3916), .A3(n3915), .ZN(n3926) );
  OAI22_X1 U4102 ( .A1(n3919), .A2(n3990), .B1(n3918), .B2(n4021), .ZN(n3920)
         );
  OAI21_X1 U4103 ( .B1(n3921), .B2(n3920), .A(operand_a_i[20]), .ZN(n3925) );
  NAND2_X1 U4104 ( .A1(n3923), .A2(n3922), .ZN(n3924) );
  NAND4_X1 U4105 ( .A1(n3927), .A2(n3926), .A3(n3925), .A4(n3924), .ZN(n3928)
         );
  AOI21_X1 U4106 ( .B1(result_div[20]), .B2(n3988), .A(n3928), .ZN(n3929) );
  INV_X1 U4107 ( .A(n3929), .ZN(n3930) );
  AOI21_X1 U4108 ( .B1(n3321), .B2(n4014), .A(n3930), .ZN(n3932) );
  OAI211_X1 U4109 ( .C1(n3934), .C2(n4184), .A(n3933), .B(n3932), .ZN(n3935)
         );
  NAND2_X1 U4110 ( .A1(n4123), .A2(n4007), .ZN(n3936) );
  NAND2_X1 U4111 ( .A1(n3936), .A2(n4151), .ZN(n3943) );
  OAI22_X1 U4112 ( .A1(n4310), .A2(n3937), .B1(n3990), .B2(n4115), .ZN(n3938)
         );
  NAND2_X1 U4115 ( .A1(result_div[31]), .A2(n3988), .ZN(n3968) );
  AOI22_X1 U4116 ( .A1(n3944), .A2(n4316), .B1(n4123), .B2(n4014), .ZN(n3967)
         );
  MUX2_X1 U4117 ( .A(n4017), .B(n4016), .S(operand_b_i[31]), .Z(n3964) );
  NAND2_X1 U4118 ( .A1(n4023), .A2(n4304), .ZN(n3962) );
  INV_X1 U4119 ( .A(n3945), .ZN(n3973) );
  AOI22_X1 U4120 ( .A1(n4027), .A2(n3973), .B1(n4029), .B2(n3981), .ZN(n3947)
         );
  AOI22_X1 U4121 ( .A1(n4031), .A2(n3975), .B1(n4025), .B2(n3974), .ZN(n3946)
         );
  OAI211_X1 U4122 ( .C1(n4034), .C2(n3948), .A(n3947), .B(n3946), .ZN(n3958)
         );
  NAND2_X1 U4123 ( .A1(n4036), .A2(operand_a_i[7]), .ZN(n3956) );
  OAI22_X1 U4124 ( .A1(n4038), .A2(n3950), .B1(n148), .B2(n4021), .ZN(n3951)
         );
  AOI21_X1 U4125 ( .B1(n3952), .B2(operand_c_i[31]), .A(n3951), .ZN(n3955) );
  NAND2_X1 U4126 ( .A1(n4045), .A2(n3972), .ZN(n3954) );
  NAND2_X1 U4127 ( .A1(n4043), .A2(n3971), .ZN(n3953) );
  NAND4_X1 U4128 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(n3957)
         );
  NOR2_X1 U4129 ( .A1(n3958), .A2(n3957), .ZN(n3961) );
  NAND2_X1 U4130 ( .A1(n4052), .A2(n3959), .ZN(n3960) );
  NAND4_X1 U4131 ( .A1(n3962), .A2(n3961), .A3(n4054), .A4(n3960), .ZN(n3963)
         );
  NOR2_X1 U4132 ( .A1(n3964), .A2(n3963), .ZN(n3966) );
  MUX2_X1 U4133 ( .A(n4179), .B(n4178), .S(operand_b_i[7]), .Z(n3996) );
  AOI22_X1 U4134 ( .A1(n4154), .A2(n3971), .B1(n4139), .B2(n3970), .ZN(n3985)
         );
  AOI22_X1 U4135 ( .A1(n4133), .A2(n3973), .B1(n4144), .B2(n3972), .ZN(n3984)
         );
  AOI22_X1 U4136 ( .A1(n4136), .A2(n3975), .B1(n4142), .B2(n3974), .ZN(n3983)
         );
  INV_X1 U4137 ( .A(n3976), .ZN(n3977) );
  OAI22_X1 U4138 ( .A1(n3979), .A2(n3978), .B1(n4038), .B2(n3977), .ZN(n3980)
         );
  AOI21_X1 U4139 ( .B1(n4138), .B2(n3981), .A(n3980), .ZN(n3982) );
  NAND4_X1 U4140 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3987)
         );
  AOI211_X1 U4141 ( .C1(n3988), .C2(result_div[7]), .A(n3987), .B(n3986), .ZN(
        n3995) );
  OAI22_X1 U4142 ( .A1(n4004), .A2(n3990), .B1(n588), .B2(n3989), .ZN(n3991)
         );
  OAI21_X1 U4143 ( .B1(n4124), .B2(n3991), .A(operand_a_i[7]), .ZN(n3994) );
  NAND2_X1 U4144 ( .A1(n4177), .A2(n3992), .ZN(n3993) );
  NAND4_X1 U4145 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n3998)
         );
  NOR2_X1 U4146 ( .A1(n4000), .A2(n4121), .ZN(n3997) );
  AOI211_X1 U4147 ( .C1(n4012), .C2(n3999), .A(n3998), .B(n3997), .ZN(n4003)
         );
  OAI21_X1 U4148 ( .B1(n4000), .B2(n4122), .A(n4151), .ZN(n4001) );
  AOI22_X1 U4149 ( .A1(n4001), .A2(n4004), .B1(n4059), .B2(n4015), .ZN(n4002)
         );
  OAI211_X1 U4150 ( .C1(n4005), .C2(n4004), .A(n4003), .B(n4002), .ZN(
        result_o[7]) );
  AOI21_X1 U4151 ( .B1(n4015), .B2(n4007), .A(n4006), .ZN(n4008) );
  INV_X1 U4152 ( .A(n4008), .ZN(n4011) );
  NAND2_X1 U4154 ( .A1(n4013), .A2(n4012), .ZN(n4064) );
  NAND2_X1 U4155 ( .A1(n4015), .A2(n4014), .ZN(n4063) );
  MUX2_X1 U4156 ( .A(n4017), .B(n4016), .S(n110), .Z(n4058) );
  NAND2_X1 U4157 ( .A1(n4018), .A2(n4126), .ZN(n4019) );
  OAI21_X1 U4158 ( .B1(n4021), .B2(n4020), .A(n4019), .ZN(n4022) );
  OAI21_X1 U4159 ( .B1(n4023), .B2(n4022), .A(operand_a_i[25]), .ZN(n4056) );
  AOI22_X1 U4160 ( .A1(n4027), .A2(n4026), .B1(n4025), .B2(n4024), .ZN(n4033)
         );
  AOI22_X1 U4161 ( .A1(n4031), .A2(n4030), .B1(n4029), .B2(n4028), .ZN(n4032)
         );
  OAI211_X1 U4162 ( .C1(n4035), .C2(n4034), .A(n4033), .B(n4032), .ZN(n4050)
         );
  NAND2_X1 U4163 ( .A1(n4036), .A2(n4225), .ZN(n4048) );
  OAI22_X1 U4164 ( .A1(n4040), .A2(n4039), .B1(n4038), .B2(n4037), .ZN(n4041)
         );
  AOI21_X1 U4165 ( .B1(n4043), .B2(n4042), .A(n4041), .ZN(n4047) );
  NAND2_X1 U4166 ( .A1(n4045), .A2(n4044), .ZN(n4046) );
  NAND3_X1 U4167 ( .A1(n4048), .A2(n4047), .A3(n4046), .ZN(n4049) );
  NOR2_X1 U4168 ( .A1(n4050), .A2(n4049), .ZN(n4055) );
  NAND2_X1 U4169 ( .A1(n4052), .A2(n4051), .ZN(n4053) );
  NAND4_X1 U4170 ( .A1(n4056), .A2(n4055), .A3(n4054), .A4(n4053), .ZN(n4057)
         );
  AOI211_X1 U4171 ( .C1(result_div[25]), .C2(n3988), .A(n4058), .B(n4057), 
        .ZN(n4062) );
  NAND2_X1 U4172 ( .A1(n4305), .A2(n4059), .ZN(n4061) );
  NAND4_X1 U4173 ( .A1(n4064), .A2(n4063), .A3(n4062), .A4(n4061), .ZN(n4065)
         );
  MUX2_X1 U4174 ( .A(n4085), .B(n4099), .S(operand_a_i[24]), .Z(n4066) );
  OAI21_X1 U4175 ( .B1(n4226), .B2(n2543), .A(n4066), .ZN(ff_input[7]) );
  OAI21_X1 U4176 ( .B1(n4088), .B2(n4069), .A(n4068), .ZN(ff_input[11]) );
  MUX2_X1 U4177 ( .A(n4085), .B(n4228), .S(operand_a_i[25]), .Z(n4070) );
  OAI21_X1 U4178 ( .B1(n4088), .B2(n4071), .A(n4070), .ZN(ff_input[6]) );
  INV_X1 U4179 ( .A(operand_a_i[9]), .ZN(n4074) );
  OAI21_X1 U4180 ( .B1(n4227), .B2(n4074), .A(n4073), .ZN(ff_input[9]) );
  OAI21_X1 U4181 ( .B1(n4227), .B2(n2570), .A(n4076), .ZN(ff_input[10]) );
  OAI21_X1 U4182 ( .B1(n4088), .B2(n4106), .A(n4077), .ZN(ff_input[8]) );
  OAI21_X1 U4183 ( .B1(n4116), .B2(n4079), .A(n4078), .ZN(ff_input[5]) );
  OAI21_X1 U4184 ( .B1(n4116), .B2(n4108), .A(n4080), .ZN(ff_input[4]) );
  OAI21_X1 U4185 ( .B1(n4227), .B2(n3011), .A(n4081), .ZN(ff_input[3]) );
  MUX2_X1 U4186 ( .A(n4099), .B(n4113), .S(n4112), .Z(n4083) );
  OAI21_X1 U4187 ( .B1(n4116), .B2(n2546), .A(n4083), .ZN(ff_input[1]) );
  OAI21_X1 U4188 ( .B1(n4088), .B2(n4087), .A(n4086), .ZN(ff_input[2]) );
  INV_X1 U4189 ( .A(n4089), .ZN(n4090) );
  NOR2_X1 U4190 ( .A1(n4090), .A2(n4092), .ZN(n4093) );
  MUX2_X1 U4191 ( .A(n4093), .B(n4092), .S(n4091), .Z(div_shift[5]) );
  MUX2_X1 U4192 ( .A(n4085), .B(n4228), .S(operand_a_i[16]), .Z(n4094) );
  OAI21_X1 U4193 ( .B1(n4226), .B2(n4095), .A(n4094), .ZN(ff_input[15]) );
  OAI21_X1 U4194 ( .B1(n4227), .B2(n4097), .A(n4096), .ZN(ff_input[16]) );
  MUX2_X1 U4195 ( .A(n4229), .B(n4113), .S(n4098), .Z(n4100) );
  OAI21_X1 U4196 ( .B1(n4088), .B2(n71), .A(n4102), .ZN(ff_input[18]) );
  OAI21_X1 U4197 ( .B1(n4116), .B2(n4105), .A(n4104), .ZN(ff_input[19]) );
  MUX2_X1 U4198 ( .A(n4228), .B(n4113), .S(n4106), .Z(n4107) );
  OAI21_X1 U4199 ( .B1(n4116), .B2(n585), .A(n4107), .ZN(ff_input[23]) );
  MUX2_X1 U4200 ( .A(n4228), .B(n4085), .S(n4108), .Z(n4109) );
  OAI21_X1 U4201 ( .B1(n4227), .B2(n2521), .A(n4109), .ZN(ff_input[27]) );
  MUX2_X1 U4202 ( .A(n4085), .B(n4228), .S(n48), .Z(n4110) );
  OAI21_X1 U4203 ( .B1(n4116), .B2(n2522), .A(n4110), .ZN(ff_input[28]) );
  MUX2_X1 U4204 ( .A(n4229), .B(n4085), .S(n2546), .Z(n4111) );
  OAI21_X1 U4205 ( .B1(n4227), .B2(n4112), .A(n4111), .ZN(ff_input[30]) );
  MUX2_X1 U4206 ( .A(n4229), .B(n4113), .S(n4127), .Z(n4114) );
  OAI21_X1 U4207 ( .B1(n4116), .B2(n4115), .A(n4114), .ZN(ff_input[31]) );
  NAND2_X1 U4208 ( .A1(n4120), .A2(n4119), .ZN(n4150) );
  OAI21_X1 U4209 ( .B1(n4122), .B2(n4150), .A(n4121), .ZN(n4188) );
  INV_X1 U4210 ( .A(n4123), .ZN(n4183) );
  INV_X1 U4211 ( .A(n4124), .ZN(n4129) );
  AOI22_X1 U4212 ( .A1(n4126), .A2(n4150), .B1(n4125), .B2(operand_b_i[0]), 
        .ZN(n4128) );
  AOI21_X1 U4213 ( .B1(n4129), .B2(n4128), .A(n4127), .ZN(n4175) );
  MUX2_X1 U4214 ( .A(n4131), .B(n4130), .S(n4283), .Z(n4173) );
  INV_X1 U4215 ( .A(n4132), .ZN(n4134) );
  AOI22_X1 U4216 ( .A1(n4136), .A2(n4135), .B1(n4134), .B2(n4133), .ZN(n4158)
         );
  AOI22_X1 U4217 ( .A1(n4140), .A2(n4139), .B1(n4138), .B2(n4137), .ZN(n4157)
         );
  AOI22_X1 U4218 ( .A1(n4144), .A2(n4143), .B1(n4142), .B2(n4141), .ZN(n4156)
         );
  AOI22_X1 U4219 ( .A1(n4146), .A2(n4145), .B1(n3988), .B2(result_div[0]), 
        .ZN(n4149) );
  NAND2_X1 U4220 ( .A1(n4147), .A2(operand_c_i[0]), .ZN(n4148) );
  OAI211_X1 U4221 ( .C1(n4151), .C2(n4150), .A(n4149), .B(n4148), .ZN(n4152)
         );
  AOI21_X1 U4222 ( .B1(n4154), .B2(n4153), .A(n4152), .ZN(n4155) );
  NAND4_X1 U4223 ( .A1(n4158), .A2(n4157), .A3(n4156), .A4(n4155), .ZN(n4168)
         );
  NAND3_X1 U4224 ( .A1(n4161), .A2(n4160), .A3(n4159), .ZN(n4166) );
  MUX2_X1 U4225 ( .A(n4163), .B(n4162), .S(n4337), .Z(n4165) );
  INV_X1 U4226 ( .A(n2832), .ZN(n4164) );
  AOI21_X1 U4227 ( .B1(n4166), .B2(n4165), .A(n4164), .ZN(n4167) );
  AOI211_X1 U4228 ( .C1(n4169), .C2(cnt_result[0]), .A(n4168), .B(n4167), .ZN(
        n4170) );
  OAI211_X1 U4229 ( .C1(n4173), .C2(n4172), .A(n4171), .B(n4170), .ZN(n4174)
         );
  AOI211_X1 U4230 ( .C1(n4177), .C2(n4176), .A(n4175), .B(n4174), .ZN(n4181)
         );
  MUX2_X1 U4231 ( .A(n4179), .B(n4178), .S(operand_b_i[0]), .Z(n4180) );
  OAI211_X1 U4232 ( .C1(n4183), .C2(n4182), .A(n4181), .B(n4180), .ZN(n4187)
         );
  NOR2_X1 U4233 ( .A1(n4185), .A2(n4184), .ZN(n4186) );
  OR2_X2 U170 ( .A1(n2329), .A2(n2130), .ZN(n2170) );
  OR2_X2 U942 ( .A1(n2120), .A2(n1794), .ZN(n2155) );
  NOR2_X2 U2580 ( .A1(n2333), .A2(n2290), .ZN(n2296) );
  AOI21_X2 U183 ( .B1(n478), .B2(n82), .A(n1287), .ZN(n1944) );
  NOR2_X2 U122 ( .A1(n638), .A2(n637), .ZN(n979) );
  alu_popcnt alu_popcnt_i ( .in_i({n4304, operand_a_i[30], n54, 
        operand_a_i[28:19], n72, operand_a_i[17:15], n4300, operand_a_i[13], 
        n163, operand_a_i[11], n167, operand_a_i[9], n149, operand_a_i[7:4], 
        n48, operand_a_i[2], n4225, n4198}), .result_o(cnt_result) );
  alu_ff alu_ff_i ( .in_i(ff_input), .first_one_o(ff1_result), .no_ones_o(
        ff_no_one) );
  riscv_alu_div int_div_div_i ( .Clk_CI(clk), .Rst_RBI(rst_n), .OpA_DI({
        operand_b_i[31:28], n64, n170, n110, n4340, operand_b_i[23:19], n4194, 
        n4328, operand_b_i[16:12], n150, operand_b_i[10], n4195, n4196, 
        operand_b_i[7:0]}), .OpB_DI({n2421, n2420, n2419, n2418, n2417, n2416, 
        n2415, n2414, n2413, n2412, n2411, n2410, n2409, n4224, n2407, n2406, 
        n2405, n2404, n2403, n4275, n4284, n2400, n2399, n2398, n2397, n2396, 
        n2395, n2394, n2393, n2392, n2391, n2390}), .OpBShift_DI({
        div_shift[5:4], n2844, div_shift[2:0]}), .OpBIsZero_SI(n2389), 
        .OpBSign_SI(int_div_div_op_a_signed), .OpCode_SI({n4337, n52}), 
        .InVld_SI(div_valid), .OutRdy_SI(ex_ready_i), .OutVld_SO(ready_o), 
        .Res_DO(result_div) );
  BUF_X2 U1148 ( .A(n587), .Z(n775) );
  MUX2_X2 U476 ( .A(n2401), .B(n2410), .S(n91), .Z(n3321) );
  AOI21_X1 U212 ( .B1(n866), .B2(n672), .A(n136), .ZN(n783) );
  AND3_X2 U2348 ( .A1(n1760), .A2(n1759), .A3(n1758), .ZN(n2214) );
  INV_X2 U679 ( .A(n4118), .ZN(n3642) );
  BUF_X2 U176 ( .A(n1587), .Z(n1702) );
  OAI21_X1 U119 ( .B1(n1312), .B2(n1306), .A(n1307), .ZN(n1290) );
  AND2_X1 U40 ( .A1(n1684), .A2(n1678), .ZN(n42) );
  NOR2_X1 U32 ( .A1(n2495), .A2(n3380), .ZN(n397) );
  INV_X1 U1172 ( .A(operand_a_i[28]), .ZN(n2522) );
  BUF_X1 U52 ( .A(operand_a_i[3]), .Z(n48) );
  INV_X1 U15 ( .A(bmask_b_i[2]), .ZN(n1076) );
  OR2_X2 U247 ( .A1(operator_i[0]), .A2(operator_i[1]), .ZN(n3380) );
  INV_X2 U1197 ( .A(operand_a_i[21]), .ZN(n4075) );
  INV_X1 U1241 ( .A(operand_a_i[31]), .ZN(n4115) );
  INV_X1 U882 ( .A(operand_a_i[23]), .ZN(n585) );
  INV_X1 U557 ( .A(operand_a_i[27]), .ZN(n2521) );
  INV_X1 U16 ( .A(bmask_a_i[4]), .ZN(n2369) );
  CLKBUF_X1 U20 ( .A(operand_b_i[8]), .Z(n4196) );
  INV_X1 U240 ( .A(n1218), .ZN(n1171) );
  AND2_X1 U81 ( .A1(n497), .A2(operator_i[2]), .ZN(n2647) );
  NAND2_X1 U990 ( .A1(n4337), .A2(n52), .ZN(n3683) );
  OR2_X1 U572 ( .A1(n2495), .A2(n504), .ZN(n532) );
  AND4_X1 U53 ( .A1(n3533), .A2(n2821), .A3(n3950), .A4(n3295), .ZN(n283) );
  INV_X2 U126 ( .A(n532), .ZN(n82) );
  CLKBUF_X1 U128 ( .A(n218), .Z(n2660) );
  BUF_X2 U1038 ( .A(n558), .Z(n1205) );
  BUF_X2 U47 ( .A(n558), .Z(n704) );
  OR2_X1 U906 ( .A1(n2662), .A2(n2495), .ZN(n546) );
  CLKBUF_X2 U77 ( .A(n3840), .Z(n4113) );
  INV_X1 U340 ( .A(n3882), .ZN(n4088) );
  NOR2_X1 U101 ( .A1(n670), .A2(n671), .ZN(n872) );
  OR2_X1 U224 ( .A1(n575), .A2(n82), .ZN(n1545) );
  NOR2_X1 U221 ( .A1(n645), .A2(n644), .ZN(n923) );
  CLKBUF_X1 U343 ( .A(n2753), .Z(n154) );
  AND2_X1 U90 ( .A1(n91), .A2(n2784), .ZN(n1605) );
  NOR2_X1 U316 ( .A1(n745), .A2(n748), .ZN(n770) );
  OR2_X1 U64 ( .A1(n3242), .A2(n1030), .ZN(n1536) );
  NOR2_X1 U339 ( .A1(ff1_result[0]), .A2(ff1_result[1]), .ZN(n492) );
  INV_X1 U198 ( .A(n4017), .ZN(n4179) );
  INV_X1 U2036 ( .A(n1458), .ZN(n1543) );
  OAI21_X1 U116 ( .B1(n518), .B2(n90), .A(n432), .ZN(n2169) );
  INV_X1 U721 ( .A(n1788), .ZN(n1620) );
  AOI21_X1 U24 ( .B1(n1584), .B2(n1605), .A(n1583), .ZN(n2151) );
  NAND2_X1 U186 ( .A1(n392), .A2(n395), .ZN(n2000) );
  CLKBUF_X1 U171 ( .A(n1629), .Z(n1776) );
  AND4_X1 U165 ( .A1(n1799), .A2(n1798), .A3(n1800), .A4(n1797), .ZN(n2269) );
  MUX2_X1 U2751 ( .A(n2416), .B(n2395), .S(n2376), .Z(n3794) );
  AND2_X1 U140 ( .A1(bmask_a_i[0]), .A2(bmask_a_i[1]), .ZN(n2372) );
  INV_X2 U1036 ( .A(is_subrot_i), .ZN(n540) );
  NOR2_X1 U1067 ( .A1(bmask_a_i[0]), .A2(bmask_a_i[1]), .ZN(n2368) );
  CLKBUF_X1 U13 ( .A(operand_b_i[25]), .Z(n110) );
  BUF_X1 U56 ( .A(operator_i[0]), .Z(n52) );
  AND3_X1 U699 ( .A1(n283), .A2(n284), .A3(n3860), .ZN(n2604) );
  CLKBUF_X2 U231 ( .A(n3840), .Z(n4085) );
  CLKBUF_X2 U558 ( .A(n587), .Z(n1128) );
  INV_X2 U124 ( .A(n2106), .ZN(n92) );
  BUF_X2 U97 ( .A(n575), .Z(n91) );
  INV_X1 U12 ( .A(n91), .ZN(n1544) );
  OR2_X1 U121 ( .A1(n1532), .A2(n505), .ZN(n1871) );
  BUF_X2 U115 ( .A(n1270), .Z(n1315) );
  AOI21_X1 U181 ( .B1(n358), .B2(n82), .A(n1305), .ZN(n2194) );
  MUX2_X1 U2540 ( .A(n2001), .B(n2058), .S(n2000), .Z(n2289) );
  OR2_X1 U95 ( .A1(n3833), .A2(n3832), .ZN(n4099) );
  BUF_X1 U5 ( .A(n3145), .Z(n3558) );
  BUF_X1 U6 ( .A(n2310), .Z(n4233) );
  OR2_X1 U8 ( .A1(n2323), .A2(n1845), .ZN(n2162) );
  BUF_X1 U10 ( .A(n85), .Z(n4287) );
  OR2_X1 U17 ( .A1(n3833), .A2(n3832), .ZN(n4228) );
  OR2_X1 U18 ( .A1(n3833), .A2(n3832), .ZN(n4229) );
  BUF_X1 U21 ( .A(operator_i[2]), .Z(n2648) );
  NAND2_X1 U28 ( .A1(ff1_result[0]), .A2(n112), .ZN(n494) );
  AND2_X2 U35 ( .A1(n4356), .A2(n4355), .ZN(n1321) );
  BUF_X1 U37 ( .A(operator_i[5]), .Z(n4307) );
  INV_X2 U38 ( .A(n2178), .ZN(n2174) );
  INV_X2 U39 ( .A(n2105), .ZN(n2305) );
  INV_X1 U46 ( .A(n3882), .ZN(n4226) );
  INV_X1 U51 ( .A(n3882), .ZN(n4227) );
  INV_X2 U54 ( .A(n3882), .ZN(n4116) );
  AND2_X2 U55 ( .A1(n3740), .A2(n295), .ZN(n3882) );
  BUF_X1 U58 ( .A(n2151), .Z(n4230) );
  BUF_X1 U59 ( .A(n2151), .Z(n4231) );
  AOI21_X2 U62 ( .B1(n639), .B2(n996), .A(n209), .ZN(n890) );
  CLKBUF_X1 U63 ( .A(n2310), .Z(n4232) );
  NOR2_X1 U65 ( .A1(n2288), .A2(n2000), .ZN(n2310) );
  NOR2_X2 U68 ( .A1(n67), .A2(is_subrot_i), .ZN(n1181) );
  OAI211_X2 U71 ( .C1(n1041), .C2(n1458), .A(n1039), .B(n1040), .ZN(n1322) );
  CLKBUF_X1 U75 ( .A(n3672), .Z(n4365) );
  BUF_X1 U78 ( .A(n85), .Z(n4288) );
  NAND2_X1 U84 ( .A1(n1320), .A2(n2695), .ZN(n2288) );
  AND2_X1 U85 ( .A1(n4342), .A2(n4343), .ZN(n1458) );
  CLKBUF_X2 U87 ( .A(n679), .Z(n75) );
  CLKBUF_X2 U88 ( .A(n679), .Z(n76) );
  BUF_X1 U89 ( .A(n77), .Z(n169) );
  CLKBUF_X1 U91 ( .A(n2565), .Z(n4302) );
  CLKBUF_X2 U92 ( .A(n540), .Z(n83) );
  CLKBUF_X1 U94 ( .A(operand_b_i[17]), .Z(n4328) );
  CLKBUF_X2 U98 ( .A(operand_b_i[9]), .Z(n4195) );
  CLKBUF_X1 U100 ( .A(n3177), .Z(n4309) );
  CLKBUF_X1 U106 ( .A(n4060), .Z(n4305) );
  MUX2_X1 U109 ( .A(n2397), .B(n2414), .S(n91), .Z(n3999) );
  CLKBUF_X1 U117 ( .A(n2236), .Z(n4278) );
  BUF_X1 U120 ( .A(n2261), .Z(n4298) );
  AND2_X1 U125 ( .A1(n1404), .A2(n1403), .ZN(n4334) );
  OR2_X1 U127 ( .A1(n2288), .A2(n1933), .ZN(n2207) );
  BUF_X2 U129 ( .A(n1261), .Z(n1657) );
  BUF_X1 U132 ( .A(n2169), .Z(n1884) );
  OAI21_X1 U134 ( .B1(n175), .B2(n1600), .A(n1599), .ZN(n2120) );
  BUF_X2 U135 ( .A(n1261), .Z(n1730) );
  NAND2_X1 U137 ( .A1(n527), .A2(n526), .ZN(n4294) );
  OAI21_X1 U139 ( .B1(div_shift[1]), .B2(n299), .A(n297), .ZN(n527) );
  OR2_X1 U141 ( .A1(n3095), .A2(n1033), .ZN(n1461) );
  AND2_X1 U143 ( .A1(n3992), .A2(n1015), .ZN(n1018) );
  CLKBUF_X1 U150 ( .A(n1158), .Z(n4308) );
  NOR2_X1 U155 ( .A1(n3296), .A2(n4310), .ZN(n4364) );
  NAND4_X1 U157 ( .A1(n3079), .A2(n3499), .A3(n2582), .A4(n2563), .ZN(n278) );
  CLKBUF_X1 U160 ( .A(operand_a_i[31]), .Z(n4304) );
  CLKBUF_X1 U169 ( .A(operator_i[6]), .Z(n4306) );
  BUF_X2 U172 ( .A(operator_i[1]), .Z(n4337) );
  CLKBUF_X1 U173 ( .A(n3120), .Z(n60) );
  INV_X1 U182 ( .A(operand_b_i[28]), .ZN(n4335) );
  AND2_X1 U184 ( .A1(operand_a_i[28]), .A2(n4335), .ZN(n2531) );
  INV_X1 U185 ( .A(n918), .ZN(n1223) );
  AND2_X1 U188 ( .A1(operator_i[1]), .A2(n2648), .ZN(n386) );
  INV_X1 U189 ( .A(n386), .ZN(n3831) );
  OR2_X1 U206 ( .A1(n4327), .A2(n4325), .ZN(n1373) );
  AND2_X1 U209 ( .A1(n219), .A2(n398), .ZN(n3740) );
  CLKBUF_X1 U216 ( .A(operand_a_i[1]), .Z(n4225) );
  CLKBUF_X1 U219 ( .A(operand_a_i[8]), .Z(n149) );
  OAI22_X1 U229 ( .A1(n1545), .A2(n4115), .B1(n1544), .B2(n4127), .ZN(n1257)
         );
  INV_X1 U237 ( .A(n1545), .ZN(n1532) );
  INV_X1 U239 ( .A(n137), .ZN(n1011) );
  NAND2_X1 U242 ( .A1(n91), .A2(n3387), .ZN(n1594) );
  CLKBUF_X1 U244 ( .A(n2547), .Z(n4087) );
  INV_X1 U246 ( .A(bmask_b_i[3]), .ZN(n1109) );
  CLKBUF_X2 U249 ( .A(n3837), .Z(n3988) );
  INV_X1 U253 ( .A(n3889), .ZN(n3144) );
  CLKBUF_X1 U254 ( .A(operand_b_i[18]), .Z(n4194) );
  AND2_X2 U266 ( .A1(vector_mode_i[1]), .A2(vector_mode_i[0]), .ZN(n3387) );
  INV_X1 U268 ( .A(n1871), .ZN(n90) );
  AOI211_X1 U275 ( .C1(n4316), .C2(n4188), .A(n4187), .B(n4186), .ZN(n4190) );
  NAND4_X1 U284 ( .A1(n884), .A2(n883), .A3(n882), .A4(n881), .ZN(n3000) );
  OR2_X1 U285 ( .A1(n2280), .A2(n2279), .ZN(n4303) );
  CLKBUF_X1 U289 ( .A(n1894), .Z(n4292) );
  AND4_X1 U290 ( .A1(n4329), .A2(n460), .A3(n3968), .A4(n4236), .ZN(n244) );
  CLKBUF_X1 U308 ( .A(operand_b_i[26]), .Z(n170) );
  CLKBUF_X1 U309 ( .A(operand_b_i[24]), .Z(n4340) );
  INV_X1 U321 ( .A(n2150), .ZN(n4332) );
  INV_X1 U326 ( .A(n2207), .ZN(n2108) );
  OR2_X1 U341 ( .A1(n4310), .A2(n3534), .ZN(n4234) );
  INV_X2 U342 ( .A(n91), .ZN(n2376) );
  AND2_X1 U359 ( .A1(n1680), .A2(n92), .ZN(n4235) );
  INV_X1 U362 ( .A(n2149), .ZN(n4331) );
  NAND2_X1 U389 ( .A1(n3943), .A2(n246), .ZN(n4236) );
  AND2_X1 U395 ( .A1(n264), .A2(n2372), .ZN(n4237) );
  INV_X1 U401 ( .A(n2169), .ZN(n2290) );
  NOR2_X1 U427 ( .A1(n3172), .A2(n4238), .ZN(n4252) );
  NAND2_X1 U430 ( .A1(n3180), .A2(n4354), .ZN(n4238) );
  NAND3_X2 U435 ( .A1(n325), .A2(n326), .A3(n324), .ZN(n2132) );
  OAI211_X1 U436 ( .C1(n4285), .C2(n1919), .A(n1563), .B(n192), .ZN(n2184) );
  NAND2_X1 U437 ( .A1(n84), .A2(n4242), .ZN(n4239) );
  AND2_X1 U450 ( .A1(n4239), .A2(n4240), .ZN(result_o[28]) );
  OR2_X1 U480 ( .A1(n4241), .A2(n1142), .ZN(n4240) );
  INV_X1 U487 ( .A(n226), .ZN(n4241) );
  AND2_X1 U549 ( .A1(n4344), .A2(n226), .ZN(n4242) );
  NAND2_X1 U553 ( .A1(n3181), .A2(n3180), .ZN(n4243) );
  NOR2_X1 U559 ( .A1(n4244), .A2(n4245), .ZN(result_o[20]) );
  AND2_X1 U596 ( .A1(n3642), .A2(n4262), .ZN(n4244) );
  NOR2_X1 U606 ( .A1(n4261), .A2(n699), .ZN(n4245) );
  NAND2_X1 U615 ( .A1(n3642), .A2(n4249), .ZN(n4246) );
  AND2_X1 U617 ( .A1(n4246), .A2(n4247), .ZN(result_o[27]) );
  OR2_X1 U632 ( .A1(n4248), .A2(n2875), .ZN(n4247) );
  INV_X1 U638 ( .A(n2880), .ZN(n4248) );
  AND2_X1 U639 ( .A1(n4349), .A2(n2880), .ZN(n4249) );
  NAND2_X1 U640 ( .A1(n3642), .A2(n4252), .ZN(n4250) );
  AND2_X1 U648 ( .A1(n4250), .A2(n4251), .ZN(result_o[18]) );
  OR2_X1 U649 ( .A1(n4243), .A2(n3174), .ZN(n4251) );
  NOR2_X1 U651 ( .A1(n4253), .A2(n4254), .ZN(result_o[13]) );
  AND2_X1 U652 ( .A1(n3642), .A2(n4264), .ZN(n4253) );
  NOR2_X1 U656 ( .A1(n4263), .A2(n3591), .ZN(n4254) );
  NAND2_X1 U672 ( .A1(n3642), .A2(n4258), .ZN(n4255) );
  AND2_X1 U686 ( .A1(n4255), .A2(n4256), .ZN(result_o[19]) );
  OR2_X1 U687 ( .A1(n4257), .A2(n768), .ZN(n4256) );
  INV_X1 U692 ( .A(n3039), .ZN(n4257) );
  AND2_X1 U693 ( .A1(n4348), .A2(n3039), .ZN(n4258) );
  NOR2_X1 U720 ( .A1(n4259), .A2(n4260), .ZN(result_o[22]) );
  AND2_X1 U739 ( .A1(n84), .A2(n4270), .ZN(n4259) );
  NOR2_X1 U787 ( .A1(n4269), .A2(n839), .ZN(n4260) );
  INV_X1 U799 ( .A(n220), .ZN(n4261) );
  AND2_X1 U829 ( .A1(n4352), .A2(n220), .ZN(n4262) );
  INV_X1 U904 ( .A(n229), .ZN(n4263) );
  AND2_X1 U949 ( .A1(n183), .A2(n229), .ZN(n4264) );
  NAND2_X1 U976 ( .A1(n3642), .A2(n4268), .ZN(n4265) );
  AND2_X1 U979 ( .A1(n4265), .A2(n4266), .ZN(result_o[23]) );
  OR2_X1 U982 ( .A1(n4267), .A2(n855), .ZN(n4266) );
  INV_X1 U1001 ( .A(n2964), .ZN(n4267) );
  AND2_X1 U1022 ( .A1(n4351), .A2(n2964), .ZN(n4268) );
  INV_X1 U1049 ( .A(n40), .ZN(n4269) );
  AND2_X1 U1061 ( .A1(n4361), .A2(n40), .ZN(n4270) );
  AND4_X1 U1064 ( .A1(n250), .A2(n251), .A3(n249), .A4(n248), .ZN(n2382) );
  AND4_X2 U1102 ( .A1(n2381), .A2(n2382), .A3(n2384), .A4(n2383), .ZN(n4118)
         );
  AOI21_X1 U1126 ( .B1(n1445), .B2(n1018), .A(n1017), .ZN(n4271) );
  OAI211_X1 U1183 ( .C1(n2028), .C2(n1751), .A(n1405), .B(n4334), .ZN(n2294)
         );
  INV_X1 U1203 ( .A(n4285), .ZN(n4272) );
  NAND2_X2 U1232 ( .A1(n1788), .A2(n1619), .ZN(n1764) );
  AND2_X1 U1315 ( .A1(n3337), .A2(n1020), .ZN(n4273) );
  INV_X1 U1528 ( .A(n4273), .ZN(n1518) );
  NAND2_X1 U1544 ( .A1(n492), .A2(n482), .ZN(n4274) );
  NOR2_X1 U1665 ( .A1(n492), .A2(n491), .ZN(n3686) );
  NAND4_X1 U1666 ( .A1(n2088), .A2(n2087), .A3(n2086), .A4(n2085), .ZN(n4275)
         );
  NAND2_X1 U1667 ( .A1(n338), .A2(n336), .ZN(n4276) );
  MUX2_X1 U1670 ( .A(n2413), .B(n2398), .S(n91), .Z(n3280) );
  MUX2_X1 U1671 ( .A(n2413), .B(n2398), .S(n2376), .Z(n3672) );
  OAI211_X1 U1682 ( .C1(n1927), .C2(n4294), .A(n1748), .B(n1747), .ZN(n4277)
         );
  OR2_X1 U1697 ( .A1(n2017), .A2(n1702), .ZN(n2236) );
  INV_X1 U1730 ( .A(n2152), .ZN(n4333) );
  MUX2_X2 U1762 ( .A(n2399), .B(n2412), .S(n91), .Z(n3595) );
  INV_X1 U1763 ( .A(n1377), .ZN(n4326) );
  CLKBUF_X1 U1869 ( .A(n4013), .Z(n4279) );
  XNOR2_X1 U1875 ( .A(n1134), .B(n4280), .ZN(n2864) );
  AND2_X1 U1912 ( .A1(n1132), .A2(n1148), .ZN(n4280) );
  OAI21_X1 U1917 ( .B1(n2000), .B2(n1842), .A(n1784), .ZN(n4281) );
  INV_X1 U1920 ( .A(n1614), .ZN(n4282) );
  BUF_X2 U1921 ( .A(n1562), .Z(n1821) );
  CLKBUF_X1 U1924 ( .A(ff1_result[0]), .Z(n4283) );
  CLKBUF_X1 U1929 ( .A(n2401), .Z(n4284) );
  MUX2_X1 U1955 ( .A(n1842), .B(n2070), .S(n1933), .Z(n2227) );
  NAND2_X1 U1964 ( .A1(n4356), .A2(n4355), .ZN(n4285) );
  AND4_X2 U1984 ( .A1(n2381), .A2(n2382), .A3(n2384), .A4(n2383), .ZN(n4286)
         );
  INV_X1 U1985 ( .A(n1657), .ZN(n4355) );
  OR2_X1 U1987 ( .A1(n4286), .A2(n4323), .ZN(n4010) );
  INV_X1 U2128 ( .A(n2333), .ZN(n85) );
  NOR2_X1 U2166 ( .A1(n3350), .A2(n2642), .ZN(n4289) );
  NOR2_X1 U2178 ( .A1(n3350), .A2(n2642), .ZN(n4290) );
  OAI211_X1 U2183 ( .C1(n2289), .C2(n2288), .A(n2286), .B(n2287), .ZN(n2414)
         );
  MUX2_X1 U2283 ( .A(n2397), .B(n2414), .S(n2376), .Z(n4060) );
  INV_X1 U2411 ( .A(n1143), .ZN(n4291) );
  INV_X1 U2415 ( .A(n1143), .ZN(n1126) );
  OR2_X1 U2500 ( .A1(n646), .A2(n647), .ZN(n4293) );
  NAND2_X1 U2621 ( .A1(n527), .A2(n526), .ZN(n1788) );
  MUX2_X1 U2632 ( .A(n1935), .B(n1934), .S(n1933), .Z(n2188) );
  INV_X1 U2633 ( .A(n1788), .ZN(n4356) );
  OAI21_X1 U2696 ( .B1(n1162), .B2(n1161), .A(n1160), .ZN(n4295) );
  INV_X1 U2697 ( .A(n1274), .ZN(n4296) );
  INV_X1 U2731 ( .A(n966), .ZN(n4297) );
  BUF_X1 U2734 ( .A(n1143), .Z(n1162) );
  INV_X1 U2744 ( .A(n4230), .ZN(n2103) );
  NOR2_X1 U2944 ( .A1(n626), .A2(n625), .ZN(n950) );
  AOI21_X1 U2955 ( .B1(n452), .B2(n82), .A(n1310), .ZN(n2261) );
  AND2_X1 U2965 ( .A1(n3642), .A2(n4345), .ZN(n3213) );
  MUX2_X1 U2971 ( .A(n2261), .B(n2256), .S(n1657), .Z(n1824) );
  CLKBUF_X1 U3005 ( .A(n1258), .Z(n4299) );
  INV_X1 U3137 ( .A(n4098), .ZN(n4300) );
  OR2_X1 U3147 ( .A1(n1050), .A2(n1051), .ZN(n4301) );
  NOR2_X1 U3151 ( .A1(n2952), .A2(n1052), .ZN(n1359) );
  OAI211_X1 U3247 ( .C1(n2278), .C2(n2277), .A(n2283), .B(n4303), .ZN(n2284)
         );
  NAND2_X1 U3248 ( .A1(n1620), .A2(n2230), .ZN(n2178) );
  INV_X1 U3249 ( .A(n4117), .ZN(n4310) );
  INV_X1 U3288 ( .A(n4117), .ZN(n4009) );
  NAND2_X1 U3290 ( .A1(n1636), .A2(n4235), .ZN(n128) );
  CLKBUF_X1 U3291 ( .A(n3320), .Z(n4311) );
  CLKBUF_X1 U3375 ( .A(n2334), .Z(n4312) );
  CLKBUF_X1 U3377 ( .A(n2743), .Z(n2606) );
  CLKBUF_X1 U3378 ( .A(n1768), .Z(n4313) );
  INV_X1 U3423 ( .A(n1515), .ZN(n4314) );
  CLKBUF_X1 U3424 ( .A(n2636), .Z(n4315) );
  AOI21_X1 U3449 ( .B1(n1445), .B2(n1018), .A(n1017), .ZN(n1524) );
  BUF_X1 U3450 ( .A(n4189), .Z(n4316) );
  MUX2_X1 U3451 ( .A(n2390), .B(n2421), .S(n2376), .Z(n4189) );
  INV_X1 U3475 ( .A(n1322), .ZN(n1395) );
  AND2_X1 U3476 ( .A1(n2636), .A2(n1016), .ZN(n1017) );
  CLKBUF_X1 U3519 ( .A(operator_i[3]), .Z(n487) );
  NAND2_X1 U3520 ( .A1(n375), .A2(n4317), .ZN(n2586) );
  AND2_X1 U3548 ( .A1(n374), .A2(n2585), .ZN(n4317) );
  AND2_X1 U3549 ( .A1(n335), .A2(operator_i[4]), .ZN(n4353) );
  AND2_X1 U3592 ( .A1(n421), .A2(n425), .ZN(n1587) );
  NAND2_X1 U3593 ( .A1(n649), .A2(n888), .ZN(n651) );
  NAND2_X1 U3594 ( .A1(n4318), .A2(n3066), .ZN(n3072) );
  NAND2_X1 U3617 ( .A1(n84), .A2(n4319), .ZN(n4318) );
  OR2_X1 U3619 ( .A1(n3044), .A2(n4310), .ZN(n4319) );
  NAND4_X1 U3660 ( .A1(n4320), .A2(n2762), .A3(n2760), .A4(n2761), .ZN(
        comparison_result_o) );
  NAND2_X1 U3686 ( .A1(n2743), .A2(n2742), .ZN(n4320) );
  NAND2_X1 U3687 ( .A1(n4321), .A2(n3214), .ZN(n3256) );
  NAND2_X1 U3709 ( .A1(n3642), .A2(n4322), .ZN(n4321) );
  OR2_X1 U3710 ( .A1(n3230), .A2(n4310), .ZN(n4322) );
  INV_X1 U3815 ( .A(n4350), .ZN(n4323) );
  NAND3_X1 U3866 ( .A1(n2574), .A2(n2573), .A3(n2572), .ZN(n2578) );
  OAI211_X1 U4063 ( .C1(n2539), .C2(n2538), .A(n2537), .B(n2536), .ZN(n2540)
         );
  NAND3_X1 U4087 ( .A1(n4324), .A2(n256), .A3(n257), .ZN(n251) );
  NAND2_X1 U4113 ( .A1(n3889), .A2(n4237), .ZN(n4324) );
  MUX2_X1 U4114 ( .A(n2401), .B(n2410), .S(n2376), .Z(n3889) );
  MUX2_X2 U4153 ( .A(n2402), .B(n2409), .S(n91), .Z(n3217) );
  NAND2_X1 U4234 ( .A1(n407), .A2(n2072), .ZN(n2409) );
  NAND3_X1 U4235 ( .A1(n1682), .A2(n42), .A3(n1679), .ZN(n1859) );
  NAND2_X1 U4236 ( .A1(n1929), .A2(n1930), .ZN(n1931) );
  MUX2_X1 U4237 ( .A(n2194), .B(n2261), .S(n1657), .Z(n1929) );
  NAND4_X1 U4238 ( .A1(operator_i[1]), .A2(n4353), .A3(n2647), .A4(n2651), 
        .ZN(n2503) );
  INV_X1 U4239 ( .A(n1018), .ZN(n1451) );
  AND2_X1 U4240 ( .A1(n4326), .A2(n1322), .ZN(n4325) );
  INV_X1 U4241 ( .A(n1378), .ZN(n4327) );
  NAND2_X1 U4242 ( .A1(n2603), .A2(n2595), .ZN(n2596) );
  NAND2_X1 U4243 ( .A1(n285), .A2(n62), .ZN(n214) );
  AND2_X1 U4244 ( .A1(n3967), .A2(n3966), .ZN(n4329) );
  NAND4_X1 U4245 ( .A1(n4330), .A2(n252), .A3(n2361), .A4(n2360), .ZN(n249) );
  NAND2_X1 U4246 ( .A1(n3010), .A2(n2725), .ZN(n4330) );
  NAND2_X1 U4247 ( .A1(n542), .A2(n543), .ZN(n616) );
  NAND2_X1 U4248 ( .A1(n541), .A2(n465), .ZN(n542) );
  AOI22_X1 U4249 ( .A1(n4333), .A2(n2103), .B1(n4332), .B2(n4331), .ZN(n2168)
         );
  NAND2_X1 U4250 ( .A1(n4336), .A2(n2140), .ZN(n2407) );
  NAND2_X1 U4251 ( .A1(n2125), .A2(n2292), .ZN(n4336) );
  NAND3_X1 U4252 ( .A1(n129), .A2(n131), .A3(n4313), .ZN(n1909) );
  OR2_X1 U4253 ( .A1(n4286), .A2(n3938), .ZN(n3942) );
  NAND2_X1 U4254 ( .A1(n4338), .A2(n3105), .ZN(n3110) );
  NAND2_X1 U4255 ( .A1(n3642), .A2(n4339), .ZN(n4338) );
  OR2_X1 U4256 ( .A1(n3086), .A2(n4310), .ZN(n4339) );
  OR2_X1 U4257 ( .A1(n4286), .A2(n4364), .ZN(n4363) );
  NAND3_X1 U4258 ( .A1(n218), .A2(n66), .A3(n52), .ZN(n67) );
  NAND2_X1 U4259 ( .A1(n84), .A2(n4341), .ZN(n2765) );
  OR2_X1 U4260 ( .A1(n2822), .A2(n4310), .ZN(n4341) );
  NAND2_X1 U4261 ( .A1(n1025), .A2(n1443), .ZN(n4342) );
  INV_X1 U4262 ( .A(n1024), .ZN(n4343) );
  OR2_X1 U4263 ( .A1(n3861), .A2(n4310), .ZN(n4344) );
  OR2_X1 U4264 ( .A1(n3191), .A2(n4310), .ZN(n4345) );
  NAND2_X1 U4265 ( .A1(n4346), .A2(n3000), .ZN(n3006) );
  NAND2_X1 U4266 ( .A1(n3642), .A2(n4347), .ZN(n4346) );
  OR2_X1 U4267 ( .A1(n2980), .A2(n4310), .ZN(n4347) );
  OR2_X1 U4268 ( .A1(n3013), .A2(n4310), .ZN(n4348) );
  OR2_X1 U4269 ( .A1(n2858), .A2(n4310), .ZN(n4349) );
  OR2_X1 U4270 ( .A1(n4039), .A2(n4310), .ZN(n4350) );
  OR2_X1 U4271 ( .A1(n2921), .A2(n4310), .ZN(n4351) );
  OR2_X1 U4272 ( .A1(n3903), .A2(n4310), .ZN(n4352) );
  OR2_X1 U4273 ( .A1(n3155), .A2(n4310), .ZN(n4354) );
  NAND2_X1 U4274 ( .A1(n1321), .A2(n1756), .ZN(n1698) );
  NAND2_X1 U4275 ( .A1(n84), .A2(n4357), .ZN(n3257) );
  OR2_X1 U4276 ( .A1(n3262), .A2(n4310), .ZN(n4357) );
  NAND3_X1 U4277 ( .A1(n4358), .A2(n3316), .A3(n3317), .ZN(result_o[30]) );
  NAND2_X1 U4278 ( .A1(n4363), .A2(n3313), .ZN(n4358) );
  NAND2_X1 U4279 ( .A1(n4359), .A2(n3347), .ZN(n104) );
  NAND2_X1 U4280 ( .A1(n3642), .A2(n4360), .ZN(n4359) );
  OR2_X1 U4281 ( .A1(n3325), .A2(n4310), .ZN(n4360) );
  OR2_X1 U4282 ( .A1(n3111), .A2(n4310), .ZN(n4361) );
  AOI21_X1 U4283 ( .B1(n4362), .B2(n1059), .A(n1058), .ZN(n1270) );
  OAI211_X1 U4284 ( .C1(n1041), .C2(n1458), .A(n1039), .B(n1040), .ZN(n4362)
         );
  OAI21_X1 U4285 ( .B1(n930), .B2(n117), .A(n631), .ZN(n137) );
  NAND3_X1 U4286 ( .A1(n218), .A2(n66), .A3(n52), .ZN(n217) );
  AND2_X1 U4287 ( .A1(n84), .A2(n4234), .ZN(n4366) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_12 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_11 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_10 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_9 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_8 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_7 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_6 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_5 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_4 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_3 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_2 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_1 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_0 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module riscv_hwloop_regs_N_REGS2 ( clk, rst_n, hwlp_start_data_i, 
        hwlp_end_data_i, hwlp_cnt_data_i, hwlp_we_i, hwlp_regid_i, valid_i, 
        hwlp_dec_cnt_i, hwlp_start_addr_o, hwlp_end_addr_o, hwlp_counter_o );
  input [31:0] hwlp_start_data_i;
  input [31:0] hwlp_end_data_i;
  input [31:0] hwlp_cnt_data_i;
  input [2:0] hwlp_we_i;
  input [0:0] hwlp_regid_i;
  input [1:0] hwlp_dec_cnt_i;
  output [63:0] hwlp_start_addr_o;
  output [63:0] hwlp_end_addr_o;
  output [63:0] hwlp_counter_o;
  input clk, rst_n, valid_i;
  wire   n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n537, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n582, n583, n584,
         n585, n586, n587, n588, n589, n962, n964, n965, n967, n969, n971;

  INV_X1 U17 ( .A(hwlp_we_i[2]), .ZN(n1) );
  OR2_X1 U18 ( .A1(hwlp_counter_o[1]), .A2(hwlp_counter_o[0]), .ZN(n51) );
  INV_X1 U19 ( .A(n51), .ZN(n3) );
  NOR2_X1 U20 ( .A1(hwlp_counter_o[2]), .A2(hwlp_counter_o[3]), .ZN(n2) );
  NAND2_X1 U21 ( .A1(n3), .A2(n2), .ZN(n64) );
  INV_X1 U22 ( .A(n64), .ZN(n5) );
  NOR2_X1 U23 ( .A1(hwlp_counter_o[5]), .A2(hwlp_counter_o[4]), .ZN(n4) );
  NAND2_X1 U24 ( .A1(n5), .A2(n4), .ZN(n73) );
  OR2_X1 U25 ( .A1(hwlp_counter_o[7]), .A2(hwlp_counter_o[6]), .ZN(n6) );
  NOR2_X1 U26 ( .A1(n73), .A2(n6), .ZN(n79) );
  NOR2_X1 U27 ( .A1(hwlp_counter_o[9]), .A2(hwlp_counter_o[8]), .ZN(n7) );
  AND2_X1 U28 ( .A1(n79), .A2(n7), .ZN(n89) );
  NOR2_X1 U29 ( .A1(hwlp_counter_o[11]), .A2(hwlp_counter_o[10]), .ZN(n8) );
  NAND2_X1 U30 ( .A1(n89), .A2(n8), .ZN(n98) );
  OR2_X1 U31 ( .A1(hwlp_counter_o[13]), .A2(hwlp_counter_o[12]), .ZN(n9) );
  NOR2_X1 U32 ( .A1(n98), .A2(n9), .ZN(n107) );
  NOR2_X1 U33 ( .A1(hwlp_counter_o[15]), .A2(hwlp_counter_o[14]), .ZN(n10) );
  NAND2_X1 U34 ( .A1(n107), .A2(n10), .ZN(n117) );
  OR2_X1 U35 ( .A1(hwlp_counter_o[17]), .A2(hwlp_counter_o[16]), .ZN(n11) );
  NOR2_X1 U36 ( .A1(n117), .A2(n11), .ZN(n125) );
  NOR2_X1 U37 ( .A1(hwlp_counter_o[19]), .A2(hwlp_counter_o[18]), .ZN(n12) );
  AND2_X1 U38 ( .A1(n125), .A2(n12), .ZN(n134) );
  NOR2_X1 U39 ( .A1(hwlp_counter_o[21]), .A2(hwlp_counter_o[20]), .ZN(n13) );
  AND2_X1 U40 ( .A1(n134), .A2(n13), .ZN(n143) );
  NOR2_X1 U41 ( .A1(hwlp_counter_o[23]), .A2(hwlp_counter_o[22]), .ZN(n14) );
  AND2_X1 U42 ( .A1(n143), .A2(n14), .ZN(n344) );
  NOR2_X1 U43 ( .A1(hwlp_counter_o[25]), .A2(hwlp_counter_o[24]), .ZN(n15) );
  AND2_X1 U44 ( .A1(n344), .A2(n15), .ZN(n353) );
  NOR2_X1 U45 ( .A1(hwlp_counter_o[27]), .A2(hwlp_counter_o[26]), .ZN(n16) );
  AND2_X1 U46 ( .A1(n353), .A2(n16), .ZN(n361) );
  INV_X1 U47 ( .A(n361), .ZN(n18) );
  AND2_X1 U48 ( .A1(valid_i), .A2(hwlp_dec_cnt_i[0]), .ZN(n48) );
  OR2_X1 U49 ( .A1(n378), .A2(n48), .ZN(n372) );
  INV_X1 U50 ( .A(n372), .ZN(n354) );
  AOI21_X1 U51 ( .B1(n17), .B2(n18), .A(n354), .ZN(n365) );
  NAND2_X1 U52 ( .A1(n361), .A2(n548), .ZN(n371) );
  OR2_X1 U53 ( .A1(n366), .A2(n371), .ZN(n367) );
  OAI21_X1 U54 ( .B1(n365), .B2(n548), .A(n367), .ZN(n19) );
  OR2_X1 U57 ( .A1(hwlp_counter_o[33]), .A2(hwlp_counter_o[32]), .ZN(n390) );
  INV_X1 U58 ( .A(n390), .ZN(n22) );
  NOR2_X1 U59 ( .A1(hwlp_counter_o[34]), .A2(hwlp_counter_o[35]), .ZN(n21) );
  NAND2_X1 U60 ( .A1(n22), .A2(n21), .ZN(n403) );
  INV_X1 U61 ( .A(n403), .ZN(n24) );
  NOR2_X1 U62 ( .A1(hwlp_counter_o[37]), .A2(hwlp_counter_o[36]), .ZN(n23) );
  NAND2_X1 U63 ( .A1(n24), .A2(n23), .ZN(n412) );
  OR2_X1 U64 ( .A1(hwlp_counter_o[39]), .A2(hwlp_counter_o[38]), .ZN(n25) );
  NOR2_X1 U65 ( .A1(n412), .A2(n25), .ZN(n418) );
  NOR2_X1 U66 ( .A1(hwlp_counter_o[41]), .A2(hwlp_counter_o[40]), .ZN(n26) );
  AND2_X1 U67 ( .A1(n418), .A2(n26), .ZN(n428) );
  NOR2_X1 U68 ( .A1(hwlp_counter_o[43]), .A2(hwlp_counter_o[42]), .ZN(n27) );
  NAND2_X1 U69 ( .A1(n428), .A2(n27), .ZN(n437) );
  OR2_X1 U70 ( .A1(hwlp_counter_o[45]), .A2(hwlp_counter_o[44]), .ZN(n28) );
  NOR2_X1 U71 ( .A1(n437), .A2(n28), .ZN(n447) );
  NOR2_X1 U72 ( .A1(hwlp_counter_o[47]), .A2(hwlp_counter_o[46]), .ZN(n29) );
  NAND2_X1 U73 ( .A1(n447), .A2(n29), .ZN(n457) );
  OR2_X1 U74 ( .A1(hwlp_counter_o[49]), .A2(hwlp_counter_o[48]), .ZN(n30) );
  NOR2_X1 U75 ( .A1(n457), .A2(n30), .ZN(n465) );
  NOR2_X1 U76 ( .A1(hwlp_counter_o[51]), .A2(hwlp_counter_o[50]), .ZN(n31) );
  AND2_X1 U77 ( .A1(n465), .A2(n31), .ZN(n474) );
  NOR2_X1 U78 ( .A1(hwlp_counter_o[53]), .A2(hwlp_counter_o[52]), .ZN(n32) );
  AND2_X1 U79 ( .A1(n474), .A2(n32), .ZN(n483) );
  NOR2_X1 U80 ( .A1(hwlp_counter_o[55]), .A2(hwlp_counter_o[54]), .ZN(n33) );
  AND2_X1 U81 ( .A1(n483), .A2(n33), .ZN(n492) );
  NOR2_X1 U82 ( .A1(hwlp_counter_o[57]), .A2(hwlp_counter_o[56]), .ZN(n34) );
  AND2_X1 U83 ( .A1(n492), .A2(n34), .ZN(n501) );
  NOR2_X1 U84 ( .A1(hwlp_counter_o[59]), .A2(hwlp_counter_o[58]), .ZN(n35) );
  AND2_X1 U85 ( .A1(n501), .A2(n35), .ZN(n509) );
  INV_X1 U86 ( .A(n509), .ZN(n37) );
  NAND2_X1 U87 ( .A1(valid_i), .A2(hwlp_dec_cnt_i[1]), .ZN(n388) );
  NAND2_X1 U88 ( .A1(n36), .A2(n388), .ZN(n520) );
  INV_X1 U89 ( .A(n520), .ZN(n502) );
  AOI21_X1 U90 ( .B1(n36), .B2(n37), .A(n502), .ZN(n513) );
  NAND2_X1 U91 ( .A1(n520), .A2(n36), .ZN(n514) );
  NAND2_X1 U92 ( .A1(n509), .A2(n549), .ZN(n519) );
  OR2_X1 U93 ( .A1(n514), .A2(n519), .ZN(n515) );
  OAI21_X1 U94 ( .B1(n513), .B2(n549), .A(n515), .ZN(n38) );
  OAI21_X1 U97 ( .B1(n360), .B2(n79), .A(n372), .ZN(n86) );
  AOI21_X1 U98 ( .B1(hwlp_counter_o[8]), .B2(n17), .A(n86), .ZN(n40) );
  NAND2_X1 U99 ( .A1(n381), .A2(n89), .ZN(n91) );
  OAI21_X1 U100 ( .B1(n40), .B2(n573), .A(n91), .ZN(n41) );
  AOI21_X1 U101 ( .B1(hwlp_cnt_data_i[9]), .B2(n360), .A(n41), .ZN(n42) );
  INV_X1 U102 ( .A(n42), .ZN(n168) );
  OAI21_X1 U103 ( .B1(n508), .B2(n418), .A(n520), .ZN(n425) );
  AOI21_X1 U104 ( .B1(hwlp_counter_o[40]), .B2(n36), .A(n425), .ZN(n43) );
  NAND2_X1 U106 ( .A1(n528), .A2(n428), .ZN(n430) );
  OAI21_X1 U107 ( .B1(n43), .B2(n574), .A(n430), .ZN(n44) );
  AOI21_X1 U108 ( .B1(hwlp_cnt_data_i[9]), .B2(n508), .A(n44), .ZN(n45) );
  INV_X1 U109 ( .A(n45), .ZN(n200) );
  NAND2_X1 U110 ( .A1(hwlp_cnt_data_i[0]), .A2(n575), .ZN(n47) );
  MUX2_X1 U111 ( .A(n366), .B(n372), .S(hwlp_counter_o[0]), .Z(n46) );
  NAND2_X1 U112 ( .A1(n47), .A2(n46), .ZN(n177) );
  NAND2_X1 U113 ( .A1(hwlp_cnt_data_i[1]), .A2(n360), .ZN(n53) );
  INV_X1 U114 ( .A(n48), .ZN(n49) );
  NOR2_X1 U115 ( .A1(n49), .A2(hwlp_counter_o[0]), .ZN(n50) );
  NOR2_X1 U116 ( .A1(n360), .A2(n50), .ZN(n54) );
  NOR2_X1 U117 ( .A1(n366), .A2(n51), .ZN(n56) );
  AOI21_X1 U118 ( .B1(hwlp_counter_o[1]), .B2(n54), .A(n56), .ZN(n52) );
  NAND2_X1 U119 ( .A1(n53), .A2(n52), .ZN(n176) );
  NAND2_X1 U120 ( .A1(hwlp_cnt_data_i[2]), .A2(n360), .ZN(n59) );
  INV_X1 U121 ( .A(n54), .ZN(n55) );
  OAI21_X1 U122 ( .B1(n366), .B2(n572), .A(n55), .ZN(n61) );
  AND2_X1 U123 ( .A1(n56), .A2(n542), .ZN(n57) );
  AOI21_X1 U124 ( .B1(hwlp_counter_o[2]), .B2(n61), .A(n57), .ZN(n58) );
  NAND2_X1 U125 ( .A1(n59), .A2(n58), .ZN(n175) );
  NAND2_X1 U126 ( .A1(hwlp_cnt_data_i[3]), .A2(n360), .ZN(n63) );
  OAI21_X1 U127 ( .B1(n542), .B2(n570), .A(n64), .ZN(n60) );
  AOI22_X1 U128 ( .A1(n61), .A2(hwlp_counter_o[3]), .B1(n381), .B2(n60), .ZN(
        n62) );
  NAND2_X1 U129 ( .A1(n63), .A2(n62), .ZN(n174) );
  NAND2_X1 U130 ( .A1(hwlp_cnt_data_i[4]), .A2(n360), .ZN(n68) );
  AOI21_X1 U131 ( .B1(n17), .B2(n64), .A(n354), .ZN(n69) );
  INV_X1 U132 ( .A(n69), .ZN(n66) );
  NOR3_X1 U133 ( .A1(n366), .A2(hwlp_counter_o[4]), .A3(n64), .ZN(n65) );
  AOI21_X1 U134 ( .B1(n66), .B2(hwlp_counter_o[4]), .A(n65), .ZN(n67) );
  NAND2_X1 U135 ( .A1(n68), .A2(n67), .ZN(n173) );
  NAND2_X1 U136 ( .A1(hwlp_cnt_data_i[5]), .A2(n575), .ZN(n72) );
  OAI21_X1 U137 ( .B1(n360), .B2(n550), .A(n69), .ZN(n70) );
  NOR2_X1 U138 ( .A1(n366), .A2(n73), .ZN(n75) );
  AOI21_X1 U139 ( .B1(n70), .B2(hwlp_counter_o[5]), .A(n75), .ZN(n71) );
  NAND2_X1 U140 ( .A1(n72), .A2(n71), .ZN(n172) );
  NAND2_X1 U141 ( .A1(hwlp_cnt_data_i[6]), .A2(n360), .ZN(n77) );
  AOI21_X1 U142 ( .B1(n17), .B2(n73), .A(n354), .ZN(n78) );
  NOR2_X1 U143 ( .A1(n78), .A2(n544), .ZN(n74) );
  AOI21_X1 U144 ( .B1(n75), .B2(n544), .A(n74), .ZN(n76) );
  NAND2_X1 U145 ( .A1(n77), .A2(n76), .ZN(n171) );
  NAND2_X1 U146 ( .A1(hwlp_cnt_data_i[7]), .A2(n360), .ZN(n83) );
  OAI21_X1 U147 ( .B1(n360), .B2(n544), .A(n78), .ZN(n81) );
  NAND2_X1 U148 ( .A1(n381), .A2(n79), .ZN(n84) );
  INV_X1 U149 ( .A(n84), .ZN(n80) );
  AOI21_X1 U150 ( .B1(hwlp_counter_o[7]), .B2(n81), .A(n80), .ZN(n82) );
  NAND2_X1 U151 ( .A1(n83), .A2(n82), .ZN(n170) );
  NAND2_X1 U152 ( .A1(hwlp_cnt_data_i[8]), .A2(n360), .ZN(n88) );
  NOR2_X1 U153 ( .A1(n84), .A2(hwlp_counter_o[8]), .ZN(n85) );
  AOI21_X1 U154 ( .B1(hwlp_counter_o[8]), .B2(n86), .A(n85), .ZN(n87) );
  NAND2_X1 U155 ( .A1(n88), .A2(n87), .ZN(n169) );
  NAND2_X1 U156 ( .A1(hwlp_cnt_data_i[10]), .A2(n575), .ZN(n93) );
  INV_X1 U157 ( .A(n89), .ZN(n90) );
  AOI21_X1 U158 ( .B1(n17), .B2(n90), .A(n354), .ZN(n94) );
  MUX2_X1 U159 ( .A(n91), .B(n94), .S(hwlp_counter_o[10]), .Z(n92) );
  NAND2_X1 U160 ( .A1(n93), .A2(n92), .ZN(n167) );
  NAND2_X1 U161 ( .A1(hwlp_cnt_data_i[11]), .A2(n575), .ZN(n97) );
  OAI21_X1 U162 ( .B1(n360), .B2(n554), .A(n94), .ZN(n95) );
  NOR2_X1 U163 ( .A1(n366), .A2(n98), .ZN(n100) );
  AOI21_X1 U164 ( .B1(n95), .B2(hwlp_counter_o[11]), .A(n100), .ZN(n96) );
  NAND2_X1 U165 ( .A1(n97), .A2(n96), .ZN(n166) );
  NAND2_X1 U166 ( .A1(hwlp_cnt_data_i[12]), .A2(n360), .ZN(n102) );
  AOI21_X1 U167 ( .B1(n17), .B2(n98), .A(n354), .ZN(n103) );
  NOR2_X1 U168 ( .A1(n103), .A2(n546), .ZN(n99) );
  AOI21_X1 U169 ( .B1(n100), .B2(n546), .A(n99), .ZN(n101) );
  NAND2_X1 U170 ( .A1(n102), .A2(n101), .ZN(n165) );
  NAND2_X1 U171 ( .A1(hwlp_cnt_data_i[13]), .A2(n360), .ZN(n106) );
  NAND2_X1 U172 ( .A1(n381), .A2(n107), .ZN(n109) );
  OAI21_X1 U173 ( .B1(n378), .B2(n546), .A(n103), .ZN(n104) );
  NAND2_X1 U174 ( .A1(n104), .A2(hwlp_counter_o[13]), .ZN(n105) );
  NAND3_X1 U175 ( .A1(n106), .A2(n109), .A3(n105), .ZN(n164) );
  NAND2_X1 U176 ( .A1(hwlp_cnt_data_i[14]), .A2(n575), .ZN(n111) );
  INV_X1 U177 ( .A(n107), .ZN(n108) );
  AOI21_X1 U178 ( .B1(n17), .B2(n108), .A(n354), .ZN(n113) );
  MUX2_X1 U179 ( .A(n109), .B(n113), .S(hwlp_counter_o[14]), .Z(n110) );
  NAND2_X1 U180 ( .A1(n111), .A2(n110), .ZN(n163) );
  NAND2_X1 U181 ( .A1(hwlp_cnt_data_i[15]), .A2(n360), .ZN(n116) );
  INV_X1 U182 ( .A(n117), .ZN(n112) );
  NAND2_X1 U183 ( .A1(n381), .A2(n112), .ZN(n118) );
  OAI21_X1 U184 ( .B1(n360), .B2(n566), .A(n113), .ZN(n114) );
  NAND2_X1 U185 ( .A1(n114), .A2(hwlp_counter_o[15]), .ZN(n115) );
  NAND3_X1 U186 ( .A1(n116), .A2(n118), .A3(n115), .ZN(n162) );
  NAND2_X1 U187 ( .A1(hwlp_cnt_data_i[16]), .A2(n575), .ZN(n120) );
  AOI21_X1 U188 ( .B1(n17), .B2(n117), .A(n354), .ZN(n121) );
  MUX2_X1 U189 ( .A(n118), .B(n121), .S(hwlp_counter_o[16]), .Z(n119) );
  NAND2_X1 U190 ( .A1(n120), .A2(n119), .ZN(n161) );
  NAND2_X1 U191 ( .A1(hwlp_cnt_data_i[17]), .A2(n575), .ZN(n124) );
  NAND2_X1 U192 ( .A1(n381), .A2(n125), .ZN(n127) );
  OAI21_X1 U193 ( .B1(n575), .B2(n563), .A(n121), .ZN(n122) );
  NAND2_X1 U194 ( .A1(n122), .A2(hwlp_counter_o[17]), .ZN(n123) );
  NAND3_X1 U195 ( .A1(n124), .A2(n127), .A3(n123), .ZN(n160) );
  NAND2_X1 U196 ( .A1(hwlp_cnt_data_i[18]), .A2(n575), .ZN(n129) );
  INV_X1 U197 ( .A(n125), .ZN(n126) );
  AOI21_X1 U198 ( .B1(n17), .B2(n126), .A(n354), .ZN(n130) );
  MUX2_X1 U199 ( .A(n127), .B(n130), .S(hwlp_counter_o[18]), .Z(n128) );
  NAND2_X1 U200 ( .A1(n129), .A2(n128), .ZN(n159) );
  NAND2_X1 U201 ( .A1(hwlp_cnt_data_i[19]), .A2(n575), .ZN(n133) );
  NAND2_X1 U202 ( .A1(n381), .A2(n134), .ZN(n136) );
  OAI21_X1 U203 ( .B1(n360), .B2(n557), .A(n130), .ZN(n131) );
  NAND2_X1 U204 ( .A1(n131), .A2(hwlp_counter_o[19]), .ZN(n132) );
  NAND3_X1 U205 ( .A1(n133), .A2(n136), .A3(n132), .ZN(n158) );
  NAND2_X1 U206 ( .A1(hwlp_cnt_data_i[20]), .A2(n575), .ZN(n138) );
  INV_X1 U207 ( .A(n134), .ZN(n135) );
  AOI21_X1 U208 ( .B1(n17), .B2(n135), .A(n354), .ZN(n139) );
  MUX2_X1 U209 ( .A(n136), .B(n139), .S(hwlp_counter_o[20]), .Z(n137) );
  NAND2_X1 U210 ( .A1(n138), .A2(n137), .ZN(n157) );
  NAND2_X1 U211 ( .A1(hwlp_cnt_data_i[21]), .A2(n575), .ZN(n142) );
  NAND2_X1 U212 ( .A1(n381), .A2(n143), .ZN(n145) );
  OAI21_X1 U213 ( .B1(n360), .B2(n562), .A(n139), .ZN(n140) );
  NAND2_X1 U214 ( .A1(n140), .A2(hwlp_counter_o[21]), .ZN(n141) );
  NAND3_X1 U215 ( .A1(n142), .A2(n145), .A3(n141), .ZN(n156) );
  NAND2_X1 U216 ( .A1(hwlp_cnt_data_i[22]), .A2(n575), .ZN(n339) );
  INV_X1 U217 ( .A(n143), .ZN(n144) );
  AOI21_X1 U218 ( .B1(n17), .B2(n144), .A(n354), .ZN(n340) );
  MUX2_X1 U219 ( .A(n145), .B(n340), .S(hwlp_counter_o[22]), .Z(n338) );
  NAND2_X1 U220 ( .A1(n339), .A2(n338), .ZN(n155) );
  NAND2_X1 U221 ( .A1(hwlp_cnt_data_i[23]), .A2(n575), .ZN(n343) );
  NAND2_X1 U222 ( .A1(n381), .A2(n344), .ZN(n346) );
  OAI21_X1 U223 ( .B1(n360), .B2(n567), .A(n340), .ZN(n341) );
  NAND2_X1 U224 ( .A1(n341), .A2(hwlp_counter_o[23]), .ZN(n342) );
  NAND3_X1 U225 ( .A1(n343), .A2(n346), .A3(n342), .ZN(n154) );
  NAND2_X1 U226 ( .A1(hwlp_cnt_data_i[24]), .A2(n575), .ZN(n348) );
  INV_X1 U227 ( .A(n344), .ZN(n345) );
  AOI21_X1 U228 ( .B1(n17), .B2(n345), .A(n354), .ZN(n349) );
  MUX2_X1 U229 ( .A(n346), .B(n349), .S(hwlp_counter_o[24]), .Z(n347) );
  NAND2_X1 U230 ( .A1(n348), .A2(n347), .ZN(n153) );
  NAND2_X1 U231 ( .A1(hwlp_cnt_data_i[25]), .A2(n575), .ZN(n352) );
  NAND2_X1 U232 ( .A1(n381), .A2(n353), .ZN(n356) );
  OAI21_X1 U233 ( .B1(n360), .B2(n560), .A(n349), .ZN(n350) );
  NAND2_X1 U234 ( .A1(n350), .A2(hwlp_counter_o[25]), .ZN(n351) );
  NAND3_X1 U235 ( .A1(n352), .A2(n356), .A3(n351), .ZN(n152) );
  NAND2_X1 U236 ( .A1(hwlp_cnt_data_i[26]), .A2(n575), .ZN(n358) );
  INV_X1 U237 ( .A(n353), .ZN(n355) );
  AOI21_X1 U238 ( .B1(n17), .B2(n355), .A(n354), .ZN(n359) );
  MUX2_X1 U239 ( .A(n356), .B(n359), .S(hwlp_counter_o[26]), .Z(n357) );
  NAND2_X1 U240 ( .A1(n358), .A2(n357), .ZN(n151) );
  NAND2_X1 U241 ( .A1(hwlp_cnt_data_i[27]), .A2(n575), .ZN(n364) );
  OAI21_X1 U242 ( .B1(n360), .B2(n558), .A(n359), .ZN(n362) );
  AOI22_X1 U243 ( .A1(n362), .A2(hwlp_counter_o[27]), .B1(n381), .B2(n361), 
        .ZN(n363) );
  NAND2_X1 U244 ( .A1(n364), .A2(n363), .ZN(n150) );
  NAND2_X1 U245 ( .A1(hwlp_cnt_data_i[29]), .A2(n575), .ZN(n370) );
  OAI21_X1 U246 ( .B1(n366), .B2(n548), .A(n365), .ZN(n368) );
  NOR2_X1 U247 ( .A1(n367), .A2(hwlp_counter_o[29]), .ZN(n374) );
  AOI21_X1 U248 ( .B1(hwlp_counter_o[29]), .B2(n368), .A(n374), .ZN(n369) );
  NAND2_X1 U249 ( .A1(n370), .A2(n369), .ZN(n148) );
  NAND2_X1 U250 ( .A1(hwlp_cnt_data_i[30]), .A2(n575), .ZN(n377) );
  OAI21_X1 U251 ( .B1(hwlp_counter_o[29]), .B2(n371), .A(n381), .ZN(n373) );
  NAND2_X1 U252 ( .A1(n373), .A2(n372), .ZN(n380) );
  INV_X1 U253 ( .A(n374), .ZN(n375) );
  NOR2_X1 U254 ( .A1(n375), .A2(hwlp_counter_o[30]), .ZN(n379) );
  AOI21_X1 U255 ( .B1(hwlp_counter_o[30]), .B2(n380), .A(n379), .ZN(n376) );
  NAND2_X1 U256 ( .A1(n377), .A2(n376), .ZN(n147) );
  NAND2_X1 U257 ( .A1(hwlp_cnt_data_i[31]), .A2(n575), .ZN(n385) );
  INV_X1 U258 ( .A(n379), .ZN(n383) );
  AOI21_X1 U259 ( .B1(n381), .B2(hwlp_counter_o[30]), .A(n380), .ZN(n382) );
  MUX2_X1 U260 ( .A(n383), .B(n382), .S(hwlp_counter_o[31]), .Z(n384) );
  NAND2_X1 U261 ( .A1(n385), .A2(n384), .ZN(n146) );
  NAND2_X1 U262 ( .A1(hwlp_cnt_data_i[0]), .A2(n446), .ZN(n387) );
  MUX2_X1 U263 ( .A(n514), .B(n520), .S(hwlp_counter_o[32]), .Z(n386) );
  NAND2_X1 U264 ( .A1(n387), .A2(n386), .ZN(n209) );
  NAND2_X1 U265 ( .A1(hwlp_cnt_data_i[1]), .A2(n446), .ZN(n392) );
  INV_X1 U266 ( .A(n388), .ZN(n389) );
  AOI21_X1 U267 ( .B1(n389), .B2(n552), .A(n508), .ZN(n393) );
  NOR2_X1 U268 ( .A1(n514), .A2(n390), .ZN(n395) );
  AOI21_X1 U269 ( .B1(hwlp_counter_o[33]), .B2(n393), .A(n395), .ZN(n391) );
  NAND2_X1 U270 ( .A1(n392), .A2(n391), .ZN(n208) );
  NAND2_X1 U271 ( .A1(hwlp_cnt_data_i[2]), .A2(n446), .ZN(n398) );
  INV_X1 U272 ( .A(n393), .ZN(n394) );
  OAI21_X1 U273 ( .B1(n561), .B2(n514), .A(n394), .ZN(n400) );
  AND2_X1 U274 ( .A1(n395), .A2(n543), .ZN(n396) );
  AOI21_X1 U275 ( .B1(hwlp_counter_o[34]), .B2(n400), .A(n396), .ZN(n397) );
  NAND2_X1 U276 ( .A1(n398), .A2(n397), .ZN(n207) );
  NAND2_X1 U277 ( .A1(hwlp_cnt_data_i[3]), .A2(n446), .ZN(n402) );
  OAI21_X1 U278 ( .B1(n543), .B2(n571), .A(n403), .ZN(n399) );
  AOI22_X1 U279 ( .A1(n400), .A2(hwlp_counter_o[35]), .B1(n528), .B2(n399), 
        .ZN(n401) );
  NAND2_X1 U280 ( .A1(n402), .A2(n401), .ZN(n206) );
  NAND2_X1 U281 ( .A1(hwlp_cnt_data_i[4]), .A2(n446), .ZN(n407) );
  AOI21_X1 U282 ( .B1(n36), .B2(n403), .A(n502), .ZN(n408) );
  INV_X1 U283 ( .A(n408), .ZN(n405) );
  NOR3_X1 U284 ( .A1(n514), .A2(hwlp_counter_o[36]), .A3(n403), .ZN(n404) );
  AOI21_X1 U285 ( .B1(n405), .B2(hwlp_counter_o[36]), .A(n404), .ZN(n406) );
  NAND2_X1 U286 ( .A1(n407), .A2(n406), .ZN(n205) );
  NAND2_X1 U287 ( .A1(hwlp_cnt_data_i[5]), .A2(n446), .ZN(n411) );
  OAI21_X1 U288 ( .B1(n508), .B2(n551), .A(n408), .ZN(n409) );
  NOR2_X1 U289 ( .A1(n514), .A2(n412), .ZN(n414) );
  AOI21_X1 U290 ( .B1(n409), .B2(hwlp_counter_o[37]), .A(n414), .ZN(n410) );
  NAND2_X1 U291 ( .A1(n411), .A2(n410), .ZN(n204) );
  NAND2_X1 U292 ( .A1(hwlp_cnt_data_i[6]), .A2(n446), .ZN(n416) );
  AOI21_X1 U293 ( .B1(n36), .B2(n412), .A(n502), .ZN(n417) );
  NOR2_X1 U294 ( .A1(n417), .A2(n545), .ZN(n413) );
  AOI21_X1 U295 ( .B1(n414), .B2(n545), .A(n413), .ZN(n415) );
  NAND2_X1 U296 ( .A1(n416), .A2(n415), .ZN(n203) );
  NAND2_X1 U297 ( .A1(hwlp_cnt_data_i[7]), .A2(n446), .ZN(n422) );
  OAI21_X1 U298 ( .B1(n508), .B2(n545), .A(n417), .ZN(n420) );
  NAND2_X1 U299 ( .A1(n528), .A2(n418), .ZN(n423) );
  INV_X1 U300 ( .A(n423), .ZN(n419) );
  AOI21_X1 U301 ( .B1(hwlp_counter_o[39]), .B2(n420), .A(n419), .ZN(n421) );
  NAND2_X1 U302 ( .A1(n422), .A2(n421), .ZN(n202) );
  NAND2_X1 U303 ( .A1(hwlp_cnt_data_i[8]), .A2(n446), .ZN(n427) );
  NOR2_X1 U304 ( .A1(n423), .A2(hwlp_counter_o[40]), .ZN(n424) );
  AOI21_X1 U305 ( .B1(hwlp_counter_o[40]), .B2(n425), .A(n424), .ZN(n426) );
  NAND2_X1 U306 ( .A1(n427), .A2(n426), .ZN(n201) );
  NAND2_X1 U307 ( .A1(hwlp_cnt_data_i[10]), .A2(n446), .ZN(n432) );
  INV_X1 U308 ( .A(n428), .ZN(n429) );
  AOI21_X1 U309 ( .B1(n36), .B2(n429), .A(n502), .ZN(n433) );
  MUX2_X1 U310 ( .A(n430), .B(n433), .S(hwlp_counter_o[42]), .Z(n431) );
  NAND2_X1 U311 ( .A1(n432), .A2(n431), .ZN(n199) );
  NAND2_X1 U312 ( .A1(hwlp_cnt_data_i[11]), .A2(n446), .ZN(n436) );
  OAI21_X1 U313 ( .B1(n508), .B2(n555), .A(n433), .ZN(n434) );
  NOR2_X1 U314 ( .A1(n514), .A2(n437), .ZN(n439) );
  AOI21_X1 U315 ( .B1(n434), .B2(hwlp_counter_o[43]), .A(n439), .ZN(n435) );
  NAND2_X1 U316 ( .A1(n436), .A2(n435), .ZN(n198) );
  NAND2_X1 U317 ( .A1(hwlp_cnt_data_i[12]), .A2(n446), .ZN(n441) );
  AOI21_X1 U318 ( .B1(n36), .B2(n437), .A(n502), .ZN(n442) );
  NOR2_X1 U319 ( .A1(n442), .A2(n547), .ZN(n438) );
  AOI21_X1 U320 ( .B1(n439), .B2(n547), .A(n438), .ZN(n440) );
  NAND2_X1 U321 ( .A1(n441), .A2(n440), .ZN(n197) );
  NAND2_X1 U322 ( .A1(hwlp_cnt_data_i[13]), .A2(n446), .ZN(n445) );
  NAND2_X1 U323 ( .A1(n528), .A2(n447), .ZN(n449) );
  OAI21_X1 U324 ( .B1(n446), .B2(n547), .A(n442), .ZN(n443) );
  NAND2_X1 U325 ( .A1(n443), .A2(hwlp_counter_o[45]), .ZN(n444) );
  NAND3_X1 U326 ( .A1(n445), .A2(n449), .A3(n444), .ZN(n196) );
  NAND2_X1 U327 ( .A1(hwlp_cnt_data_i[14]), .A2(n446), .ZN(n451) );
  INV_X1 U328 ( .A(n447), .ZN(n448) );
  AOI21_X1 U329 ( .B1(n36), .B2(n448), .A(n502), .ZN(n453) );
  MUX2_X1 U330 ( .A(n449), .B(n453), .S(hwlp_counter_o[46]), .Z(n450) );
  NAND2_X1 U331 ( .A1(n451), .A2(n450), .ZN(n195) );
  NAND2_X1 U332 ( .A1(hwlp_cnt_data_i[15]), .A2(n446), .ZN(n456) );
  INV_X1 U333 ( .A(n457), .ZN(n452) );
  NAND2_X1 U334 ( .A1(n528), .A2(n452), .ZN(n458) );
  OAI21_X1 U335 ( .B1(n508), .B2(n568), .A(n453), .ZN(n454) );
  NAND2_X1 U336 ( .A1(n454), .A2(hwlp_counter_o[47]), .ZN(n455) );
  NAND3_X1 U337 ( .A1(n456), .A2(n458), .A3(n455), .ZN(n194) );
  NAND2_X1 U338 ( .A1(hwlp_cnt_data_i[16]), .A2(n446), .ZN(n460) );
  AOI21_X1 U339 ( .B1(n36), .B2(n457), .A(n502), .ZN(n461) );
  MUX2_X1 U340 ( .A(n458), .B(n461), .S(hwlp_counter_o[48]), .Z(n459) );
  NAND2_X1 U341 ( .A1(n460), .A2(n459), .ZN(n193) );
  NAND2_X1 U342 ( .A1(hwlp_cnt_data_i[17]), .A2(n446), .ZN(n464) );
  NAND2_X1 U343 ( .A1(n528), .A2(n465), .ZN(n467) );
  OAI21_X1 U344 ( .B1(n446), .B2(n564), .A(n461), .ZN(n462) );
  NAND2_X1 U345 ( .A1(n462), .A2(hwlp_counter_o[49]), .ZN(n463) );
  NAND3_X1 U346 ( .A1(n464), .A2(n467), .A3(n463), .ZN(n192) );
  NAND2_X1 U347 ( .A1(hwlp_cnt_data_i[18]), .A2(n508), .ZN(n469) );
  INV_X1 U348 ( .A(n465), .ZN(n466) );
  AOI21_X1 U349 ( .B1(n36), .B2(n466), .A(n502), .ZN(n470) );
  MUX2_X1 U350 ( .A(n467), .B(n470), .S(hwlp_counter_o[50]), .Z(n468) );
  NAND2_X1 U351 ( .A1(n469), .A2(n468), .ZN(n191) );
  NAND2_X1 U352 ( .A1(hwlp_cnt_data_i[19]), .A2(n446), .ZN(n473) );
  NAND2_X1 U353 ( .A1(n528), .A2(n474), .ZN(n476) );
  OAI21_X1 U354 ( .B1(n508), .B2(n559), .A(n470), .ZN(n471) );
  NAND2_X1 U355 ( .A1(n471), .A2(hwlp_counter_o[51]), .ZN(n472) );
  NAND3_X1 U356 ( .A1(n473), .A2(n476), .A3(n472), .ZN(n190) );
  NAND2_X1 U357 ( .A1(hwlp_cnt_data_i[20]), .A2(n508), .ZN(n478) );
  INV_X1 U358 ( .A(n474), .ZN(n475) );
  AOI21_X1 U359 ( .B1(n36), .B2(n475), .A(n502), .ZN(n479) );
  MUX2_X1 U360 ( .A(n476), .B(n479), .S(hwlp_counter_o[52]), .Z(n477) );
  NAND2_X1 U361 ( .A1(n478), .A2(n477), .ZN(n189) );
  NAND2_X1 U362 ( .A1(hwlp_cnt_data_i[21]), .A2(n446), .ZN(n482) );
  NAND2_X1 U363 ( .A1(n528), .A2(n483), .ZN(n485) );
  OAI21_X1 U364 ( .B1(n508), .B2(n565), .A(n479), .ZN(n480) );
  NAND2_X1 U365 ( .A1(n480), .A2(hwlp_counter_o[53]), .ZN(n481) );
  NAND3_X1 U366 ( .A1(n482), .A2(n485), .A3(n481), .ZN(n188) );
  NAND2_X1 U367 ( .A1(hwlp_cnt_data_i[22]), .A2(n508), .ZN(n487) );
  INV_X1 U368 ( .A(n483), .ZN(n484) );
  AOI21_X1 U369 ( .B1(n36), .B2(n484), .A(n502), .ZN(n488) );
  MUX2_X1 U370 ( .A(n485), .B(n488), .S(hwlp_counter_o[54]), .Z(n486) );
  NAND2_X1 U371 ( .A1(n487), .A2(n486), .ZN(n187) );
  NAND2_X1 U372 ( .A1(hwlp_cnt_data_i[23]), .A2(n446), .ZN(n491) );
  NAND2_X1 U373 ( .A1(n528), .A2(n492), .ZN(n494) );
  OAI21_X1 U374 ( .B1(n508), .B2(n569), .A(n488), .ZN(n489) );
  NAND2_X1 U375 ( .A1(n489), .A2(hwlp_counter_o[55]), .ZN(n490) );
  NAND3_X1 U376 ( .A1(n491), .A2(n494), .A3(n490), .ZN(n186) );
  NAND2_X1 U377 ( .A1(hwlp_cnt_data_i[24]), .A2(n508), .ZN(n496) );
  INV_X1 U378 ( .A(n492), .ZN(n493) );
  AOI21_X1 U379 ( .B1(n36), .B2(n493), .A(n502), .ZN(n497) );
  MUX2_X1 U380 ( .A(n494), .B(n497), .S(hwlp_counter_o[56]), .Z(n495) );
  NAND2_X1 U381 ( .A1(n496), .A2(n495), .ZN(n185) );
  NAND2_X1 U382 ( .A1(hwlp_cnt_data_i[25]), .A2(n446), .ZN(n500) );
  NAND2_X1 U383 ( .A1(n528), .A2(n501), .ZN(n504) );
  OAI21_X1 U384 ( .B1(n508), .B2(n556), .A(n497), .ZN(n498) );
  NAND2_X1 U385 ( .A1(n498), .A2(hwlp_counter_o[57]), .ZN(n499) );
  NAND3_X1 U386 ( .A1(n500), .A2(n504), .A3(n499), .ZN(n184) );
  NAND2_X1 U387 ( .A1(hwlp_cnt_data_i[26]), .A2(n508), .ZN(n506) );
  INV_X1 U388 ( .A(n501), .ZN(n503) );
  AOI21_X1 U389 ( .B1(n36), .B2(n503), .A(n502), .ZN(n507) );
  MUX2_X1 U390 ( .A(n504), .B(n507), .S(hwlp_counter_o[58]), .Z(n505) );
  NAND2_X1 U391 ( .A1(n506), .A2(n505), .ZN(n183) );
  NAND2_X1 U392 ( .A1(hwlp_cnt_data_i[27]), .A2(n508), .ZN(n512) );
  OAI21_X1 U393 ( .B1(n508), .B2(n553), .A(n507), .ZN(n510) );
  AOI22_X1 U394 ( .A1(n510), .A2(hwlp_counter_o[59]), .B1(n528), .B2(n509), 
        .ZN(n511) );
  NAND2_X1 U395 ( .A1(n512), .A2(n511), .ZN(n182) );
  NAND2_X1 U396 ( .A1(hwlp_cnt_data_i[29]), .A2(n508), .ZN(n518) );
  OAI21_X1 U397 ( .B1(n514), .B2(n549), .A(n513), .ZN(n516) );
  NOR2_X1 U398 ( .A1(n515), .A2(hwlp_counter_o[61]), .ZN(n522) );
  AOI21_X1 U399 ( .B1(hwlp_counter_o[61]), .B2(n516), .A(n522), .ZN(n517) );
  NAND2_X1 U400 ( .A1(n518), .A2(n517), .ZN(n180) );
  NAND2_X1 U401 ( .A1(hwlp_cnt_data_i[30]), .A2(n508), .ZN(n525) );
  OAI21_X1 U402 ( .B1(hwlp_counter_o[61]), .B2(n519), .A(n528), .ZN(n521) );
  NAND2_X1 U403 ( .A1(n521), .A2(n520), .ZN(n527) );
  INV_X1 U404 ( .A(n522), .ZN(n523) );
  NOR2_X1 U405 ( .A1(n523), .A2(hwlp_counter_o[62]), .ZN(n526) );
  AOI21_X1 U406 ( .B1(hwlp_counter_o[62]), .B2(n527), .A(n526), .ZN(n524) );
  NAND2_X1 U407 ( .A1(n525), .A2(n524), .ZN(n179) );
  NAND2_X1 U408 ( .A1(hwlp_cnt_data_i[31]), .A2(n508), .ZN(n532) );
  INV_X1 U409 ( .A(n526), .ZN(n530) );
  AOI21_X1 U410 ( .B1(n528), .B2(hwlp_counter_o[62]), .A(n527), .ZN(n529) );
  MUX2_X1 U411 ( .A(n530), .B(n529), .S(hwlp_counter_o[63]), .Z(n531) );
  NAND2_X1 U412 ( .A1(n532), .A2(n531), .ZN(n178) );
  INV_X1 U413 ( .A(hwlp_we_i[1]), .ZN(n533) );
  INV_X1 U462 ( .A(hwlp_regid_i[0]), .ZN(n537) );
  SDFFR_X1 hwlp_start_q_reg_1__31_ ( .D(hwlp_start_data_i[31]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[63]) );
  SDFFR_X1 hwlp_start_q_reg_1__30_ ( .D(hwlp_start_data_i[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[62]) );
  SDFFR_X1 hwlp_start_q_reg_1__29_ ( .D(hwlp_start_data_i[29]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[61]) );
  SDFFR_X1 hwlp_start_q_reg_1__28_ ( .D(hwlp_start_data_i[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[60]) );
  SDFFR_X1 hwlp_start_q_reg_1__27_ ( .D(hwlp_start_data_i[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[59]) );
  SDFFR_X1 hwlp_start_q_reg_1__26_ ( .D(hwlp_start_data_i[26]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[58]) );
  SDFFR_X1 hwlp_start_q_reg_1__25_ ( .D(hwlp_start_data_i[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[57]) );
  SDFFR_X1 hwlp_start_q_reg_1__24_ ( .D(hwlp_start_data_i[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[56]) );
  SDFFR_X1 hwlp_start_q_reg_1__23_ ( .D(hwlp_start_data_i[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[55]) );
  SDFFR_X1 hwlp_start_q_reg_1__22_ ( .D(hwlp_start_data_i[22]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[54]) );
  SDFFR_X1 hwlp_start_q_reg_1__21_ ( .D(hwlp_start_data_i[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[53]) );
  SDFFR_X1 hwlp_start_q_reg_1__20_ ( .D(hwlp_start_data_i[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[52]) );
  SDFFR_X1 hwlp_start_q_reg_1__19_ ( .D(hwlp_start_data_i[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[51]) );
  SDFFR_X1 hwlp_start_q_reg_1__18_ ( .D(hwlp_start_data_i[18]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[50]) );
  SDFFR_X1 hwlp_start_q_reg_1__17_ ( .D(hwlp_start_data_i[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[49]) );
  SDFFR_X1 hwlp_start_q_reg_1__16_ ( .D(hwlp_start_data_i[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[48]) );
  SDFFR_X1 hwlp_start_q_reg_1__15_ ( .D(hwlp_start_data_i[15]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[47]) );
  SDFFR_X1 hwlp_start_q_reg_1__14_ ( .D(hwlp_start_data_i[14]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[46]) );
  SDFFR_X1 hwlp_start_q_reg_1__13_ ( .D(hwlp_start_data_i[13]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[45]) );
  SDFFR_X1 hwlp_start_q_reg_1__12_ ( .D(hwlp_start_data_i[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[44]) );
  SDFFR_X1 hwlp_start_q_reg_1__10_ ( .D(hwlp_start_data_i[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[42]) );
  SDFFR_X1 hwlp_start_q_reg_1__9_ ( .D(hwlp_start_data_i[9]), .SI(1'b0), .SE(
        1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[41]) );
  SDFFR_X1 hwlp_start_q_reg_1__8_ ( .D(hwlp_start_data_i[8]), .SI(1'b0), .SE(
        1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[40]) );
  SDFFR_X1 hwlp_start_q_reg_1__7_ ( .D(hwlp_start_data_i[7]), .SI(1'b0), .SE(
        1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[39]) );
  SDFFR_X1 hwlp_start_q_reg_1__6_ ( .D(hwlp_start_data_i[6]), .SI(1'b0), .SE(
        1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[38]) );
  SDFFR_X1 hwlp_start_q_reg_1__5_ ( .D(hwlp_start_data_i[5]), .SI(1'b0), .SE(
        1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[37]) );
  SDFFR_X1 hwlp_start_q_reg_1__4_ ( .D(hwlp_start_data_i[4]), .SI(1'b0), .SE(
        1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[36]) );
  SDFFR_X1 hwlp_start_q_reg_1__3_ ( .D(hwlp_start_data_i[3]), .SI(1'b0), .SE(
        1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[35]) );
  SDFFR_X1 hwlp_start_q_reg_1__2_ ( .D(hwlp_start_data_i[2]), .SI(1'b0), .SE(
        1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[34]) );
  SDFFR_X1 hwlp_start_q_reg_1__1_ ( .D(hwlp_start_data_i[1]), .SI(1'b0), .SE(
        1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[33]) );
  SDFFR_X1 hwlp_start_q_reg_1__0_ ( .D(hwlp_start_data_i[0]), .SI(1'b0), .SE(
        1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[32]) );
  SDFFR_X1 hwlp_start_q_reg_0__31_ ( .D(hwlp_start_data_i[31]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[31]) );
  SDFFR_X1 hwlp_start_q_reg_0__30_ ( .D(hwlp_start_data_i[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[30]) );
  SDFFR_X1 hwlp_start_q_reg_0__29_ ( .D(hwlp_start_data_i[29]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[29]) );
  SDFFR_X1 hwlp_start_q_reg_0__28_ ( .D(hwlp_start_data_i[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[28]) );
  SDFFR_X1 hwlp_start_q_reg_0__27_ ( .D(hwlp_start_data_i[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[27]) );
  SDFFR_X1 hwlp_start_q_reg_0__26_ ( .D(hwlp_start_data_i[26]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[26]) );
  SDFFR_X1 hwlp_start_q_reg_0__25_ ( .D(hwlp_start_data_i[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[25]) );
  SDFFR_X1 hwlp_start_q_reg_0__24_ ( .D(hwlp_start_data_i[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[24]) );
  SDFFR_X1 hwlp_start_q_reg_0__23_ ( .D(hwlp_start_data_i[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[23]) );
  SDFFR_X1 hwlp_start_q_reg_0__22_ ( .D(hwlp_start_data_i[22]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[22]) );
  SDFFR_X1 hwlp_start_q_reg_0__21_ ( .D(hwlp_start_data_i[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[21]) );
  SDFFR_X1 hwlp_start_q_reg_0__20_ ( .D(hwlp_start_data_i[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[20]) );
  SDFFR_X1 hwlp_start_q_reg_0__19_ ( .D(hwlp_start_data_i[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[19]) );
  SDFFR_X1 hwlp_start_q_reg_0__18_ ( .D(hwlp_start_data_i[18]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[18]) );
  SDFFR_X1 hwlp_start_q_reg_0__17_ ( .D(hwlp_start_data_i[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[17]) );
  SDFFR_X1 hwlp_start_q_reg_0__16_ ( .D(hwlp_start_data_i[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[16]) );
  SDFFR_X1 hwlp_start_q_reg_0__15_ ( .D(hwlp_start_data_i[15]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[15]) );
  SDFFR_X1 hwlp_start_q_reg_0__14_ ( .D(hwlp_start_data_i[14]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[14]) );
  SDFFR_X1 hwlp_start_q_reg_0__13_ ( .D(hwlp_start_data_i[13]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[13]) );
  SDFFR_X1 hwlp_start_q_reg_0__12_ ( .D(hwlp_start_data_i[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[12]) );
  SDFFR_X1 hwlp_start_q_reg_0__11_ ( .D(hwlp_start_data_i[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[11]) );
  SDFFR_X1 hwlp_start_q_reg_0__10_ ( .D(hwlp_start_data_i[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[10]) );
  SDFFR_X1 hwlp_start_q_reg_0__9_ ( .D(hwlp_start_data_i[9]), .SI(1'b0), .SE(
        1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[9]) );
  SDFFR_X1 hwlp_start_q_reg_0__8_ ( .D(hwlp_start_data_i[8]), .SI(1'b0), .SE(
        1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[8]) );
  SDFFR_X1 hwlp_start_q_reg_0__7_ ( .D(hwlp_start_data_i[7]), .SI(1'b0), .SE(
        1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[7]) );
  SDFFR_X1 hwlp_start_q_reg_0__6_ ( .D(hwlp_start_data_i[6]), .SI(1'b0), .SE(
        1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[6]) );
  SDFFR_X1 hwlp_start_q_reg_0__5_ ( .D(hwlp_start_data_i[5]), .SI(1'b0), .SE(
        1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[5]) );
  SDFFR_X1 hwlp_start_q_reg_0__4_ ( .D(hwlp_start_data_i[4]), .SI(1'b0), .SE(
        1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[4]) );
  SDFFR_X1 hwlp_start_q_reg_0__3_ ( .D(hwlp_start_data_i[3]), .SI(1'b0), .SE(
        1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[3]) );
  SDFFR_X1 hwlp_start_q_reg_0__1_ ( .D(hwlp_start_data_i[1]), .SI(1'b0), .SE(
        1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[1]) );
  SDFFR_X1 hwlp_start_q_reg_0__0_ ( .D(hwlp_start_data_i[0]), .SI(1'b0), .SE(
        1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[0]) );
  SDFFR_X1 hwlp_end_q_reg_1__31_ ( .D(hwlp_end_data_i[31]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[63]) );
  SDFFR_X1 hwlp_end_q_reg_1__30_ ( .D(hwlp_end_data_i[30]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[62]) );
  SDFFR_X1 hwlp_end_q_reg_1__29_ ( .D(hwlp_end_data_i[29]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[61]) );
  SDFFR_X1 hwlp_end_q_reg_1__28_ ( .D(hwlp_end_data_i[28]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[60]) );
  SDFFR_X1 hwlp_end_q_reg_1__27_ ( .D(hwlp_end_data_i[27]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[59]) );
  SDFFR_X1 hwlp_end_q_reg_1__26_ ( .D(hwlp_end_data_i[26]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[58]) );
  SDFFR_X1 hwlp_end_q_reg_1__25_ ( .D(hwlp_end_data_i[25]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[57]) );
  SDFFR_X1 hwlp_end_q_reg_1__24_ ( .D(hwlp_end_data_i[24]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[56]) );
  SDFFR_X1 hwlp_end_q_reg_1__23_ ( .D(hwlp_end_data_i[23]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[55]) );
  SDFFR_X1 hwlp_end_q_reg_1__22_ ( .D(hwlp_end_data_i[22]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[54]) );
  SDFFR_X1 hwlp_end_q_reg_1__21_ ( .D(hwlp_end_data_i[21]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[53]) );
  SDFFR_X1 hwlp_end_q_reg_1__20_ ( .D(hwlp_end_data_i[20]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[52]) );
  SDFFR_X1 hwlp_end_q_reg_1__19_ ( .D(hwlp_end_data_i[19]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[51]) );
  SDFFR_X1 hwlp_end_q_reg_1__18_ ( .D(hwlp_end_data_i[18]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[50]) );
  SDFFR_X1 hwlp_end_q_reg_1__17_ ( .D(hwlp_end_data_i[17]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[49]) );
  SDFFR_X1 hwlp_end_q_reg_1__16_ ( .D(hwlp_end_data_i[16]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[48]) );
  SDFFR_X1 hwlp_end_q_reg_1__15_ ( .D(hwlp_end_data_i[15]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[47]) );
  SDFFR_X1 hwlp_end_q_reg_1__14_ ( .D(hwlp_end_data_i[14]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[46]) );
  SDFFR_X1 hwlp_end_q_reg_1__13_ ( .D(hwlp_end_data_i[13]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[45]) );
  SDFFR_X1 hwlp_end_q_reg_1__12_ ( .D(hwlp_end_data_i[12]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[44]) );
  SDFFR_X1 hwlp_end_q_reg_1__11_ ( .D(hwlp_end_data_i[11]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[43]) );
  SDFFR_X1 hwlp_end_q_reg_1__10_ ( .D(hwlp_end_data_i[10]), .SI(1'b0), .SE(
        1'b0), .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[42]) );
  SDFFR_X1 hwlp_end_q_reg_1__9_ ( .D(hwlp_end_data_i[9]), .SI(1'b0), .SE(1'b0), 
        .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[41]) );
  SDFFR_X1 hwlp_end_q_reg_1__8_ ( .D(hwlp_end_data_i[8]), .SI(1'b0), .SE(1'b0), 
        .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[40]) );
  SDFFR_X1 hwlp_end_q_reg_1__7_ ( .D(hwlp_end_data_i[7]), .SI(1'b0), .SE(1'b0), 
        .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[39]) );
  SDFFR_X1 hwlp_end_q_reg_1__6_ ( .D(hwlp_end_data_i[6]), .SI(1'b0), .SE(1'b0), 
        .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[38]) );
  SDFFR_X1 hwlp_end_q_reg_1__5_ ( .D(hwlp_end_data_i[5]), .SI(1'b0), .SE(1'b0), 
        .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[37]) );
  SDFFR_X1 hwlp_end_q_reg_1__4_ ( .D(hwlp_end_data_i[4]), .SI(1'b0), .SE(1'b0), 
        .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[36]) );
  SDFFR_X1 hwlp_end_q_reg_1__3_ ( .D(hwlp_end_data_i[3]), .SI(1'b0), .SE(1'b0), 
        .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[35]) );
  SDFFR_X1 hwlp_end_q_reg_1__2_ ( .D(hwlp_end_data_i[2]), .SI(1'b0), .SE(1'b0), 
        .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[34]) );
  SDFFR_X1 hwlp_end_q_reg_1__1_ ( .D(hwlp_end_data_i[1]), .SI(1'b0), .SE(1'b0), 
        .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[33]) );
  SDFFR_X1 hwlp_end_q_reg_1__0_ ( .D(hwlp_end_data_i[0]), .SI(1'b0), .SE(1'b0), 
        .CK(n967), .RN(rst_n), .Q(hwlp_end_addr_o[32]) );
  SDFFR_X1 hwlp_end_q_reg_0__31_ ( .D(hwlp_end_data_i[31]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[31]) );
  SDFFR_X1 hwlp_end_q_reg_0__30_ ( .D(hwlp_end_data_i[30]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[30]) );
  SDFFR_X1 hwlp_end_q_reg_0__29_ ( .D(hwlp_end_data_i[29]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[29]) );
  SDFFR_X1 hwlp_end_q_reg_0__28_ ( .D(hwlp_end_data_i[28]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[28]) );
  SDFFR_X1 hwlp_end_q_reg_0__27_ ( .D(hwlp_end_data_i[27]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[27]) );
  SDFFR_X1 hwlp_end_q_reg_0__26_ ( .D(hwlp_end_data_i[26]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[26]) );
  SDFFR_X1 hwlp_end_q_reg_0__25_ ( .D(hwlp_end_data_i[25]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[25]) );
  SDFFR_X1 hwlp_end_q_reg_0__24_ ( .D(hwlp_end_data_i[24]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[24]) );
  SDFFR_X1 hwlp_end_q_reg_0__23_ ( .D(hwlp_end_data_i[23]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[23]) );
  SDFFR_X1 hwlp_end_q_reg_0__22_ ( .D(hwlp_end_data_i[22]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[22]) );
  SDFFR_X1 hwlp_end_q_reg_0__21_ ( .D(hwlp_end_data_i[21]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[21]) );
  SDFFR_X1 hwlp_end_q_reg_0__20_ ( .D(hwlp_end_data_i[20]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[20]) );
  SDFFR_X1 hwlp_end_q_reg_0__19_ ( .D(hwlp_end_data_i[19]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[19]) );
  SDFFR_X1 hwlp_end_q_reg_0__18_ ( .D(hwlp_end_data_i[18]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[18]) );
  SDFFR_X1 hwlp_end_q_reg_0__17_ ( .D(hwlp_end_data_i[17]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[17]) );
  SDFFR_X1 hwlp_end_q_reg_0__16_ ( .D(hwlp_end_data_i[16]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[16]) );
  SDFFR_X1 hwlp_end_q_reg_0__15_ ( .D(hwlp_end_data_i[15]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[15]) );
  SDFFR_X1 hwlp_end_q_reg_0__14_ ( .D(hwlp_end_data_i[14]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[14]) );
  SDFFR_X1 hwlp_end_q_reg_0__13_ ( .D(hwlp_end_data_i[13]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[13]) );
  SDFFR_X1 hwlp_end_q_reg_0__12_ ( .D(hwlp_end_data_i[12]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[12]) );
  SDFFR_X1 hwlp_end_q_reg_0__11_ ( .D(hwlp_end_data_i[11]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[11]) );
  SDFFR_X1 hwlp_end_q_reg_0__10_ ( .D(hwlp_end_data_i[10]), .SI(1'b0), .SE(
        1'b0), .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[10]) );
  SDFFR_X1 hwlp_end_q_reg_0__9_ ( .D(hwlp_end_data_i[9]), .SI(1'b0), .SE(1'b0), 
        .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[9]) );
  SDFFR_X1 hwlp_end_q_reg_0__8_ ( .D(hwlp_end_data_i[8]), .SI(1'b0), .SE(1'b0), 
        .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[8]) );
  SDFFR_X1 hwlp_end_q_reg_0__7_ ( .D(hwlp_end_data_i[7]), .SI(1'b0), .SE(1'b0), 
        .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[7]) );
  SDFFR_X1 hwlp_end_q_reg_0__6_ ( .D(hwlp_end_data_i[6]), .SI(1'b0), .SE(1'b0), 
        .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[6]) );
  SDFFR_X1 hwlp_end_q_reg_0__5_ ( .D(hwlp_end_data_i[5]), .SI(1'b0), .SE(1'b0), 
        .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[5]) );
  SDFFR_X1 hwlp_end_q_reg_0__4_ ( .D(hwlp_end_data_i[4]), .SI(1'b0), .SE(1'b0), 
        .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[4]) );
  SDFFR_X1 hwlp_end_q_reg_0__3_ ( .D(hwlp_end_data_i[3]), .SI(1'b0), .SE(1'b0), 
        .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[3]) );
  SDFFR_X1 hwlp_end_q_reg_0__2_ ( .D(hwlp_end_data_i[2]), .SI(1'b0), .SE(1'b0), 
        .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[2]) );
  SDFFR_X1 hwlp_end_q_reg_0__1_ ( .D(hwlp_end_data_i[1]), .SI(1'b0), .SE(1'b0), 
        .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[1]) );
  SDFFR_X1 hwlp_end_q_reg_0__0_ ( .D(hwlp_end_data_i[0]), .SI(1'b0), .SE(1'b0), 
        .CK(n965), .RN(rst_n), .Q(hwlp_end_addr_o[0]) );
  SDFFR_X1 hwlp_counter_q_reg_1__31_ ( .D(n178), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[63]) );
  SDFFR_X1 hwlp_counter_q_reg_1__30_ ( .D(n179), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[62]) );
  SDFFR_X1 hwlp_counter_q_reg_1__29_ ( .D(n180), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[61]) );
  SDFFR_X1 hwlp_counter_q_reg_1__27_ ( .D(n182), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[59]) );
  SDFFR_X1 hwlp_counter_q_reg_1__24_ ( .D(n185), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[56]), .QN(n556) );
  SDFFR_X1 hwlp_counter_q_reg_1__23_ ( .D(n186), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[55]) );
  SDFFR_X1 hwlp_counter_q_reg_1__22_ ( .D(n187), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[54]), .QN(n569) );
  SDFFR_X1 hwlp_counter_q_reg_1__21_ ( .D(n188), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[53]) );
  SDFFR_X1 hwlp_counter_q_reg_1__20_ ( .D(n189), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[52]), .QN(n565) );
  SDFFR_X1 hwlp_counter_q_reg_1__19_ ( .D(n190), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[51]) );
  SDFFR_X1 hwlp_counter_q_reg_1__18_ ( .D(n191), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[50]), .QN(n559) );
  SDFFR_X1 hwlp_counter_q_reg_1__17_ ( .D(n192), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[49]) );
  SDFFR_X1 hwlp_counter_q_reg_1__16_ ( .D(n193), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[48]), .QN(n564) );
  SDFFR_X1 hwlp_counter_q_reg_1__15_ ( .D(n194), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[47]) );
  SDFFR_X1 hwlp_counter_q_reg_1__14_ ( .D(n195), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[46]), .QN(n568) );
  SDFFR_X1 hwlp_counter_q_reg_1__13_ ( .D(n196), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[45]) );
  SDFFR_X1 hwlp_counter_q_reg_1__11_ ( .D(n198), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[43]) );
  SDFFR_X1 hwlp_counter_q_reg_1__10_ ( .D(n199), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[42]), .QN(n555) );
  SDFFR_X1 hwlp_counter_q_reg_1__9_ ( .D(n200), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[41]), .QN(n574) );
  SDFFR_X1 hwlp_counter_q_reg_1__8_ ( .D(n201), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[40]) );
  SDFFR_X1 hwlp_counter_q_reg_1__7_ ( .D(n202), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[39]) );
  SDFFR_X1 hwlp_counter_q_reg_1__6_ ( .D(n203), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[38]), .QN(n545) );
  SDFFR_X1 hwlp_counter_q_reg_1__5_ ( .D(n204), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[37]) );
  SDFFR_X1 hwlp_counter_q_reg_1__3_ ( .D(n206), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[35]), .QN(n571) );
  SDFFR_X1 hwlp_counter_q_reg_1__2_ ( .D(n207), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[34]), .QN(n543) );
  SDFFR_X1 hwlp_counter_q_reg_1__1_ ( .D(n208), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[33]), .QN(n561) );
  SDFFR_X1 hwlp_counter_q_reg_1__0_ ( .D(n209), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[32]), .QN(n552) );
  SDFFR_X1 hwlp_counter_q_reg_0__31_ ( .D(n146), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[31]) );
  SDFFR_X1 hwlp_counter_q_reg_0__30_ ( .D(n147), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[30]) );
  SDFFR_X1 hwlp_counter_q_reg_0__29_ ( .D(n148), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[29]) );
  SDFFR_X1 hwlp_counter_q_reg_0__27_ ( .D(n150), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[27]) );
  SDFFR_X1 hwlp_counter_q_reg_0__26_ ( .D(n151), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[26]), .QN(n558) );
  SDFFR_X1 hwlp_counter_q_reg_0__24_ ( .D(n153), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[24]), .QN(n560) );
  SDFFR_X1 hwlp_counter_q_reg_0__23_ ( .D(n154), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[23]) );
  SDFFR_X1 hwlp_counter_q_reg_0__22_ ( .D(n155), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[22]), .QN(n567) );
  SDFFR_X1 hwlp_counter_q_reg_0__21_ ( .D(n156), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[21]) );
  SDFFR_X1 hwlp_counter_q_reg_0__20_ ( .D(n157), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[20]), .QN(n562) );
  SDFFR_X1 hwlp_counter_q_reg_0__19_ ( .D(n158), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[19]) );
  SDFFR_X1 hwlp_counter_q_reg_0__18_ ( .D(n159), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[18]), .QN(n557) );
  SDFFR_X1 hwlp_counter_q_reg_0__17_ ( .D(n160), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[17]) );
  SDFFR_X1 hwlp_counter_q_reg_0__16_ ( .D(n161), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[16]), .QN(n563) );
  SDFFR_X1 hwlp_counter_q_reg_0__15_ ( .D(n162), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[15]) );
  SDFFR_X1 hwlp_counter_q_reg_0__14_ ( .D(n163), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[14]), .QN(n566) );
  SDFFR_X1 hwlp_counter_q_reg_0__13_ ( .D(n164), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[13]) );
  SDFFR_X1 hwlp_counter_q_reg_0__12_ ( .D(n165), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[12]), .QN(n546) );
  SDFFR_X1 hwlp_counter_q_reg_0__11_ ( .D(n166), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[11]) );
  SDFFR_X1 hwlp_counter_q_reg_0__10_ ( .D(n167), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[10]), .QN(n554) );
  SDFFR_X1 hwlp_counter_q_reg_0__9_ ( .D(n168), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[9]), .QN(n573) );
  SDFFR_X1 hwlp_counter_q_reg_0__8_ ( .D(n169), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[8]) );
  SDFFR_X1 hwlp_counter_q_reg_0__7_ ( .D(n170), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[7]) );
  SDFFR_X1 hwlp_counter_q_reg_0__6_ ( .D(n171), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[6]), .QN(n544) );
  SDFFR_X1 hwlp_counter_q_reg_0__5_ ( .D(n172), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[5]) );
  SDFFR_X1 hwlp_counter_q_reg_0__4_ ( .D(n173), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[4]), .QN(n550) );
  SDFFR_X1 hwlp_counter_q_reg_0__3_ ( .D(n174), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[3]), .QN(n570) );
  SDFFR_X1 hwlp_counter_q_reg_0__2_ ( .D(n175), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[2]), .QN(n542) );
  SDFFR_X1 hwlp_counter_q_reg_0__1_ ( .D(n176), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[1]), .QN(n572) );
  SDFFR_X1 hwlp_counter_q_reg_0__0_ ( .D(n177), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[0]) );
  SNPS_CLOCK_GATE_HIGH_riscv_hwloop_regs_N_REGS2_0 clk_gate_hwlp_start_q_reg_1__0_ ( 
        .CLK(clk), .EN(n589), .ENCLK(n971), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_hwloop_regs_N_REGS2_1 clk_gate_hwlp_start_q_reg_0__2_ ( 
        .CLK(clk), .EN(n588), .ENCLK(n969), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_hwloop_regs_N_REGS2_2 clk_gate_hwlp_end_q_reg_1__0_ ( 
        .CLK(clk), .EN(n587), .ENCLK(n967), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_hwloop_regs_N_REGS2_3 clk_gate_hwlp_end_q_reg_0__0_ ( 
        .CLK(clk), .EN(n586), .ENCLK(n965), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_hwloop_regs_N_REGS2_4 clk_gate_hwlp_counter_q_reg_1__9_ ( 
        .CLK(clk), .EN(n964), .ENCLK(n962), .TE(1'b0) );
  SDFFR_X2 hwlp_counter_q_reg_1__25_ ( .D(n184), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[57]) );
  SDFFR_X2 hwlp_counter_q_reg_0__25_ ( .D(n152), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[25]) );
  SDFFR_X1 hwlp_counter_q_reg_0__28_ ( .D(n149), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[28]), .QN(n548) );
  SDFFR_X1 hwlp_counter_q_reg_1__26_ ( .D(n183), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[58]), .QN(n553) );
  SDFFR_X2 hwlp_start_q_reg_0__2_ ( .D(hwlp_start_data_i[2]), .SI(1'b0), .SE(
        1'b0), .CK(n969), .RN(rst_n), .Q(hwlp_start_addr_o[2]) );
  SDFFR_X2 hwlp_counter_q_reg_1__4_ ( .D(n205), .SI(1'b0), .SE(1'b0), .CK(n962), .RN(rst_n), .Q(hwlp_counter_o[36]), .QN(n551) );
  SDFFR_X2 hwlp_counter_q_reg_1__12_ ( .D(n197), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[44]), .QN(n547) );
  SDFFR_X1 hwlp_counter_q_reg_1__28_ ( .D(n181), .SI(1'b0), .SE(1'b0), .CK(
        n962), .RN(rst_n), .Q(hwlp_counter_o[60]), .QN(n549) );
  INV_X1 U12 ( .A(n36), .ZN(n508) );
  INV_X1 U13 ( .A(n17), .ZN(n360) );
  NAND2_X1 U14 ( .A1(n372), .A2(n17), .ZN(n366) );
  INV_X1 U105 ( .A(n514), .ZN(n528) );
  SDFFR_X1 hwlp_start_q_reg_1__11_ ( .D(hwlp_start_data_i[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n971), .RN(rst_n), .Q(hwlp_start_addr_o[43]) );
  OR2_X1 U3 ( .A1(hwlp_regid_i[0]), .A2(n1), .ZN(n17) );
  INV_X1 U4 ( .A(n366), .ZN(n381) );
  NAND2_X1 U5 ( .A1(hwlp_regid_i[0]), .A2(hwlp_we_i[2]), .ZN(n36) );
  BUF_X1 U6 ( .A(n378), .Z(n575) );
  INV_X1 U7 ( .A(n36), .ZN(n446) );
  INV_X1 U8 ( .A(n17), .ZN(n378) );
  NAND2_X1 U56 ( .A1(n583), .A2(n582), .ZN(n181) );
  INV_X1 U95 ( .A(n38), .ZN(n582) );
  NAND2_X1 U96 ( .A1(hwlp_cnt_data_i[28]), .A2(n508), .ZN(n583) );
  NAND2_X1 U414 ( .A1(n585), .A2(n584), .ZN(n149) );
  INV_X1 U415 ( .A(n19), .ZN(n584) );
  NAND2_X1 U416 ( .A1(hwlp_cnt_data_i[28]), .A2(n360), .ZN(n585) );
  NOR2_X1 U417 ( .A1(hwlp_regid_i[0]), .A2(n533), .ZN(n586) );
  AND2_X1 U418 ( .A1(hwlp_regid_i[0]), .A2(hwlp_we_i[1]), .ZN(n587) );
  AND2_X1 U419 ( .A1(hwlp_we_i[0]), .A2(n537), .ZN(n588) );
  AND2_X1 U420 ( .A1(hwlp_regid_i[0]), .A2(hwlp_we_i[0]), .ZN(n589) );
  OR2_X1 U794 ( .A1(valid_i), .A2(hwlp_we_i[2]), .ZN(n964) );
endmodule


module riscv_int_controller_PULP_SECURE1 ( clk, rst_n, irq_req_ctrl_o, 
        irq_sec_ctrl_o, irq_id_ctrl_o, ctrl_kill_i, irq_i, irq_sec_i, irq_id_i, 
        m_IE_i, u_IE_i, current_priv_lvl_i, ctrl_ack_i_BAR );
  output [4:0] irq_id_ctrl_o;
  input [4:0] irq_id_i;
  input [1:0] current_priv_lvl_i;
  input clk, rst_n, ctrl_kill_i, irq_i, irq_sec_i, m_IE_i, u_IE_i,
         ctrl_ack_i_BAR;
  output irq_req_ctrl_o, irq_sec_ctrl_o;
  wire   n20, n21, n22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n23, n40, n42;
  wire   [1:0] exc_ctrl_cs;

  INV_X1 U26 ( .A(rst_n) );
  INV_X1 U3 ( .A(ctrl_kill_i), .ZN(n7) );
  AOI21_X1 U4 ( .B1(n7), .B2(ctrl_ack_i_BAR), .A(exc_ctrl_cs[1]), .ZN(n5) );
  INV_X1 U5 ( .A(current_priv_lvl_i[1]), .ZN(n1) );
  OAI21_X1 U6 ( .B1(u_IE_i), .B2(irq_sec_i), .A(n1), .ZN(n3) );
  NAND3_X1 U7 ( .A1(current_priv_lvl_i[0]), .A2(current_priv_lvl_i[1]), .A3(
        m_IE_i), .ZN(n2) );
  OAI21_X1 U8 ( .B1(current_priv_lvl_i[0]), .B2(n3), .A(n2), .ZN(n4) );
  NAND2_X1 U9 ( .A1(irq_i), .A2(n4), .ZN(n9) );
  OR3_X1 U10 ( .A1(n9), .A2(exc_ctrl_cs[0]), .A3(exc_ctrl_cs[1]), .ZN(n11) );
  OAI21_X1 U11 ( .B1(n5), .B2(n13), .A(n11), .ZN(n22) );
  INV_X1 U12 ( .A(ctrl_ack_i_BAR), .ZN(n6) );
  AOI21_X1 U13 ( .B1(n7), .B2(n6), .A(exc_ctrl_cs[1]), .ZN(n8) );
  NOR2_X1 U14 ( .A1(n8), .A2(n13), .ZN(n21) );
  AOI21_X1 U20 ( .B1(n9), .B2(n14), .A(exc_ctrl_cs[0]), .ZN(n12) );
  INV_X1 U21 ( .A(irq_sec_i), .ZN(n10) );
  OAI22_X1 U22 ( .A1(n12), .A2(n23), .B1(n11), .B2(n10), .ZN(n20) );
  NOR2_X1 U23 ( .A1(n13), .A2(exc_ctrl_cs[1]), .ZN(irq_req_ctrl_o) );
  SDFFR_X1 exc_ctrl_cs_reg_0_ ( .D(n22), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(exc_ctrl_cs[0]), .QN(n13) );
  SDFFR_X1 exc_ctrl_cs_reg_1_ ( .D(n21), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(exc_ctrl_cs[1]), .QN(n14) );
  SDFFR_X1 irq_sec_q_reg ( .D(n20), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(rst_n), 
        .Q(irq_sec_ctrl_o), .QN(n23) );
  SDFFR_X1 irq_id_q_reg_4_ ( .D(irq_id_i[4]), .SI(1'b0), .SE(1'b0), .CK(n40), 
        .RN(rst_n), .Q(irq_id_ctrl_o[4]) );
  SDFFR_X1 irq_id_q_reg_3_ ( .D(irq_id_i[3]), .SI(1'b0), .SE(1'b0), .CK(n40), 
        .RN(rst_n), .Q(irq_id_ctrl_o[3]) );
  SDFFR_X1 irq_id_q_reg_2_ ( .D(irq_id_i[2]), .SI(1'b0), .SE(1'b0), .CK(n40), 
        .RN(rst_n), .Q(irq_id_ctrl_o[2]) );
  SDFFR_X1 irq_id_q_reg_1_ ( .D(irq_id_i[1]), .SI(1'b0), .SE(1'b0), .CK(n40), 
        .RN(rst_n), .Q(irq_id_ctrl_o[1]) );
  SDFFR_X1 irq_id_q_reg_0_ ( .D(irq_id_i[0]), .SI(1'b0), .SE(1'b0), .CK(n40), 
        .RN(rst_n), .Q(irq_id_ctrl_o[0]) );
  SNPS_CLOCK_GATE_HIGH_riscv_int_controller_PULP_SECURE1_0 clk_gate_irq_id_q_reg_0_ ( 
        .CLK(clk), .EN(n42), .ENCLK(n40), .TE(1'b0) );
  INV_X1 U37 ( .A(n11), .ZN(n42) );
endmodule


module riscv_controller_FPU0 ( clk, rst_n, fetch_enable_i, ctrl_busy_o, 
        first_fetch_o, is_fetch_failed_i, deassert_we_o, illegal_insn_i, 
        ecall_insn_i, mret_insn_i, uret_insn_i, dret_insn_i, mret_dec_i, 
        uret_dec_i, dret_dec_i, pipe_flush_i, ebrk_insn_i, fencei_insn_i, 
        csr_status_i, instr_multicycle_i, instr_valid_i, instr_req_o, pc_set_o, 
        pc_mux_o, exc_pc_mux_o, trap_addr_mux_o, data_req_ex_i, data_we_ex_i, 
        data_misaligned_i, data_load_event_i, mult_multicycle_i, apu_en_i, 
        apu_read_dep_i, apu_write_dep_i, apu_stall_o, branch_taken_ex_i, 
        jump_in_id_i, jump_in_dec_i, irq_i, irq_req_ctrl_i, irq_sec_ctrl_i, 
        irq_id_ctrl_i, m_IE_i, u_IE_i, current_priv_lvl_i, irq_id_o, 
        exc_cause_o, exc_kill_o, debug_mode_o, debug_cause_o, debug_csr_save_o, 
        debug_req_i, debug_single_step_i, debug_ebreakm_i, debug_ebreaku_i, 
        csr_save_if_o, csr_save_id_o, csr_irq_sec_o, csr_restore_mret_id_o, 
        csr_restore_uret_id_o, csr_restore_dret_id_o, csr_save_cause_o, 
        regfile_we_id_i, regfile_alu_waddr_id_i, regfile_we_ex_i, 
        regfile_waddr_ex_i, regfile_we_wb_i, regfile_alu_we_fw_i, 
        operand_a_fw_mux_sel_o, operand_b_fw_mux_sel_o, reg_d_ex_is_reg_a_i, 
        reg_d_ex_is_reg_b_i, reg_d_ex_is_reg_c_i, reg_d_wb_is_reg_a_i, 
        reg_d_wb_is_reg_b_i, reg_d_wb_is_reg_c_i, reg_d_alu_is_reg_a_i, 
        reg_d_alu_is_reg_b_i, reg_d_alu_is_reg_c_i, halt_if_o, 
        misaligned_stall_o, jr_stall_o, load_stall_o, ex_valid_i, wb_ready_i, 
        perf_jump_o, perf_jr_stall_o, perf_ld_stall_o, perf_pipeline_stall_o, 
        irq_ack_o_BAR, exc_ack_o_BAR, csr_cause_o_5__BAR, csr_cause_o_4_, 
        csr_cause_o_3_, csr_cause_o_2_, csr_cause_o_0_, id_ready_i_BAR, 
        data_err_ack_o_BAR, csr_save_ex_o_BAR, data_err_i_BAR, 
        csr_cause_o_1__BAR, halt_id_o_BAR, operand_c_fw_mux_sel_o_1_, 
        operand_c_fw_mux_sel_o_0__BAR, is_decoding_o );
  output [2:0] pc_mux_o;
  output [2:0] exc_pc_mux_o;
  input [1:0] jump_in_id_i;
  input [1:0] jump_in_dec_i;
  input [4:0] irq_id_ctrl_i;
  input [1:0] current_priv_lvl_i;
  output [4:0] irq_id_o;
  output [5:0] exc_cause_o;
  output [2:0] debug_cause_o;
  input [5:0] regfile_alu_waddr_id_i;
  input [5:0] regfile_waddr_ex_i;
  output [1:0] operand_a_fw_mux_sel_o;
  output [1:0] operand_b_fw_mux_sel_o;
  input clk, rst_n, fetch_enable_i, is_fetch_failed_i, illegal_insn_i,
         ecall_insn_i, mret_insn_i, uret_insn_i, dret_insn_i, mret_dec_i,
         uret_dec_i, dret_dec_i, pipe_flush_i, ebrk_insn_i, fencei_insn_i,
         csr_status_i, instr_multicycle_i, instr_valid_i, data_req_ex_i,
         data_we_ex_i, data_misaligned_i, data_load_event_i, mult_multicycle_i,
         apu_en_i, apu_read_dep_i, apu_write_dep_i, branch_taken_ex_i, irq_i,
         irq_req_ctrl_i, irq_sec_ctrl_i, m_IE_i, u_IE_i, debug_req_i,
         debug_single_step_i, debug_ebreakm_i, debug_ebreaku_i,
         regfile_we_id_i, regfile_we_ex_i, regfile_we_wb_i,
         regfile_alu_we_fw_i, reg_d_ex_is_reg_a_i, reg_d_ex_is_reg_b_i,
         reg_d_ex_is_reg_c_i, reg_d_wb_is_reg_a_i, reg_d_wb_is_reg_b_i,
         reg_d_wb_is_reg_c_i, reg_d_alu_is_reg_a_i, reg_d_alu_is_reg_b_i,
         reg_d_alu_is_reg_c_i, ex_valid_i, wb_ready_i, id_ready_i_BAR,
         data_err_i_BAR;
  output ctrl_busy_o, first_fetch_o, deassert_we_o, instr_req_o, pc_set_o,
         trap_addr_mux_o, apu_stall_o, exc_kill_o, debug_mode_o,
         debug_csr_save_o, csr_save_if_o, csr_save_id_o, csr_irq_sec_o,
         csr_restore_mret_id_o, csr_restore_uret_id_o, csr_restore_dret_id_o,
         csr_save_cause_o, halt_if_o, misaligned_stall_o, jr_stall_o,
         load_stall_o, perf_jump_o, perf_jr_stall_o, perf_ld_stall_o,
         perf_pipeline_stall_o, irq_ack_o_BAR, exc_ack_o_BAR,
         csr_cause_o_5__BAR, csr_cause_o_4_, csr_cause_o_3_, csr_cause_o_2_,
         csr_cause_o_0_, data_err_ack_o_BAR, csr_save_ex_o_BAR,
         csr_cause_o_1__BAR, halt_id_o_BAR, operand_c_fw_mux_sel_o_1_,
         operand_c_fw_mux_sel_o_0__BAR, is_decoding_o;
  wire   n101, \exc_cause_o[4] , data_misaligned_i, load_stall_o, jump_done_q,
         illegal_insn_q, instr_valid_irq_flush_n, instr_valid_irq_flush_q,
         data_err_q, jr_stall_o, N448, csr_save_ex_o_BAR, csr_cause_o_5__BAR,
         n263, n264, n265, n266, n267, n268, n269, n103, n104, n105, n106,
         n107, n108, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182,
         is_decoding_o_BAR, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n258, n259,
         n260, n261, n262, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n417, n421;
  wire   [4:0] ctrl_fsm_cs;
  assign irq_id_o[4] = irq_id_ctrl_i[4];
  assign irq_id_o[3] = irq_id_ctrl_i[3];
  assign irq_id_o[2] = irq_id_ctrl_i[2];
  assign irq_id_o[1] = irq_id_ctrl_i[1];
  assign irq_id_o[0] = irq_id_ctrl_i[0];
  assign csr_cause_o_4_ = \exc_cause_o[4] ;
  assign exc_cause_o[4] = \exc_cause_o[4] ;
  assign misaligned_stall_o = data_misaligned_i;
  assign perf_ld_stall_o = load_stall_o;
  assign perf_jr_stall_o = jr_stall_o;
  assign data_err_ack_o_BAR = csr_save_ex_o_BAR;
  assign irq_ack_o_BAR = csr_cause_o_5__BAR;
  assign exc_ack_o_BAR = csr_cause_o_5__BAR;

  INV_X1 U320 ( .A(rst_n) );
  NAND2_X1 U4 ( .A1(n138), .A2(n111), .ZN(pc_set_o) );
  OR3_X2 U5 ( .A1(debug_req_i), .A2(n147), .A3(n107), .ZN(n113) );
  CLKBUF_X1 U7 ( .A(ecall_insn_i), .Z(n105) );
  NOR2_X1 U8 ( .A1(n191), .A2(n190), .ZN(halt_id_o_BAR) );
  AND2_X1 U9 ( .A1(n270), .A2(n204), .ZN(is_decoding_o) );
  INV_X1 U12 ( .A(n148), .ZN(n114) );
  NAND2_X1 U13 ( .A1(n122), .A2(csr_cause_o_5__BAR), .ZN(pc_mux_o[2]) );
  OR2_X1 U14 ( .A1(n204), .A2(n145), .ZN(n117) );
  NOR2_X1 U15 ( .A1(n381), .A2(n228), .ZN(n204) );
  NOR2_X1 U17 ( .A1(ctrl_fsm_cs[3]), .A2(ctrl_fsm_cs[4]), .ZN(n377) );
  OR2_X1 U18 ( .A1(n412), .A2(ctrl_fsm_cs[4]), .ZN(n403) );
  NAND4_X4 U19 ( .A1(n106), .A2(n113), .A3(n114), .A4(n108), .ZN(pc_mux_o[1])
         );
  NAND2_X1 U20 ( .A1(n104), .A2(jump_in_dec_i[1]), .ZN(n179) );
  NAND3_X1 U21 ( .A1(n123), .A2(n360), .A3(n359), .ZN(n104) );
  NAND2_X2 U22 ( .A1(n116), .A2(n115), .ZN(pc_mux_o[0]) );
  NAND2_X1 U23 ( .A1(branch_taken_ex_i), .A2(n117), .ZN(n106) );
  OR2_X1 U24 ( .A1(n142), .A2(n143), .ZN(n107) );
  AND2_X1 U25 ( .A1(n151), .A2(n108), .ZN(n115) );
  AND2_X1 U27 ( .A1(n139), .A2(n127), .ZN(n110) );
  AOI22_X1 U28 ( .A1(n178), .A2(n177), .B1(n176), .B2(n175), .ZN(load_stall_o)
         );
  OR2_X1 U29 ( .A1(n145), .A2(n137), .ZN(n112) );
  OR2_X1 U32 ( .A1(n144), .A2(n199), .ZN(n108) );
  OR4_X1 U33 ( .A1(load_stall_o), .A2(illegal_insn_i), .A3(jr_stall_o), .A4(
        is_decoding_o_BAR), .ZN(deassert_we_o) );
  NAND2_X1 U35 ( .A1(n347), .A2(n112), .ZN(n111) );
  NAND2_X1 U36 ( .A1(branch_taken_ex_i), .A2(n117), .ZN(n116) );
  NAND2_X1 U37 ( .A1(n103), .A2(n204), .ZN(n212) );
  OR2_X1 U38 ( .A1(pc_mux_o[2]), .A2(n134), .ZN(n118) );
  NOR2_X1 U39 ( .A1(n179), .A2(jump_in_dec_i[0]), .ZN(jr_stall_o) );
  NOR2_X1 U40 ( .A1(n141), .A2(ctrl_fsm_cs[1]), .ZN(n282) );
  AND2_X1 U41 ( .A1(ctrl_fsm_cs[1]), .A2(ctrl_fsm_cs[2]), .ZN(n196) );
  NAND2_X1 U42 ( .A1(n377), .A2(n196), .ZN(csr_cause_o_5__BAR) );
  NOR2_X1 U43 ( .A1(current_priv_lvl_i[1]), .A2(current_priv_lvl_i[0]), .ZN(
        n157) );
  INV_X1 U44 ( .A(n157), .ZN(n365) );
  OR2_X1 U45 ( .A1(ecall_insn_i), .A2(ebrk_insn_i), .ZN(n237) );
  NOR2_X1 U46 ( .A1(data_err_q), .A2(illegal_insn_q), .ZN(n309) );
  INV_X1 U47 ( .A(n309), .ZN(n149) );
  AND2_X1 U48 ( .A1(n410), .A2(ctrl_fsm_cs[0]), .ZN(n311) );
  OAI21_X1 U49 ( .B1(n237), .B2(n149), .A(n311), .ZN(n119) );
  OR2_X1 U50 ( .A1(n410), .A2(ctrl_fsm_cs[0]), .ZN(n322) );
  AOI21_X1 U51 ( .B1(n119), .B2(n322), .A(n408), .ZN(n121) );
  AND2_X1 U52 ( .A1(n408), .A2(ctrl_fsm_cs[2]), .ZN(n310) );
  NOR2_X1 U53 ( .A1(mret_dec_i), .A2(uret_insn_i), .ZN(n193) );
  AND2_X1 U54 ( .A1(ctrl_fsm_cs[2]), .A2(ctrl_fsm_cs[0]), .ZN(n275) );
  OR2_X1 U55 ( .A1(n275), .A2(ctrl_fsm_cs[1]), .ZN(n165) );
  NOR2_X1 U56 ( .A1(dret_dec_i), .A2(n165), .ZN(n120) );
  AOI21_X1 U57 ( .B1(n193), .B2(n120), .A(n403), .ZN(n132) );
  OAI21_X1 U58 ( .B1(n121), .B2(n310), .A(n132), .ZN(n122) );
  NAND2_X1 U59 ( .A1(reg_d_alu_is_reg_a_i), .A2(regfile_alu_we_fw_i), .ZN(n359) );
  NAND2_X1 U60 ( .A1(reg_d_wb_is_reg_a_i), .A2(regfile_we_wb_i), .ZN(n360) );
  NAND2_X1 U61 ( .A1(reg_d_ex_is_reg_a_i), .A2(regfile_we_ex_i), .ZN(n123) );
  XNOR2_X1 U62 ( .A(jump_in_dec_i[1]), .B(jump_in_dec_i[0]), .ZN(n396) );
  INV_X1 U63 ( .A(n396), .ZN(n139) );
  OAI21_X1 U64 ( .B1(u_IE_i), .B2(irq_sec_ctrl_i), .A(n157), .ZN(n125) );
  NAND3_X1 U65 ( .A1(m_IE_i), .A2(current_priv_lvl_i[1]), .A3(
        current_priv_lvl_i[0]), .ZN(n124) );
  NAND2_X1 U66 ( .A1(n125), .A2(n124), .ZN(n152) );
  AND2_X1 U67 ( .A1(n152), .A2(irq_req_ctrl_i), .ZN(n230) );
  INV_X1 U68 ( .A(n230), .ZN(n184) );
  NOR2_X1 U69 ( .A1(n184), .A2(n101), .ZN(n143) );
  NOR2_X1 U70 ( .A1(illegal_insn_i), .A2(n143), .ZN(n180) );
  NAND4_X1 U71 ( .A1(n377), .A2(ctrl_fsm_cs[0]), .A3(n408), .A4(n413), .ZN(
        n126) );
  OR2_X1 U72 ( .A1(instr_valid_i), .A2(instr_valid_irq_flush_q), .ZN(n209) );
  NAND2_X1 U73 ( .A1(data_err_i_BAR), .A2(n209), .ZN(n160) );
  NOR2_X1 U74 ( .A1(n126), .A2(n160), .ZN(n127) );
  NOR2_X1 U75 ( .A1(n128), .A2(n409), .ZN(n136) );
  NOR2_X1 U76 ( .A1(n128), .A2(debug_req_i), .ZN(n135) );
  INV_X1 U77 ( .A(fencei_insn_i), .ZN(n130) );
  OAI21_X1 U78 ( .B1(n377), .B2(ctrl_fsm_cs[1]), .A(n311), .ZN(n129) );
  AOI21_X1 U79 ( .B1(n130), .B2(ctrl_fsm_cs[1]), .A(n129), .ZN(n131) );
  OAI21_X1 U80 ( .B1(n132), .B2(n408), .A(n131), .ZN(n133) );
  INV_X1 U81 ( .A(n133), .ZN(n134) );
  NOR3_X1 U82 ( .A1(n136), .A2(n135), .A3(n118), .ZN(n138) );
  OR2_X1 U83 ( .A1(ctrl_fsm_cs[2]), .A2(ctrl_fsm_cs[0]), .ZN(n206) );
  INV_X1 U84 ( .A(n206), .ZN(n295) );
  NOR2_X1 U85 ( .A1(ctrl_fsm_cs[1]), .A2(ctrl_fsm_cs[3]), .ZN(n294) );
  NAND3_X1 U86 ( .A1(n295), .A2(ctrl_fsm_cs[4]), .A3(n294), .ZN(n404) );
  INV_X1 U87 ( .A(n404), .ZN(n145) );
  AND2_X1 U88 ( .A1(n408), .A2(ctrl_fsm_cs[0]), .ZN(n401) );
  AND2_X1 U89 ( .A1(n401), .A2(n377), .ZN(n137) );
  INV_X1 U90 ( .A(data_err_i_BAR), .ZN(n417) );
  NAND2_X1 U91 ( .A1(n139), .A2(n209), .ZN(n140) );
  OR2_X1 U92 ( .A1(illegal_insn_i), .A2(n140), .ZN(n147) );
  INV_X1 U93 ( .A(n377), .ZN(n381) );
  INV_X1 U94 ( .A(n275), .ZN(n141) );
  INV_X1 U95 ( .A(n282), .ZN(n228) );
  INV_X1 U96 ( .A(n204), .ZN(n153) );
  NOR2_X1 U97 ( .A1(n153), .A2(n417), .ZN(n211) );
  INV_X1 U98 ( .A(n211), .ZN(n142) );
  INV_X1 U99 ( .A(dret_dec_i), .ZN(n144) );
  NOR2_X1 U100 ( .A1(n322), .A2(ctrl_fsm_cs[1]), .ZN(n231) );
  INV_X1 U101 ( .A(n403), .ZN(n350) );
  NAND2_X1 U102 ( .A1(n231), .A2(n350), .ZN(n199) );
  NAND2_X1 U103 ( .A1(n211), .A2(n101), .ZN(n146) );
  INV_X1 U104 ( .A(uret_insn_i), .ZN(n362) );
  OAI22_X1 U105 ( .A1(n147), .A2(n146), .B1(n199), .B2(n362), .ZN(n148) );
  NOR2_X1 U106 ( .A1(uret_insn_i), .A2(n199), .ZN(n150) );
  NAND2_X1 U107 ( .A1(n311), .A2(ctrl_fsm_cs[1]), .ZN(n227) );
  OR2_X1 U108 ( .A1(n227), .A2(n403), .ZN(n308) );
  NOR2_X1 U109 ( .A1(n308), .A2(n149), .ZN(n388) );
  AOI22_X1 U110 ( .A1(n150), .A2(mret_dec_i), .B1(fencei_insn_i), .B2(n388), 
        .ZN(n151) );
  NOR2_X1 U111 ( .A1(n322), .A2(n408), .ZN(n378) );
  AND2_X1 U112 ( .A1(n378), .A2(n350), .ZN(n383) );
  INV_X1 U113 ( .A(n383), .ZN(n380) );
  NAND2_X1 U114 ( .A1(n282), .A2(n350), .ZN(n158) );
  NAND2_X1 U115 ( .A1(n380), .A2(n158), .ZN(exc_pc_mux_o[1]) );
  AND2_X1 U116 ( .A1(irq_i), .A2(n152), .ZN(n235) );
  NOR3_X1 U117 ( .A1(n235), .A2(n417), .A3(n206), .ZN(n288) );
  AND3_X1 U118 ( .A1(n288), .A2(n350), .A3(n408), .ZN(instr_valid_irq_flush_n)
         );
  OR2_X1 U119 ( .A1(n103), .A2(data_err_i_BAR), .ZN(n271) );
  NOR2_X1 U120 ( .A1(n271), .A2(n153), .ZN(n187) );
  AND2_X1 U121 ( .A1(n275), .A2(ctrl_fsm_cs[1]), .ZN(n351) );
  INV_X1 U122 ( .A(n351), .ZN(n382) );
  OR2_X1 U123 ( .A1(n403), .A2(data_err_i_BAR), .ZN(n163) );
  AOI21_X1 U124 ( .B1(n382), .B2(n206), .A(n163), .ZN(n154) );
  AND2_X1 U125 ( .A1(current_priv_lvl_i[1]), .A2(current_priv_lvl_i[0]), .ZN(
        n155) );
  AND2_X1 U126 ( .A1(debug_ebreakm_i), .A2(n155), .ZN(n156) );
  AOI21_X1 U127 ( .B1(n157), .B2(debug_ebreaku_i), .A(n156), .ZN(n219) );
  INV_X1 U128 ( .A(ebrk_insn_i), .ZN(n407) );
  OR3_X1 U129 ( .A1(n219), .A2(n101), .A3(n407), .ZN(n159) );
  AOI21_X1 U130 ( .B1(n273), .B2(n159), .A(n158), .ZN(n376) );
  OR2_X1 U131 ( .A1(n376), .A2(n383), .ZN(debug_csr_save_o) );
  OAI21_X1 U132 ( .B1(n421), .B2(n230), .A(n409), .ZN(n326) );
  NAND2_X1 U133 ( .A1(n326), .A2(is_decoding_o), .ZN(n387) );
  INV_X1 U134 ( .A(n219), .ZN(n161) );
  NOR2_X1 U135 ( .A1(n161), .A2(n101), .ZN(n259) );
  AND2_X1 U136 ( .A1(n259), .A2(ebrk_insn_i), .ZN(n364) );
  NOR3_X1 U137 ( .A1(illegal_insn_i), .A2(n105), .A3(n364), .ZN(n162) );
  NOR2_X1 U138 ( .A1(n387), .A2(n162), .ZN(n375) );
  INV_X1 U139 ( .A(n196), .ZN(n286) );
  AND2_X1 U140 ( .A1(n206), .A2(n286), .ZN(n280) );
  OAI21_X1 U141 ( .B1(n163), .B2(n280), .A(csr_cause_o_5__BAR), .ZN(n164) );
  AND2_X1 U142 ( .A1(n410), .A2(ctrl_fsm_cs[1]), .ZN(n239) );
  NAND2_X1 U143 ( .A1(n239), .A2(n309), .ZN(n341) );
  NOR2_X1 U144 ( .A1(n237), .A2(n341), .ZN(n279) );
  NOR2_X1 U145 ( .A1(n206), .A2(n408), .ZN(n241) );
  NAND2_X1 U146 ( .A1(n165), .A2(n350), .ZN(n166) );
  OR4_X1 U147 ( .A1(n279), .A2(n241), .A3(n351), .A4(n166), .ZN(
        exc_pc_mux_o[0]) );
  NAND2_X1 U148 ( .A1(regfile_alu_we_fw_i), .A2(reg_d_alu_is_reg_b_i), .ZN(
        n405) );
  INV_X1 U149 ( .A(data_misaligned_i), .ZN(n358) );
  AND4_X1 U150 ( .A1(regfile_we_wb_i), .A2(reg_d_wb_is_reg_b_i), .A3(n405), 
        .A4(n358), .ZN(operand_b_fw_mux_sel_o[1]) );
  AOI22_X1 U151 ( .A1(regfile_alu_we_fw_i), .A2(reg_d_alu_is_reg_c_i), .B1(
        mult_multicycle_i), .B2(n358), .ZN(operand_c_fw_mux_sel_o_0__BAR) );
  AND3_X1 U152 ( .A1(regfile_we_wb_i), .A2(operand_c_fw_mux_sel_o_0__BAR), 
        .A3(reg_d_wb_is_reg_c_i), .ZN(operand_c_fw_mux_sel_o_1_) );
  AND2_X1 U153 ( .A1(n231), .A2(n377), .ZN(first_fetch_o) );
  INV_X1 U154 ( .A(regfile_we_wb_i), .ZN(n167) );
  OR2_X1 U155 ( .A1(wb_ready_i), .A2(n167), .ZN(n178) );
  NAND2_X1 U156 ( .A1(regfile_we_ex_i), .A2(data_req_ex_i), .ZN(n177) );
  INV_X1 U157 ( .A(is_decoding_o), .ZN(is_decoding_o_BAR) );
  XOR2_X1 U158 ( .A(regfile_alu_waddr_id_i[1]), .B(regfile_waddr_ex_i[1]), .Z(
        n173) );
  XOR2_X1 U159 ( .A(regfile_alu_waddr_id_i[4]), .B(regfile_waddr_ex_i[4]), .Z(
        n172) );
  XNOR2_X1 U160 ( .A(regfile_alu_waddr_id_i[3]), .B(regfile_waddr_ex_i[3]), 
        .ZN(n170) );
  XNOR2_X1 U161 ( .A(regfile_alu_waddr_id_i[2]), .B(regfile_waddr_ex_i[2]), 
        .ZN(n169) );
  XNOR2_X1 U162 ( .A(regfile_alu_waddr_id_i[0]), .B(regfile_waddr_ex_i[0]), 
        .ZN(n168) );
  NAND4_X1 U163 ( .A1(n170), .A2(n169), .A3(n168), .A4(regfile_we_id_i), .ZN(
        n171) );
  NOR4_X1 U164 ( .A1(is_decoding_o_BAR), .A2(n173), .A3(n172), .A4(n171), .ZN(
        n174) );
  NOR3_X1 U165 ( .A1(n174), .A2(reg_d_ex_is_reg_a_i), .A3(reg_d_ex_is_reg_b_i), 
        .ZN(n176) );
  INV_X1 U166 ( .A(reg_d_ex_is_reg_c_i), .ZN(n175) );
  AND2_X1 U167 ( .A1(mret_insn_i), .A2(n388), .ZN(csr_restore_mret_id_o) );
  INV_X1 U168 ( .A(csr_cause_o_5__BAR), .ZN(n372) );
  AND2_X1 U169 ( .A1(n372), .A2(irq_id_ctrl_i[4]), .ZN(\exc_cause_o[4] ) );
  NAND2_X1 U170 ( .A1(n239), .A2(n377), .ZN(ctrl_busy_o) );
  AND2_X1 U171 ( .A1(n273), .A2(n180), .ZN(n327) );
  NOR2_X1 U172 ( .A1(mret_insn_i), .A2(uret_insn_i), .ZN(n221) );
  INV_X1 U173 ( .A(n221), .ZN(n181) );
  NOR2_X1 U174 ( .A1(n181), .A2(dret_insn_i), .ZN(n342) );
  NOR3_X1 U175 ( .A1(n237), .A2(fencei_insn_i), .A3(pipe_flush_i), .ZN(n182)
         );
  AND2_X1 U176 ( .A1(n342), .A2(n182), .ZN(n258) );
  AOI21_X1 U177 ( .B1(n327), .B2(n258), .A(is_decoding_o_BAR), .ZN(n191) );
  AND2_X1 U178 ( .A1(n273), .A2(n184), .ZN(n205) );
  INV_X1 U179 ( .A(first_fetch_o), .ZN(n189) );
  OR2_X1 U180 ( .A1(n403), .A2(n310), .ZN(n185) );
  OAI21_X1 U181 ( .B1(n378), .B2(n185), .A(ctrl_busy_o), .ZN(n186) );
  NOR2_X1 U182 ( .A1(n187), .A2(n186), .ZN(n188) );
  OAI21_X1 U183 ( .B1(n205), .B2(n189), .A(n188), .ZN(n190) );
  NOR4_X1 U184 ( .A1(n351), .A2(n294), .A3(ctrl_fsm_cs[4]), .A4(n410), .ZN(
        n192) );
  AND4_X1 U185 ( .A1(n193), .A2(dret_dec_i), .A3(n192), .A4(csr_cause_o_5__BAR), .ZN(n195) );
  INV_X1 U186 ( .A(exc_pc_mux_o[1]), .ZN(n194) );
  OAI21_X1 U187 ( .B1(n195), .B2(n409), .A(n194), .ZN(n267) );
  NAND3_X1 U188 ( .A1(n326), .A2(n270), .A3(illegal_insn_i), .ZN(n202) );
  MUX2_X1 U189 ( .A(n412), .B(n350), .S(n275), .Z(n197) );
  NOR3_X1 U190 ( .A1(n403), .A2(ctrl_fsm_cs[1]), .A3(ctrl_fsm_cs[2]), .ZN(n349) );
  NOR4_X1 U191 ( .A1(n197), .A2(n349), .A3(ctrl_fsm_cs[4]), .A4(n196), .ZN(
        n200) );
  NOR2_X1 U192 ( .A1(n417), .A2(n403), .ZN(n318) );
  NAND2_X1 U193 ( .A1(n318), .A2(n241), .ZN(n216) );
  INV_X1 U194 ( .A(n308), .ZN(n198) );
  NAND2_X1 U195 ( .A1(n198), .A2(data_err_q), .ZN(n393) );
  NAND4_X1 U196 ( .A1(n200), .A2(n216), .A3(n199), .A4(n393), .ZN(n201) );
  AOI21_X1 U197 ( .B1(n202), .B2(n204), .A(n201), .ZN(n203) );
  MUX2_X1 U198 ( .A(illegal_insn_q), .B(n204), .S(n203), .Z(n269) );
  NAND3_X1 U199 ( .A1(id_ready_i_BAR), .A2(n205), .A3(first_fetch_o), .ZN(n215) );
  NOR4_X1 U200 ( .A1(n421), .A2(irq_i), .A3(n101), .A4(debug_single_step_i), 
        .ZN(n208) );
  AOI211_X1 U201 ( .C1(fetch_enable_i), .C2(n408), .A(n381), .B(n206), .ZN(
        n207) );
  OAI21_X1 U202 ( .B1(n208), .B2(n408), .A(n207), .ZN(n213) );
  INV_X1 U203 ( .A(n209), .ZN(n210) );
  NAND2_X1 U204 ( .A1(n211), .A2(n210), .ZN(n346) );
  AND3_X1 U205 ( .A1(n213), .A2(n212), .A3(n346), .ZN(n214) );
  OAI211_X1 U206 ( .C1(ex_valid_i), .C2(n216), .A(n215), .B(n214), .ZN(n321)
         );
  INV_X1 U207 ( .A(n321), .ZN(n252) );
  NAND2_X1 U208 ( .A1(n409), .A2(debug_single_step_i), .ZN(n283) );
  NOR2_X1 U209 ( .A1(id_ready_i_BAR), .A2(n283), .ZN(n255) );
  INV_X1 U210 ( .A(n255), .ZN(n324) );
  INV_X1 U211 ( .A(illegal_insn_i), .ZN(n367) );
  NAND3_X1 U212 ( .A1(id_ready_i_BAR), .A2(n258), .A3(n367), .ZN(n217) );
  NAND2_X1 U213 ( .A1(n324), .A2(n217), .ZN(n325) );
  INV_X1 U214 ( .A(n258), .ZN(n218) );
  NOR3_X1 U215 ( .A1(illegal_insn_i), .A2(csr_status_i), .A3(n218), .ZN(n224)
         );
  NAND2_X1 U216 ( .A1(jump_in_id_i[1]), .A2(jump_in_id_i[0]), .ZN(n323) );
  AOI21_X1 U217 ( .B1(n219), .B2(ebrk_insn_i), .A(n105), .ZN(n220) );
  NAND2_X1 U218 ( .A1(n221), .A2(n220), .ZN(n222) );
  NOR2_X1 U219 ( .A1(illegal_insn_i), .A2(n222), .ZN(n254) );
  INV_X1 U220 ( .A(n254), .ZN(n223) );
  OAI21_X1 U221 ( .B1(n323), .B2(n223), .A(n255), .ZN(n333) );
  OAI21_X1 U222 ( .B1(n325), .B2(n224), .A(n333), .ZN(n225) );
  INV_X1 U223 ( .A(n273), .ZN(n305) );
  AOI21_X1 U224 ( .B1(n225), .B2(n326), .A(n305), .ZN(n226) );
  NAND2_X1 U225 ( .A1(n270), .A2(n282), .ZN(n332) );
  OR2_X1 U226 ( .A1(n226), .A2(n332), .ZN(n233) );
  INV_X1 U227 ( .A(n227), .ZN(n229) );
  INV_X1 U228 ( .A(n231), .ZN(n303) );
  OAI22_X1 U229 ( .A1(n273), .A2(n303), .B1(n228), .B2(n271), .ZN(n335) );
  AOI211_X1 U230 ( .C1(n231), .C2(n230), .A(n229), .B(n335), .ZN(n232) );
  AOI21_X1 U231 ( .B1(n233), .B2(n232), .A(ctrl_fsm_cs[4]), .ZN(n250) );
  NAND3_X1 U232 ( .A1(n305), .A2(n311), .A3(n408), .ZN(n234) );
  NOR2_X1 U233 ( .A1(id_ready_i_BAR), .A2(n234), .ZN(n249) );
  OAI21_X1 U234 ( .B1(n235), .B2(n417), .A(n295), .ZN(n247) );
  INV_X1 U235 ( .A(n237), .ZN(n238) );
  AOI21_X1 U236 ( .B1(n238), .B2(n415), .A(data_err_q), .ZN(n277) );
  NAND2_X1 U237 ( .A1(n277), .A2(n239), .ZN(n240) );
  NAND2_X1 U238 ( .A1(n240), .A2(n303), .ZN(n243) );
  INV_X1 U239 ( .A(n283), .ZN(n356) );
  OR2_X1 U240 ( .A1(n241), .A2(n412), .ZN(n242) );
  AOI21_X1 U241 ( .B1(n243), .B2(n356), .A(n242), .ZN(n340) );
  INV_X1 U242 ( .A(n341), .ZN(n244) );
  NAND2_X1 U243 ( .A1(pipe_flush_i), .A2(n244), .ZN(n246) );
  NOR2_X1 U244 ( .A1(data_load_event_i), .A2(n283), .ZN(n287) );
  OAI21_X1 U245 ( .B1(n287), .B2(n417), .A(n351), .ZN(n245) );
  NAND4_X1 U246 ( .A1(n247), .A2(n340), .A3(n246), .A4(n245), .ZN(n248) );
  OAI22_X1 U247 ( .A1(n250), .A2(n350), .B1(n249), .B2(n248), .ZN(n251) );
  OAI211_X1 U248 ( .C1(n252), .C2(n408), .A(n251), .B(n404), .ZN(n266) );
  AOI21_X1 U249 ( .B1(id_ready_i_BAR), .B2(csr_status_i), .A(data_load_event_i), .ZN(n272) );
  NAND2_X1 U250 ( .A1(n327), .A2(n270), .ZN(n253) );
  NOR2_X1 U251 ( .A1(n255), .A2(n253), .ZN(n261) );
  INV_X1 U252 ( .A(n261), .ZN(n300) );
  NAND4_X1 U253 ( .A1(n255), .A2(n254), .A3(n326), .A4(n323), .ZN(n256) );
  NAND2_X1 U254 ( .A1(n256), .A2(n273), .ZN(n262) );
  NOR2_X1 U255 ( .A1(csr_status_i), .A2(data_load_event_i), .ZN(n354) );
  NAND2_X1 U256 ( .A1(n354), .A2(n258), .ZN(n329) );
  OAI211_X1 U257 ( .C1(n259), .C2(n407), .A(n329), .B(n396), .ZN(n260) );
  AOI22_X1 U258 ( .A1(n270), .A2(n262), .B1(n261), .B2(n260), .ZN(n299) );
  OAI211_X1 U259 ( .C1(n272), .C2(n300), .A(n299), .B(n271), .ZN(n276) );
  INV_X1 U260 ( .A(n322), .ZN(n274) );
  AOI22_X1 U261 ( .A1(n276), .A2(n275), .B1(n274), .B2(n273), .ZN(n297) );
  OAI21_X1 U262 ( .B1(id_ready_i_BAR), .B2(n305), .A(n401), .ZN(n292) );
  AOI21_X1 U263 ( .B1(n277), .B2(n283), .A(data_err_q), .ZN(n278) );
  OAI21_X1 U264 ( .B1(n278), .B2(ctrl_fsm_cs[2]), .A(ctrl_fsm_cs[0]), .ZN(n290) );
  NAND2_X1 U265 ( .A1(n342), .A2(n279), .ZN(n285) );
  NOR2_X1 U266 ( .A1(n280), .A2(data_err_i_BAR), .ZN(n281) );
  AOI211_X1 U267 ( .C1(n310), .C2(n283), .A(n282), .B(n281), .ZN(n284) );
  OAI211_X1 U268 ( .C1(n287), .C2(n286), .A(n285), .B(n284), .ZN(n289) );
  AOI211_X1 U269 ( .C1(ctrl_fsm_cs[1]), .C2(n290), .A(n289), .B(n288), .ZN(
        n291) );
  AOI21_X1 U270 ( .B1(n292), .B2(n291), .A(n403), .ZN(n293) );
  AOI211_X1 U271 ( .C1(n295), .C2(n294), .A(n372), .B(n293), .ZN(n296) );
  OAI21_X1 U272 ( .B1(n297), .B2(n381), .A(n296), .ZN(n298) );
  MUX2_X1 U273 ( .A(n298), .B(ctrl_fsm_cs[0]), .S(n321), .Z(n263) );
  INV_X1 U274 ( .A(n299), .ZN(n302) );
  INV_X1 U275 ( .A(id_ready_i_BAR), .ZN(n400) );
  NOR3_X1 U276 ( .A1(n300), .A2(n354), .A3(n400), .ZN(n301) );
  OAI21_X1 U277 ( .B1(n302), .B2(n301), .A(n310), .ZN(n304) );
  AOI21_X1 U278 ( .B1(n304), .B2(n303), .A(ctrl_fsm_cs[4]), .ZN(n317) );
  NAND4_X1 U279 ( .A1(n400), .A2(n305), .A3(ctrl_fsm_cs[0]), .A4(n350), .ZN(
        n307) );
  AOI22_X1 U280 ( .A1(n318), .A2(n414), .B1(n377), .B2(n311), .ZN(n306) );
  AOI21_X1 U281 ( .B1(n307), .B2(n306), .A(ctrl_fsm_cs[1]), .ZN(n316) );
  AOI21_X1 U282 ( .B1(pipe_flush_i), .B2(n309), .A(n308), .ZN(n315) );
  INV_X1 U283 ( .A(n310), .ZN(n313) );
  INV_X1 U284 ( .A(n311), .ZN(n337) );
  NAND3_X1 U285 ( .A1(n337), .A2(ctrl_fsm_cs[1]), .A3(n377), .ZN(n312) );
  OAI211_X1 U286 ( .C1(n313), .C2(n403), .A(n404), .B(n312), .ZN(n314) );
  NOR4_X1 U287 ( .A1(n317), .A2(n316), .A3(n315), .A4(n314), .ZN(n320) );
  NOR2_X1 U288 ( .A1(n321), .A2(n318), .ZN(n319) );
  OAI222_X1 U289 ( .A1(n403), .A2(n322), .B1(n321), .B2(n320), .C1(n410), .C2(
        n319), .ZN(n265) );
  NOR3_X1 U290 ( .A1(n324), .A2(n323), .A3(n387), .ZN(n264) );
  INV_X1 U291 ( .A(n325), .ZN(n331) );
  INV_X1 U292 ( .A(n326), .ZN(n330) );
  INV_X1 U293 ( .A(n327), .ZN(n328) );
  OAI22_X1 U294 ( .A1(n331), .A2(n330), .B1(n329), .B2(n328), .ZN(n334) );
  AOI21_X1 U295 ( .B1(n334), .B2(n333), .A(n332), .ZN(n336) );
  NOR3_X1 U296 ( .A1(n336), .A2(ctrl_fsm_cs[3]), .A3(n335), .ZN(n345) );
  OAI21_X1 U297 ( .B1(ctrl_fsm_cs[2]), .B2(data_err_i_BAR), .A(n337), .ZN(n338) );
  AOI21_X1 U298 ( .B1(n338), .B2(n408), .A(n351), .ZN(n339) );
  OAI211_X1 U299 ( .C1(n342), .C2(n341), .A(n340), .B(n339), .ZN(n343) );
  NAND2_X1 U300 ( .A1(n343), .A2(n411), .ZN(n344) );
  OAI21_X1 U301 ( .B1(n345), .B2(n344), .A(n404), .ZN(n268) );
  NOR2_X1 U302 ( .A1(n103), .A2(n346), .ZN(n348) );
  AOI211_X1 U303 ( .C1(n351), .C2(n350), .A(n349), .B(n348), .ZN(n353) );
  INV_X1 U304 ( .A(data_load_event_i), .ZN(n352) );
  NOR2_X1 U305 ( .A1(n353), .A2(n352), .ZN(perf_pipeline_stall_o) );
  INV_X1 U306 ( .A(n354), .ZN(n355) );
  OAI21_X1 U307 ( .B1(n356), .B2(n355), .A(is_decoding_o), .ZN(n357) );
  NAND3_X1 U308 ( .A1(halt_id_o_BAR), .A2(n404), .A3(n357), .ZN(halt_if_o) );
  NAND2_X1 U309 ( .A1(n359), .A2(n358), .ZN(operand_a_fw_mux_sel_o[0]) );
  NOR2_X1 U310 ( .A1(operand_a_fw_mux_sel_o[0]), .A2(n360), .ZN(
        operand_a_fw_mux_sel_o[1]) );
  AND2_X1 U311 ( .A1(dret_insn_i), .A2(n388), .ZN(csr_restore_dret_id_o) );
  INV_X1 U312 ( .A(n388), .ZN(n361) );
  NOR2_X1 U313 ( .A1(n362), .A2(n361), .ZN(csr_restore_uret_id_o) );
  INV_X1 U314 ( .A(irq_sec_ctrl_i), .ZN(n363) );
  NOR2_X1 U315 ( .A1(csr_cause_o_5__BAR), .A2(n363), .ZN(csr_irq_sec_o) );
  NOR2_X1 U316 ( .A1(n387), .A2(illegal_insn_i), .ZN(n398) );
  INV_X1 U317 ( .A(n398), .ZN(n374) );
  AOI21_X1 U318 ( .B1(n105), .B2(n365), .A(n364), .ZN(n368) );
  NAND2_X1 U319 ( .A1(n372), .A2(irq_id_ctrl_i[0]), .ZN(n389) );
  OAI211_X1 U321 ( .C1(n374), .C2(n368), .A(csr_save_ex_o_BAR), .B(n389), .ZN(
        csr_cause_o_0_) );
  INV_X1 U322 ( .A(csr_save_ex_o_BAR), .ZN(n370) );
  INV_X1 U323 ( .A(irq_id_ctrl_i[1]), .ZN(n366) );
  NOR2_X1 U324 ( .A1(csr_cause_o_5__BAR), .A2(n366), .ZN(n390) );
  AOI21_X1 U325 ( .B1(n368), .B2(n367), .A(n387), .ZN(n369) );
  AOI211_X1 U326 ( .C1(data_we_ex_i), .C2(n370), .A(n390), .B(n369), .ZN(
        csr_cause_o_1__BAR) );
  NAND2_X1 U327 ( .A1(n372), .A2(irq_id_ctrl_i[2]), .ZN(n392) );
  NAND2_X1 U328 ( .A1(csr_save_ex_o_BAR), .A2(n392), .ZN(csr_cause_o_2_) );
  INV_X1 U329 ( .A(n105), .ZN(n373) );
  NAND2_X1 U330 ( .A1(n372), .A2(irq_id_ctrl_i[3]), .ZN(n394) );
  OAI21_X1 U331 ( .B1(n374), .B2(n373), .A(n394), .ZN(csr_cause_o_3_) );
  AOI211_X1 U332 ( .C1(n378), .C2(n377), .A(n376), .B(n375), .ZN(n379) );
  INV_X1 U333 ( .A(n379), .ZN(csr_save_id_o) );
  OAI21_X1 U334 ( .B1(n382), .B2(n381), .A(n380), .ZN(csr_save_if_o) );
  NAND3_X1 U335 ( .A1(n407), .A2(n383), .A3(debug_single_step_i), .ZN(n384) );
  NOR2_X1 U336 ( .A1(n421), .A2(n384), .ZN(debug_cause_o[2]) );
  INV_X1 U337 ( .A(irq_req_ctrl_i), .ZN(n386) );
  INV_X1 U338 ( .A(instr_valid_irq_flush_n), .ZN(n385) );
  OAI21_X1 U339 ( .B1(n387), .B2(n386), .A(n385), .ZN(exc_kill_o) );
  NAND2_X1 U340 ( .A1(n105), .A2(n388), .ZN(n395) );
  NAND3_X1 U341 ( .A1(n395), .A2(n393), .A3(n389), .ZN(exc_cause_o[0]) );
  INV_X1 U342 ( .A(n390), .ZN(n391) );
  OAI211_X1 U343 ( .C1(data_we_ex_i), .C2(n393), .A(n395), .B(n391), .ZN(
        exc_cause_o[1]) );
  NAND2_X1 U344 ( .A1(n393), .A2(n392), .ZN(exc_cause_o[2]) );
  NAND2_X1 U345 ( .A1(n395), .A2(n394), .ZN(exc_cause_o[3]) );
  NOR2_X1 U346 ( .A1(jr_stall_o), .A2(n396), .ZN(n397) );
  AOI21_X1 U347 ( .B1(n398), .B2(n397), .A(jump_done_q), .ZN(n399) );
  NOR2_X1 U348 ( .A1(n400), .A2(n399), .ZN(N448) );
  OAI21_X1 U349 ( .B1(n401), .B2(ctrl_fsm_cs[2]), .A(n411), .ZN(n402) );
  NAND3_X1 U350 ( .A1(n404), .A2(n403), .A3(n402), .ZN(instr_req_o) );
  XOR2_X1 U351 ( .A(jump_in_id_i[0]), .B(jump_in_id_i[1]), .Z(perf_jump_o) );
  NOR2_X1 U352 ( .A1(data_misaligned_i), .A2(n405), .ZN(
        operand_b_fw_mux_sel_o[0]) );
  AND3_X1 U353 ( .A1(n407), .A2(debug_csr_save_o), .A3(n421), .ZN(
        debug_cause_o[1]) );
  SDFFR_X1 data_err_q_reg ( .D(n417), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(data_err_q) );
  SDFFR_X1 illegal_insn_q_reg ( .D(n269), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(illegal_insn_q), .QN(n415) );
  SDFFR_X1 ctrl_fsm_cs_reg_4_ ( .D(n264), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(ctrl_fsm_cs[4]), .QN(n411) );
  SDFFR_X1 ctrl_fsm_cs_reg_3_ ( .D(n268), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(ctrl_fsm_cs[3]), .QN(n412) );
  SDFFR_X1 instr_valid_irq_flush_q_reg ( .D(instr_valid_irq_flush_n), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(rst_n), .Q(instr_valid_irq_flush_q) );
  SDFFR_X1 ctrl_fsm_cs_reg_0_ ( .D(n263), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(ctrl_fsm_cs[0]), .QN(n414) );
  SDFFR_X1 ctrl_fsm_cs_reg_2_ ( .D(n265), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(ctrl_fsm_cs[2]), .QN(n410) );
  SDFFR_X1 ctrl_fsm_cs_reg_1_ ( .D(n266), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(ctrl_fsm_cs[1]), .QN(n408) );
  SDFFR_X1 debug_mode_q_reg ( .D(n267), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(n101), .QN(n409) );
  SDFFR_X1 jump_done_q_reg ( .D(N448), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(jump_done_q), .QN(n413) );
  NOR3_X1 U3 ( .A1(csr_cause_o_5__BAR), .A2(irq_sec_ctrl_i), .A3(n365), .ZN(
        trap_addr_mux_o) );
  CLKBUF_X1 U10 ( .A(n347), .Z(n103) );
  OR4_X1 U31 ( .A1(debug_csr_save_o), .A2(n187), .A3(n375), .A4(n164), .ZN(
        csr_save_cause_o) );
  BUF_X1 U6 ( .A(debug_req_i), .Z(n421) );
  NAND2_X1 U11 ( .A1(n421), .A2(n409), .ZN(n273) );
  NOR2_X1 U16 ( .A1(n347), .A2(n160), .ZN(n270) );
  NOR2_X2 U26 ( .A1(n187), .A2(n154), .ZN(csr_save_ex_o_BAR) );
  CLKBUF_X1 U30 ( .A(branch_taken_ex_i), .Z(n347) );
  NAND3_X1 U355 ( .A1(n179), .A2(n180), .A3(n110), .ZN(n128) );
endmodule



    module riscv_decoder_FPU0_FP_DIVSQRT0_PULP_SECURE1_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_WOP_CPU6 ( 
        deassert_we_i, data_misaligned_i, mult_multicycle_i, 
        instr_multicycle_o, illegal_insn_o, ebrk_insn_o, mret_insn_o, 
        uret_insn_o, dret_insn_o, mret_dec_o, uret_dec_o, dret_dec_o, 
        ecall_insn_o, pipe_flush_o, fencei_insn_o, rega_used_o, regb_used_o, 
        regc_used_o, reg_fp_a_o, reg_fp_b_o, reg_fp_c_o, reg_fp_d_o, 
        bmask_a_mux_o, bmask_b_mux_o, alu_bmask_a_mux_sel_o, 
        alu_bmask_b_mux_sel_o, instr_rdata_i, illegal_c_insn_i, alu_en_o, 
        alu_operator_o, alu_op_a_mux_sel_o, alu_op_b_mux_sel_o, 
        alu_op_c_mux_sel_o, alu_vec_mode_o, scalar_replication_o, 
        scalar_replication_c_o, imm_a_mux_sel_o, imm_b_mux_sel_o, regc_mux_o, 
        is_clpx_o, is_subrot_o, mult_operator_o, mult_int_en_o, mult_dot_en_o, 
        mult_sel_subword_o, mult_signed_mode_o, mult_dot_signed_o, frm_i, 
        fpu_dst_fmt_o, fpu_src_fmt_o, fpu_int_fmt_o, apu_en_o, apu_type_o, 
        apu_op_o, apu_lat_o, apu_flags_src_o, fp_rnd_mode_o, regfile_mem_we_o, 
        regfile_alu_we_o, regfile_alu_we_dec_o, regfile_alu_waddr_sel_o, 
        csr_access_o, csr_status_o, csr_op_o, current_priv_lvl_i, data_req_o, 
        data_we_o, prepost_useincr_o, data_type_o, data_sign_extension_o, 
        data_reg_offset_o, data_load_event_o, hwloop_we_o, 
        hwloop_target_mux_sel_o, hwloop_start_mux_sel_o, hwloop_cnt_mux_sel_o, 
        jump_in_dec_o, jump_in_id_o, jump_target_mux_sel_o, 
        \mult_imm_mux_o[0]_BAR  );
  output [0:0] bmask_a_mux_o;
  output [1:0] bmask_b_mux_o;
  input [31:0] instr_rdata_i;
  output [6:0] alu_operator_o;
  output [2:0] alu_op_a_mux_sel_o;
  output [2:0] alu_op_b_mux_sel_o;
  output [1:0] alu_op_c_mux_sel_o;
  output [1:0] alu_vec_mode_o;
  output [0:0] imm_a_mux_sel_o;
  output [3:0] imm_b_mux_sel_o;
  output [1:0] regc_mux_o;
  output [2:0] mult_operator_o;
  output [1:0] mult_signed_mode_o;
  output [1:0] mult_dot_signed_o;
  input [2:0] frm_i;
  output [2:0] fpu_dst_fmt_o;
  output [2:0] fpu_src_fmt_o;
  output [1:0] fpu_int_fmt_o;
  output [1:2] apu_type_o;
  output [5:0] apu_op_o;
  output [1:0] apu_lat_o;
  output [1:2] apu_flags_src_o;
  output [2:0] fp_rnd_mode_o;
  output [1:0] csr_op_o;
  input [1:0] current_priv_lvl_i;
  output [1:0] data_type_o;
  output [1:0] data_sign_extension_o;
  output [1:0] data_reg_offset_o;
  output [2:0] hwloop_we_o;
  output [1:0] jump_in_dec_o;
  output [1:0] jump_in_id_o;
  output [1:0] jump_target_mux_sel_o;
  input deassert_we_i, data_misaligned_i, mult_multicycle_i, illegal_c_insn_i;
  output instr_multicycle_o, illegal_insn_o, ebrk_insn_o, mret_insn_o,
         uret_insn_o, dret_insn_o, mret_dec_o, uret_dec_o, dret_dec_o,
         ecall_insn_o, pipe_flush_o, fencei_insn_o, rega_used_o, regb_used_o,
         regc_used_o, reg_fp_a_o, reg_fp_b_o, reg_fp_c_o, reg_fp_d_o,
         alu_bmask_a_mux_sel_o, alu_bmask_b_mux_sel_o, alu_en_o,
         scalar_replication_o, scalar_replication_c_o, is_clpx_o, is_subrot_o,
         mult_int_en_o, mult_dot_en_o, mult_sel_subword_o, apu_en_o,
         regfile_mem_we_o, regfile_alu_we_o, regfile_alu_we_dec_o,
         regfile_alu_waddr_sel_o, csr_access_o, csr_status_o, data_req_o,
         data_we_o, prepost_useincr_o, data_load_event_o,
         hwloop_target_mux_sel_o, hwloop_start_mux_sel_o, hwloop_cnt_mux_sel_o,
         \mult_imm_mux_o[0]_BAR ;
  wire   n590, \mult_imm_mux_o[0] , n14, n17, n18, n19, n20, n21, n22, n25,
         n26, n27, n28, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n591, n592, n593, n594, n595, n596, n597, n598;
  assign \mult_imm_mux_o[0]_BAR  = n282;

  NOR2_X1 U4 ( .A1(n48), .A2(n225), .ZN(hwloop_cnt_mux_sel_o) );
  NAND3_X1 U5 ( .A1(n43), .A2(n232), .A3(n231), .ZN(rega_used_o) );
  INV_X1 U6 ( .A(n14), .ZN(n41) );
  OAI21_X1 U7 ( .B1(n230), .B2(n28), .A(n507), .ZN(n14) );
  AND2_X1 U9 ( .A1(instr_rdata_i[12]), .A2(n558), .ZN(n356) );
  NOR2_X1 U13 ( .A1(n157), .A2(n545), .ZN(n17) );
  NOR2_X1 U14 ( .A1(n157), .A2(n545), .ZN(n441) );
  OR2_X2 U15 ( .A1(n485), .A2(n50), .ZN(jump_target_mux_sel_o[0]) );
  INV_X1 U16 ( .A(instr_rdata_i[3]), .ZN(n18) );
  INV_X1 U17 ( .A(instr_rdata_i[3]), .ZN(n19) );
  CLKBUF_X1 U20 ( .A(n590), .Z(bmask_a_mux_o[0]) );
  CLKBUF_X1 U21 ( .A(n491), .Z(n38) );
  NOR2_X1 U22 ( .A1(n20), .A2(instr_rdata_i[31]), .ZN(n27) );
  AOI211_X2 U23 ( .C1(n208), .C2(n82), .A(n558), .B(n79), .ZN(
        scalar_replication_o) );
  NOR4_X1 U24 ( .A1(n435), .A2(n501), .A3(n300), .A4(n375), .ZN(n176) );
  NOR2_X1 U27 ( .A1(n228), .A2(n227), .ZN(n590) );
  OR2_X1 U28 ( .A1(n25), .A2(n242), .ZN(n230) );
  AND2_X1 U29 ( .A1(n314), .A2(n507), .ZN(n516) );
  OR2_X1 U30 ( .A1(n533), .A2(n575), .ZN(n572) );
  INV_X1 U31 ( .A(n551), .ZN(n28) );
  OR2_X1 U32 ( .A1(n197), .A2(n575), .ZN(n559) );
  OR2_X1 U34 ( .A1(n416), .A2(n575), .ZN(n491) );
  AND2_X1 U35 ( .A1(n288), .A2(instr_rdata_i[13]), .ZN(n481) );
  INV_X1 U38 ( .A(n395), .ZN(n157) );
  INV_X1 U40 ( .A(n93), .ZN(n20) );
  INV_X1 U41 ( .A(instr_rdata_i[3]), .ZN(n233) );
  NAND2_X1 U42 ( .A1(n491), .A2(jump_target_mux_sel_o[0]), .ZN(
        jump_target_mux_sel_o[1]) );
  NAND3_X1 U44 ( .A1(n148), .A2(n22), .A3(n21), .ZN(n35) );
  INV_X1 U45 ( .A(n147), .ZN(n21) );
  NAND2_X1 U46 ( .A1(n415), .A2(instr_rdata_i[27]), .ZN(n22) );
  NOR2_X2 U47 ( .A1(instr_rdata_i[29]), .A2(instr_rdata_i[28]), .ZN(n360) );
  NAND2_X1 U48 ( .A1(n488), .A2(n26), .ZN(n25) );
  AND2_X1 U49 ( .A1(n192), .A2(n483), .ZN(n26) );
  NAND2_X1 U50 ( .A1(n88), .A2(n93), .ZN(n355) );
  NAND2_X1 U51 ( .A1(n88), .A2(n27), .ZN(n551) );
  AND2_X1 U52 ( .A1(n488), .A2(n192), .ZN(n229) );
  NAND2_X1 U53 ( .A1(n533), .A2(n539), .ZN(n242) );
  NOR2_X1 U54 ( .A1(n49), .A2(instr_rdata_i[4]), .ZN(n30) );
  NOR2_X1 U55 ( .A1(n49), .A2(instr_rdata_i[4]), .ZN(n191) );
  OR2_X2 U57 ( .A1(instr_rdata_i[26]), .A2(instr_rdata_i[27]), .ZN(n76) );
  NOR2_X2 U58 ( .A1(n76), .A2(instr_rdata_i[25]), .ZN(n333) );
  INV_X1 U59 ( .A(instr_rdata_i[14]), .ZN(n395) );
  NAND2_X1 U60 ( .A1(n289), .A2(n558), .ZN(n487) );
  OR2_X1 U61 ( .A1(n193), .A2(n575), .ZN(n225) );
  OR2_X1 U62 ( .A1(n338), .A2(n184), .ZN(n44) );
  AND2_X1 U63 ( .A1(n390), .A2(n378), .ZN(n48) );
  NOR2_X1 U65 ( .A1(data_misaligned_i), .A2(n99), .ZN(alu_op_a_mux_sel_o[2])
         );
  AND2_X1 U66 ( .A1(instr_rdata_i[4]), .A2(instr_rdata_i[5]), .ZN(n51) );
  OAI21_X1 U67 ( .B1(n123), .B2(n487), .A(n36), .ZN(n170) );
  INV_X1 U68 ( .A(n44), .ZN(n47) );
  NOR3_X1 U69 ( .A1(n225), .A2(instr_rdata_i[13]), .A3(n558), .ZN(
        hwloop_start_mux_sel_o) );
  NOR2_X1 U70 ( .A1(n414), .A2(n595), .ZN(n214) );
  AND2_X1 U71 ( .A1(instr_rdata_i[6]), .A2(instr_rdata_i[2]), .ZN(n55) );
  NOR3_X1 U72 ( .A1(n246), .A2(n381), .A3(n40), .ZN(n39) );
  INV_X1 U73 ( .A(n507), .ZN(n40) );
  AOI21_X1 U74 ( .B1(n579), .B2(n584), .A(n586), .ZN(n122) );
  INV_X1 U75 ( .A(n37), .ZN(n36) );
  OAI21_X1 U76 ( .B1(n262), .B2(n245), .A(n326), .ZN(n37) );
  INV_X1 U77 ( .A(n325), .ZN(n322) );
  NOR2_X1 U78 ( .A1(instr_rdata_i[13]), .A2(instr_rdata_i[12]), .ZN(n289) );
  INV_X1 U80 ( .A(n575), .ZN(n507) );
  NOR3_X1 U81 ( .A1(n332), .A2(n185), .A3(n391), .ZN(n31) );
  AND2_X1 U82 ( .A1(n336), .A2(n47), .ZN(n32) );
  AND3_X1 U83 ( .A1(n107), .A2(n108), .A3(n407), .ZN(n33) );
  NAND3_X1 U84 ( .A1(n125), .A2(n18), .A3(n191), .ZN(n416) );
  INV_X1 U86 ( .A(instr_rdata_i[2]), .ZN(n34) );
  OAI22_X2 U87 ( .A1(n79), .A2(n411), .B1(n63), .B2(n328), .ZN(
        imm_b_mux_sel_o[3]) );
  NAND2_X1 U88 ( .A1(n55), .A2(n191), .ZN(n485) );
  NAND2_X1 U89 ( .A1(n109), .A2(n33), .ZN(n579) );
  NAND2_X1 U90 ( .A1(n245), .A2(n39), .ZN(n583) );
  INV_X1 U91 ( .A(n230), .ZN(n46) );
  OAI21_X1 U92 ( .B1(n45), .B2(n44), .A(n41), .ZN(n43) );
  NAND2_X1 U93 ( .A1(n336), .A2(instr_rdata_i[25]), .ZN(n187) );
  NAND2_X1 U94 ( .A1(n441), .A2(n342), .ZN(n390) );
  INV_X1 U95 ( .A(instr_rdata_i[5]), .ZN(n49) );
  OAI21_X1 U96 ( .B1(n250), .B2(n487), .A(n249), .ZN(hwloop_we_o[0]) );
  INV_X1 U97 ( .A(instr_rdata_i[6]), .ZN(n127) );
  OAI21_X1 U98 ( .B1(n250), .B2(n446), .A(n249), .ZN(hwloop_we_o[1]) );
  OR2_X1 U99 ( .A1(n575), .A2(instr_rdata_i[3]), .ZN(n50) );
  NOR2_X1 U101 ( .A1(instr_rdata_i[2]), .A2(instr_rdata_i[6]), .ZN(n93) );
  INV_X1 U102 ( .A(instr_rdata_i[31]), .ZN(n414) );
  NAND2_X2 U103 ( .A1(instr_rdata_i[0]), .A2(instr_rdata_i[1]), .ZN(n575) );
  NAND3_X1 U104 ( .A1(n125), .A2(n51), .A3(instr_rdata_i[3]), .ZN(n193) );
  NAND2_X1 U105 ( .A1(n198), .A2(n288), .ZN(n415) );
  INV_X1 U106 ( .A(instr_rdata_i[4]), .ZN(n151) );
  NOR2_X1 U107 ( .A1(n151), .A2(n325), .ZN(n54) );
  NAND3_X1 U108 ( .A1(n125), .A2(n54), .A3(instr_rdata_i[3]), .ZN(n539) );
  OR2_X1 U109 ( .A1(n539), .A2(n575), .ZN(n560) );
  NOR2_X1 U110 ( .A1(n560), .A2(instr_rdata_i[13]), .ZN(\mult_imm_mux_o[0] )
         );
  INV_X1 U111 ( .A(\mult_imm_mux_o[0] ), .ZN(n282) );
  AND2_X1 U112 ( .A1(n51), .A2(n233), .ZN(n88) );
  NOR2_X1 U113 ( .A1(n551), .A2(instr_rdata_i[29]), .ZN(n314) );
  NAND2_X1 U114 ( .A1(n198), .A2(n558), .ZN(n446) );
  INV_X1 U115 ( .A(n446), .ZN(n420) );
  OR2_X1 U116 ( .A1(instr_rdata_i[30]), .A2(instr_rdata_i[28]), .ZN(n345) );
  NOR2_X1 U117 ( .A1(n345), .A2(n76), .ZN(n177) );
  NAND2_X1 U118 ( .A1(n177), .A2(instr_rdata_i[25]), .ZN(n346) );
  INV_X1 U119 ( .A(n346), .ZN(n400) );
  NAND3_X1 U120 ( .A1(n516), .A2(n420), .A3(n400), .ZN(n52) );
  OAI21_X1 U121 ( .B1(n282), .B2(n414), .A(n52), .ZN(mult_signed_mode_o[1]) );
  INV_X1 U122 ( .A(deassert_we_i), .ZN(n275) );
  INV_X1 U123 ( .A(n225), .ZN(n53) );
  NAND2_X1 U124 ( .A1(n275), .A2(n53), .ZN(n250) );
  NAND2_X1 U125 ( .A1(hwloop_start_mux_sel_o), .A2(n275), .ZN(n249) );
  NAND2_X1 U126 ( .A1(n54), .A2(n19), .ZN(n89) );
  INV_X1 U127 ( .A(n55), .ZN(n56) );
  NOR2_X1 U128 ( .A1(data_misaligned_i), .A2(n572), .ZN(n317) );
  INV_X1 U129 ( .A(n317), .ZN(n79) );
  INV_X1 U130 ( .A(instr_rdata_i[27]), .ZN(n349) );
  NOR2_X1 U131 ( .A1(n349), .A2(instr_rdata_i[26]), .ZN(n464) );
  NAND2_X1 U132 ( .A1(n464), .A2(instr_rdata_i[29]), .ZN(n59) );
  AND2_X1 U133 ( .A1(instr_rdata_i[28]), .A2(instr_rdata_i[29]), .ZN(n407) );
  INV_X1 U134 ( .A(instr_rdata_i[26]), .ZN(n541) );
  NAND2_X1 U135 ( .A1(n407), .A2(n541), .ZN(n58) );
  NAND2_X1 U137 ( .A1(n408), .A2(n360), .ZN(n57) );
  NAND3_X1 U138 ( .A1(n59), .A2(n58), .A3(n57), .ZN(n60) );
  NAND2_X1 U139 ( .A1(instr_rdata_i[31]), .A2(instr_rdata_i[30]), .ZN(n353) );
  INV_X1 U140 ( .A(n353), .ZN(n78) );
  NAND2_X1 U141 ( .A1(n60), .A2(n78), .ZN(n411) );
  AND2_X1 U143 ( .A1(n390), .A2(n446), .ZN(n62) );
  NOR2_X1 U144 ( .A1(n541), .A2(instr_rdata_i[27]), .ZN(n463) );
  INV_X1 U145 ( .A(instr_rdata_i[28]), .ZN(n218) );
  OR2_X1 U146 ( .A1(n218), .A2(instr_rdata_i[30]), .ZN(n67) );
  INV_X1 U147 ( .A(n67), .ZN(n61) );
  NAND2_X1 U148 ( .A1(n463), .A2(n61), .ZN(n341) );
  OR2_X1 U149 ( .A1(n341), .A2(instr_rdata_i[25]), .ZN(n181) );
  NOR2_X1 U150 ( .A1(n62), .A2(n181), .ZN(n301) );
  INV_X1 U151 ( .A(n416), .ZN(n379) );
  AOI22_X1 U152 ( .A1(n314), .A2(n301), .B1(n379), .B2(n17), .ZN(n63) );
  AND2_X1 U153 ( .A1(instr_rdata_i[12]), .A2(instr_rdata_i[13]), .ZN(n273) );
  OR2_X1 U154 ( .A1(n273), .A2(n288), .ZN(n85) );
  OR2_X1 U155 ( .A1(n355), .A2(n85), .ZN(n64) );
  NOR2_X1 U156 ( .A1(n328), .A2(n64), .ZN(n309) );
  INV_X1 U158 ( .A(n214), .ZN(n138) );
  NOR2_X1 U159 ( .A1(n546), .A2(n138), .ZN(n65) );
  AND2_X1 U160 ( .A1(n309), .A2(n65), .ZN(alu_op_b_mux_sel_o[2]) );
  INV_X1 U161 ( .A(n360), .ZN(n581) );
  INV_X1 U162 ( .A(instr_rdata_i[30]), .ZN(n547) );
  OR2_X1 U163 ( .A1(n547), .A2(instr_rdata_i[31]), .ZN(n210) );
  NOR2_X1 U164 ( .A1(n581), .A2(n210), .ZN(n525) );
  NAND2_X1 U165 ( .A1(n464), .A2(instr_rdata_i[28]), .ZN(n66) );
  NOR2_X1 U166 ( .A1(n66), .A2(n210), .ZN(n404) );
  INV_X1 U167 ( .A(instr_rdata_i[29]), .ZN(n468) );
  NOR2_X1 U168 ( .A1(n210), .A2(n468), .ZN(n173) );
  NAND2_X1 U169 ( .A1(n173), .A2(n218), .ZN(n207) );
  NOR2_X1 U170 ( .A1(n67), .A2(n76), .ZN(n392) );
  NAND3_X1 U171 ( .A1(n392), .A2(instr_rdata_i[31]), .A3(n468), .ZN(n503) );
  OAI21_X1 U172 ( .B1(n207), .B2(n76), .A(n503), .ZN(n476) );
  OR2_X1 U173 ( .A1(n218), .A2(instr_rdata_i[29]), .ZN(n113) );
  NOR2_X1 U174 ( .A1(n210), .A2(n113), .ZN(n467) );
  AND2_X1 U175 ( .A1(n467), .A2(n408), .ZN(n526) );
  OR2_X1 U176 ( .A1(n476), .A2(n526), .ZN(n377) );
  AOI211_X1 U177 ( .C1(n525), .C2(n541), .A(n404), .B(n377), .ZN(n513) );
  INV_X1 U178 ( .A(n207), .ZN(n364) );
  INV_X1 U179 ( .A(n407), .ZN(n100) );
  NOR2_X1 U180 ( .A1(n100), .A2(n210), .ZN(n462) );
  AOI22_X1 U181 ( .A1(n364), .A2(n464), .B1(n462), .B2(n408), .ZN(n498) );
  NOR2_X1 U182 ( .A1(instr_rdata_i[31]), .A2(instr_rdata_i[30]), .ZN(n501) );
  NAND3_X1 U183 ( .A1(n360), .A2(n501), .A3(instr_rdata_i[26]), .ZN(n70) );
  NAND2_X1 U184 ( .A1(n414), .A2(instr_rdata_i[29]), .ZN(n68) );
  NOR2_X1 U185 ( .A1(n68), .A2(n345), .ZN(n524) );
  AND2_X1 U186 ( .A1(instr_rdata_i[27]), .A2(instr_rdata_i[26]), .ZN(n469) );
  NAND2_X1 U187 ( .A1(n524), .A2(n469), .ZN(n69) );
  NAND4_X1 U188 ( .A1(n513), .A2(n498), .A3(n70), .A4(n69), .ZN(n435) );
  AND2_X1 U189 ( .A1(n177), .A2(instr_rdata_i[31]), .ZN(n299) );
  INV_X1 U190 ( .A(n501), .ZN(n470) );
  NOR2_X1 U191 ( .A1(n470), .A2(n349), .ZN(n405) );
  AOI22_X1 U192 ( .A1(n299), .A2(n468), .B1(n405), .B2(n407), .ZN(n371) );
  NAND2_X1 U193 ( .A1(n525), .A2(instr_rdata_i[26]), .ZN(n72) );
  NOR2_X1 U194 ( .A1(n113), .A2(n470), .ZN(n542) );
  OAI21_X1 U195 ( .B1(n542), .B2(n524), .A(n464), .ZN(n71) );
  NAND3_X1 U196 ( .A1(n463), .A2(n407), .A3(n501), .ZN(n362) );
  NAND4_X1 U197 ( .A1(n371), .A2(n72), .A3(n71), .A4(n362), .ZN(n300) );
  NAND2_X1 U198 ( .A1(n214), .A2(n464), .ZN(n277) );
  NAND3_X1 U199 ( .A1(n407), .A2(n469), .A3(instr_rdata_i[30]), .ZN(n74) );
  NAND2_X1 U200 ( .A1(instr_rdata_i[31]), .A2(instr_rdata_i[26]), .ZN(n73) );
  AND2_X1 U201 ( .A1(n74), .A2(n73), .ZN(n529) );
  OAI21_X1 U202 ( .B1(n277), .B2(instr_rdata_i[29]), .A(n529), .ZN(n375) );
  INV_X1 U203 ( .A(n277), .ZN(n278) );
  OAI21_X1 U204 ( .B1(n278), .B2(n299), .A(instr_rdata_i[29]), .ZN(n374) );
  NAND2_X1 U205 ( .A1(n176), .A2(n374), .ZN(n83) );
  NAND2_X1 U206 ( .A1(instr_rdata_i[31]), .A2(instr_rdata_i[29]), .ZN(n77) );
  INV_X1 U207 ( .A(n77), .ZN(n75) );
  AND2_X1 U208 ( .A1(n392), .A2(n75), .ZN(n554) );
  NOR2_X1 U209 ( .A1(n83), .A2(n554), .ZN(n208) );
  NOR2_X1 U210 ( .A1(n76), .A2(instr_rdata_i[28]), .ZN(n179) );
  NAND2_X1 U211 ( .A1(n179), .A2(instr_rdata_i[30]), .ZN(n347) );
  OR2_X1 U212 ( .A1(n347), .A2(n77), .ZN(n553) );
  INV_X1 U213 ( .A(n113), .ZN(n406) );
  NAND3_X1 U214 ( .A1(n406), .A2(n408), .A3(n78), .ZN(n172) );
  NAND2_X1 U215 ( .A1(n464), .A2(n78), .ZN(n80) );
  OR2_X1 U216 ( .A1(n80), .A2(n113), .ZN(n359) );
  AND3_X1 U217 ( .A1(n553), .A2(n172), .A3(n359), .ZN(n82) );
  AND2_X1 U218 ( .A1(n467), .A2(n469), .ZN(n500) );
  INV_X1 U219 ( .A(n80), .ZN(n81) );
  NAND2_X1 U220 ( .A1(n81), .A2(n360), .ZN(n372) );
  NAND3_X1 U221 ( .A1(n82), .A2(n411), .A3(n372), .ZN(n461) );
  NOR3_X1 U222 ( .A1(n83), .A2(n500), .A3(n461), .ZN(n84) );
  INV_X1 U223 ( .A(n481), .ZN(n436) );
  NOR3_X1 U224 ( .A1(n84), .A2(n533), .A3(n436), .ZN(n91) );
  AOI21_X1 U225 ( .B1(n301), .B2(n468), .A(instr_rdata_i[31]), .ZN(n87) );
  INV_X1 U226 ( .A(n546), .ZN(n268) );
  AOI21_X1 U227 ( .B1(n268), .B2(n85), .A(n138), .ZN(n86) );
  NOR3_X1 U228 ( .A1(n87), .A2(n86), .A3(n355), .ZN(n90) );
  OR2_X1 U229 ( .A1(n485), .A2(n233), .ZN(n320) );
  NAND3_X1 U230 ( .A1(n127), .A2(n233), .A3(n594), .ZN(n134) );
  OR2_X1 U231 ( .A1(n134), .A2(n151), .ZN(n484) );
  NAND2_X1 U232 ( .A1(n320), .A2(n484), .ZN(n306) );
  NAND2_X1 U233 ( .A1(n88), .A2(n125), .ZN(n381) );
  INV_X1 U234 ( .A(n487), .ZN(n245) );
  OAI21_X1 U235 ( .B1(n381), .B2(n245), .A(n488), .ZN(n235) );
  NOR4_X1 U236 ( .A1(n91), .A2(n90), .A3(n306), .A4(n235), .ZN(n98) );
  OR2_X1 U237 ( .A1(instr_rdata_i[6]), .A2(instr_rdata_i[4]), .ZN(n92) );
  NOR2_X1 U238 ( .A1(n92), .A2(n594), .ZN(n292) );
  AND2_X1 U239 ( .A1(n292), .A2(n507), .ZN(n265) );
  NAND2_X1 U240 ( .A1(n265), .A2(n322), .ZN(n274) );
  INV_X1 U241 ( .A(n274), .ZN(n96) );
  NAND2_X1 U242 ( .A1(n481), .A2(instr_rdata_i[12]), .ZN(n331) );
  NAND2_X1 U243 ( .A1(instr_rdata_i[13]), .A2(n595), .ZN(n199) );
  NOR2_X1 U244 ( .A1(n560), .A2(n199), .ZN(n563) );
  NAND2_X1 U245 ( .A1(n30), .A2(n93), .ZN(n197) );
  INV_X1 U246 ( .A(n38), .ZN(n95) );
  INV_X1 U247 ( .A(n596), .ZN(n94) );
  AOI211_X1 U248 ( .C1(n17), .C2(n95), .A(n94), .B(data_misaligned_i), .ZN(
        n308) );
  OAI21_X1 U249 ( .B1(n288), .B2(n559), .A(n308), .ZN(n298) );
  AOI211_X1 U250 ( .C1(n96), .C2(n331), .A(n563), .B(n298), .ZN(n97) );
  OAI21_X1 U251 ( .B1(n98), .B2(n575), .A(n97), .ZN(alu_op_b_mux_sel_o[1]) );
  INV_X1 U252 ( .A(n563), .ZN(n99) );
  OAI21_X1 U253 ( .B1(current_priv_lvl_i[1]), .B2(n218), .A(n100), .ZN(n102)
         );
  INV_X1 U254 ( .A(current_priv_lvl_i[0]), .ZN(n101) );
  NAND2_X1 U255 ( .A1(n102), .A2(n101), .ZN(n103) );
  INV_X1 U256 ( .A(n289), .ZN(n271) );
  OAI211_X1 U257 ( .C1(current_priv_lvl_i[1]), .C2(n468), .A(n103), .B(n271), 
        .ZN(n262) );
  OR2_X1 U258 ( .A1(instr_rdata_i[27]), .A2(instr_rdata_i[30]), .ZN(n104) );
  NOR2_X1 U259 ( .A1(n104), .A2(instr_rdata_i[25]), .ZN(n141) );
  INV_X1 U260 ( .A(instr_rdata_i[20]), .ZN(n111) );
  INV_X1 U261 ( .A(instr_rdata_i[24]), .ZN(n105) );
  INV_X1 U262 ( .A(instr_rdata_i[22]), .ZN(n107) );
  NAND4_X1 U263 ( .A1(n141), .A2(n111), .A3(n105), .A4(n107), .ZN(n110) );
  INV_X1 U264 ( .A(instr_rdata_i[21]), .ZN(n106) );
  NOR2_X1 U265 ( .A1(n110), .A2(n106), .ZN(n580) );
  NAND2_X1 U266 ( .A1(n580), .A2(n407), .ZN(n584) );
  NAND2_X1 U267 ( .A1(instr_rdata_i[25]), .A2(instr_rdata_i[24]), .ZN(n251) );
  NOR3_X1 U268 ( .A1(n251), .A2(n106), .A3(instr_rdata_i[20]), .ZN(n109) );
  NOR2_X1 U269 ( .A1(n547), .A2(n349), .ZN(n108) );
  NAND2_X1 U270 ( .A1(current_priv_lvl_i[0]), .A2(current_priv_lvl_i[1]), .ZN(
        n586) );
  INV_X1 U271 ( .A(n110), .ZN(n256) );
  NAND2_X1 U272 ( .A1(n256), .A2(n360), .ZN(n247) );
  NOR4_X1 U273 ( .A1(n111), .A2(instr_rdata_i[24]), .A3(instr_rdata_i[22]), 
        .A4(instr_rdata_i[21]), .ZN(n112) );
  NAND3_X1 U274 ( .A1(n141), .A2(n360), .A3(n112), .ZN(n252) );
  NOR3_X1 U275 ( .A1(n113), .A2(instr_rdata_i[24]), .A3(instr_rdata_i[21]), 
        .ZN(n114) );
  NAND4_X1 U276 ( .A1(n114), .A2(n141), .A3(instr_rdata_i[22]), .A4(
        instr_rdata_i[20]), .ZN(n578) );
  NAND3_X1 U277 ( .A1(n247), .A2(n252), .A3(n578), .ZN(n121) );
  OR2_X1 U278 ( .A1(instr_rdata_i[10]), .A2(instr_rdata_i[11]), .ZN(n115) );
  NOR3_X1 U279 ( .A1(n115), .A2(instr_rdata_i[7]), .A3(instr_rdata_i[8]), .ZN(
        n119) );
  OR2_X1 U280 ( .A1(instr_rdata_i[9]), .A2(instr_rdata_i[17]), .ZN(n116) );
  NOR3_X1 U281 ( .A1(n116), .A2(instr_rdata_i[18]), .A3(instr_rdata_i[19]), 
        .ZN(n118) );
  NOR3_X1 U282 ( .A1(instr_rdata_i[23]), .A2(instr_rdata_i[15]), .A3(
        instr_rdata_i[16]), .ZN(n117) );
  NOR2_X1 U283 ( .A1(instr_rdata_i[26]), .A2(instr_rdata_i[31]), .ZN(n255) );
  NAND4_X1 U284 ( .A1(n119), .A2(n118), .A3(n117), .A4(n255), .ZN(n246) );
  INV_X1 U285 ( .A(n246), .ZN(n120) );
  OAI21_X1 U286 ( .B1(n122), .B2(n121), .A(n120), .ZN(n123) );
  INV_X1 U287 ( .A(n381), .ZN(n326) );
  INV_X1 U288 ( .A(n30), .ZN(n135) );
  MUX2_X1 U289 ( .A(n151), .B(n135), .S(n125), .Z(n133) );
  MUX2_X1 U290 ( .A(instr_rdata_i[3]), .B(instr_rdata_i[4]), .S(n593), .Z(n124) );
  NAND2_X1 U291 ( .A1(n124), .A2(n594), .ZN(n131) );
  NAND2_X1 U292 ( .A1(n125), .A2(n19), .ZN(n126) );
  NAND2_X1 U293 ( .A1(n126), .A2(instr_rdata_i[4]), .ZN(n129) );
  NAND2_X1 U294 ( .A1(n134), .A2(n127), .ZN(n128) );
  NAND2_X1 U295 ( .A1(n129), .A2(n128), .ZN(n130) );
  MUX2_X1 U296 ( .A(n131), .B(n130), .S(n322), .Z(n132) );
  OAI21_X1 U297 ( .B1(n133), .B2(n18), .A(n132), .ZN(n243) );
  OAI21_X1 U298 ( .B1(n135), .B2(n134), .A(n507), .ZN(n136) );
  NOR2_X1 U299 ( .A1(n243), .A2(n136), .ZN(n195) );
  AND2_X1 U300 ( .A1(n546), .A2(n214), .ZN(n237) );
  NOR2_X1 U301 ( .A1(n436), .A2(n353), .ZN(n137) );
  OR2_X1 U302 ( .A1(n237), .A2(n137), .ZN(n189) );
  OR2_X1 U303 ( .A1(n289), .A2(n558), .ZN(n515) );
  NOR2_X1 U304 ( .A1(n138), .A2(n515), .ZN(n139) );
  INV_X1 U305 ( .A(n355), .ZN(n548) );
  OAI21_X1 U306 ( .B1(n189), .B2(n139), .A(n548), .ZN(n140) );
  NAND2_X1 U307 ( .A1(n195), .A2(n140), .ZN(n384) );
  INV_X1 U308 ( .A(n384), .ZN(n169) );
  OAI21_X1 U309 ( .B1(n289), .B2(n273), .A(instr_rdata_i[26]), .ZN(n142) );
  NAND2_X1 U310 ( .A1(n142), .A2(n141), .ZN(n144) );
  NOR2_X1 U311 ( .A1(n446), .A2(n541), .ZN(n143) );
  MUX2_X1 U313 ( .A(n356), .B(n288), .S(instr_rdata_i[25]), .Z(n146) );
  OR2_X1 U314 ( .A1(n558), .A2(instr_rdata_i[12]), .ZN(n480) );
  NAND3_X1 U315 ( .A1(n480), .A2(n408), .A3(n545), .ZN(n145) );
  OAI21_X1 U316 ( .B1(n146), .B2(n145), .A(n595), .ZN(n148) );
  INV_X1 U317 ( .A(instr_rdata_i[25]), .ZN(n184) );
  INV_X1 U318 ( .A(n469), .ZN(n433) );
  OAI211_X1 U319 ( .C1(n408), .C2(n184), .A(n433), .B(n468), .ZN(n147) );
  NOR2_X1 U320 ( .A1(n336), .A2(n551), .ZN(n167) );
  NOR2_X1 U321 ( .A1(n546), .A2(n470), .ZN(n254) );
  NOR2_X1 U322 ( .A1(n546), .A2(n210), .ZN(n354) );
  OR2_X1 U323 ( .A1(n254), .A2(n354), .ZN(n455) );
  INV_X1 U324 ( .A(n488), .ZN(n418) );
  INV_X1 U325 ( .A(n415), .ZN(n454) );
  NAND2_X1 U326 ( .A1(n418), .A2(n454), .ZN(n150) );
  NOR2_X1 U327 ( .A1(n455), .A2(n150), .ZN(n424) );
  INV_X1 U328 ( .A(n533), .ZN(n535) );
  INV_X1 U329 ( .A(n529), .ZN(n154) );
  NOR2_X1 U330 ( .A1(n593), .A2(n325), .ZN(n152) );
  NAND4_X1 U331 ( .A1(n152), .A2(instr_rdata_i[3]), .A3(n594), .A4(n151), .ZN(
        n576) );
  NOR2_X1 U332 ( .A1(n576), .A2(n574), .ZN(n153) );
  AOI211_X1 U333 ( .C1(n535), .C2(n154), .A(illegal_c_insn_i), .B(n153), .ZN(
        n165) );
  NOR2_X1 U334 ( .A1(n485), .A2(instr_rdata_i[3]), .ZN(n156) );
  INV_X1 U335 ( .A(n193), .ZN(n155) );
  AOI22_X1 U336 ( .A1(n156), .A2(n487), .B1(n155), .B2(n481), .ZN(n164) );
  AND2_X1 U337 ( .A1(n292), .A2(n322), .ZN(n196) );
  NAND2_X1 U338 ( .A1(n345), .A2(instr_rdata_i[29]), .ZN(n158) );
  NAND4_X1 U339 ( .A1(n333), .A2(n288), .A3(n414), .A4(n158), .ZN(n159) );
  NAND2_X1 U340 ( .A1(n196), .A2(n159), .ZN(n160) );
  NAND2_X1 U341 ( .A1(n160), .A2(n197), .ZN(n161) );
  NAND2_X1 U342 ( .A1(n161), .A2(n273), .ZN(n163) );
  NOR3_X1 U345 ( .A1(n167), .A2(n424), .A3(n166), .ZN(n168) );
  OR2_X1 U347 ( .A1(n355), .A2(n575), .ZN(n227) );
  NOR3_X1 U348 ( .A1(n227), .A2(n353), .A3(n592), .ZN(alu_operator_o[6]) );
  NAND2_X1 U349 ( .A1(n574), .A2(instr_rdata_i[25]), .ZN(n171) );
  OR2_X1 U350 ( .A1(n347), .A2(n171), .ZN(n566) );
  OAI21_X1 U351 ( .B1(n346), .B2(n288), .A(n566), .ZN(n338) );
  NOR2_X1 U352 ( .A1(n551), .A2(n575), .ZN(n219) );
  NAND2_X1 U353 ( .A1(n32), .A2(n219), .ZN(regc_mux_o[0]) );
  INV_X1 U354 ( .A(n411), .ZN(n174) );
  INV_X1 U355 ( .A(n172), .ZN(n363) );
  NOR4_X1 U356 ( .A1(n174), .A2(n500), .A3(n363), .A4(n173), .ZN(n175) );
  AOI21_X1 U357 ( .B1(n176), .B2(n175), .A(n533), .ZN(n206) );
  NAND2_X1 U358 ( .A1(n400), .A2(n288), .ZN(n565) );
  INV_X1 U359 ( .A(n565), .ZN(n209) );
  NAND2_X1 U360 ( .A1(n177), .A2(n184), .ZN(n477) );
  NOR2_X1 U361 ( .A1(n477), .A2(n331), .ZN(n350) );
  INV_X1 U362 ( .A(n345), .ZN(n182) );
  NAND2_X1 U363 ( .A1(n182), .A2(n184), .ZN(n440) );
  INV_X1 U364 ( .A(n463), .ZN(n178) );
  NOR3_X1 U365 ( .A1(n440), .A2(n178), .A3(n558), .ZN(n180) );
  OR2_X1 U366 ( .A1(n487), .A2(instr_rdata_i[25]), .ZN(n393) );
  INV_X1 U367 ( .A(n179), .ZN(n450) );
  NOR2_X1 U368 ( .A1(n393), .A2(n450), .ZN(n479) );
  NOR4_X1 U369 ( .A1(n209), .A2(n350), .A3(n180), .A4(n479), .ZN(n186) );
  NAND2_X1 U370 ( .A1(n481), .A2(n342), .ZN(n389) );
  NOR2_X1 U371 ( .A1(n181), .A2(n389), .ZN(n332) );
  NAND2_X1 U372 ( .A1(n463), .A2(n182), .ZN(n183) );
  NOR2_X1 U373 ( .A1(n393), .A2(n183), .ZN(n185) );
  AND2_X1 U374 ( .A1(n392), .A2(n184), .ZN(n391) );
  OR2_X1 U375 ( .A1(n415), .A2(instr_rdata_i[25]), .ZN(n451) );
  NOR2_X1 U376 ( .A1(n451), .A2(n341), .ZN(n220) );
  NOR2_X1 U377 ( .A1(n301), .A2(n220), .ZN(n445) );
  NAND3_X1 U378 ( .A1(n186), .A2(n31), .A3(n445), .ZN(n497) );
  NOR2_X1 U379 ( .A1(n497), .A2(n187), .ZN(n291) );
  AOI21_X1 U380 ( .B1(n291), .B2(n346), .A(n551), .ZN(n205) );
  INV_X1 U381 ( .A(n356), .ZN(n188) );
  AOI21_X1 U382 ( .B1(n188), .B2(n271), .A(n353), .ZN(n190) );
  AOI211_X1 U383 ( .C1(n214), .C2(n390), .A(n190), .B(n189), .ZN(n203) );
  INV_X1 U384 ( .A(n306), .ZN(n194) );
  NAND3_X1 U385 ( .A1(n30), .A2(n593), .A3(n18), .ZN(n192) );
  AND2_X1 U386 ( .A1(n193), .A2(n576), .ZN(n382) );
  NAND4_X1 U387 ( .A1(n195), .A2(n194), .A3(n229), .A4(n382), .ZN(n293) );
  NOR2_X1 U388 ( .A1(n293), .A2(n196), .ZN(n202) );
  INV_X1 U389 ( .A(n197), .ZN(n316) );
  INV_X1 U390 ( .A(n199), .ZN(n540) );
  NOR3_X1 U391 ( .A1(n539), .A2(n198), .A3(n540), .ZN(n200) );
  AOI211_X1 U392 ( .C1(n316), .C2(n558), .A(n326), .B(n200), .ZN(n201) );
  OAI211_X1 U393 ( .C1(n203), .C2(n355), .A(n202), .B(n201), .ZN(n204) );
  OR3_X1 U394 ( .A1(n206), .A2(n205), .A3(n204), .ZN(regc_mux_o[1]) );
  NOR3_X1 U395 ( .A1(n572), .A2(n207), .A3(n433), .ZN(is_subrot_o) );
  OR3_X1 U396 ( .A1(n208), .A2(n481), .A3(n572), .ZN(n223) );
  INV_X1 U397 ( .A(n572), .ZN(n543) );
  AOI22_X1 U398 ( .A1(n516), .A2(n209), .B1(n461), .B2(n543), .ZN(n522) );
  OAI211_X1 U399 ( .C1(n38), .C2(n17), .A(n559), .B(n560), .ZN(n217) );
  INV_X1 U400 ( .A(is_subrot_o), .ZN(n213) );
  INV_X1 U401 ( .A(n210), .ZN(n211) );
  NAND4_X1 U402 ( .A1(n543), .A2(n463), .A3(n211), .A4(n581), .ZN(n212) );
  NAND2_X1 U403 ( .A1(n213), .A2(n212), .ZN(n296) );
  NOR2_X1 U404 ( .A1(n274), .A2(n331), .ZN(n269) );
  NAND2_X1 U405 ( .A1(n515), .A2(n214), .ZN(n215) );
  OR2_X1 U406 ( .A1(n546), .A2(n215), .ZN(n537) );
  NOR2_X1 U407 ( .A1(n227), .A2(n537), .ZN(n248) );
  OR3_X1 U408 ( .A1(n296), .A2(n269), .A3(n248), .ZN(n216) );
  AOI211_X1 U409 ( .C1(n219), .C2(n218), .A(n217), .B(n216), .ZN(n222) );
  OAI21_X1 U410 ( .B1(n332), .B2(n220), .A(n516), .ZN(n221) );
  NAND4_X1 U411 ( .A1(n223), .A2(n522), .A3(n222), .A4(n221), .ZN(regb_used_o)
         );
  NAND2_X1 U412 ( .A1(n487), .A2(n507), .ZN(n224) );
  NOR2_X1 U413 ( .A1(n381), .A2(n224), .ZN(csr_access_o) );
  NAND2_X1 U414 ( .A1(n289), .A2(n288), .ZN(n378) );
  OAI21_X1 U415 ( .B1(n546), .B2(n414), .A(n353), .ZN(n226) );
  INV_X1 U416 ( .A(n226), .ZN(n228) );
  INV_X1 U417 ( .A(n292), .ZN(n483) );
  AOI21_X1 U418 ( .B1(csr_access_o), .B2(n558), .A(hwloop_cnt_mux_sel_o), .ZN(
        n232) );
  INV_X1 U419 ( .A(n590), .ZN(n231) );
  NOR2_X1 U420 ( .A1(n485), .A2(n487), .ZN(n234) );
  MUX2_X1 U421 ( .A(n265), .B(n234), .S(n19), .Z(n236) );
  NOR2_X1 U422 ( .A1(n236), .A2(n235), .ZN(n240) );
  NOR2_X1 U423 ( .A1(n237), .A2(n355), .ZN(n238) );
  NOR3_X1 U424 ( .A1(n238), .A2(n306), .A3(n242), .ZN(n239) );
  AOI21_X1 U425 ( .B1(n240), .B2(n239), .A(n328), .ZN(regfile_alu_we_dec_o) );
  NAND4_X1 U426 ( .A1(n382), .A2(instr_rdata_i[3]), .A3(n507), .A4(n485), .ZN(
        n241) );
  OR3_X1 U427 ( .A1(n243), .A2(n242), .A3(n241), .ZN(regfile_alu_waddr_sel_o)
         );
  INV_X1 U428 ( .A(data_misaligned_i), .ZN(n310) );
  AND2_X1 U429 ( .A1(n310), .A2(mult_multicycle_i), .ZN(n244) );
  NOR2_X1 U430 ( .A1(n244), .A2(n559), .ZN(alu_op_c_mux_sel_o[0]) );
  NOR2_X1 U431 ( .A1(n244), .A2(n38), .ZN(alu_op_c_mux_sel_o[1]) );
  NOR2_X1 U432 ( .A1(n583), .A2(n252), .ZN(ebrk_insn_o) );
  OAI21_X1 U433 ( .B1(n596), .B2(n487), .A(n38), .ZN(jump_in_dec_o[1]) );
  OR2_X1 U434 ( .A1(n320), .A2(n575), .ZN(n304) );
  NAND2_X1 U435 ( .A1(n304), .A2(n38), .ZN(jump_in_dec_o[0]) );
  NOR3_X1 U436 ( .A1(n583), .A2(instr_rdata_i[21]), .A3(n247), .ZN(
        ecall_insn_o) );
  NAND2_X1 U437 ( .A1(n516), .A2(n391), .ZN(n518) );
  NOR2_X1 U438 ( .A1(n518), .A2(n558), .ZN(n493) );
  OR2_X1 U439 ( .A1(n493), .A2(n543), .ZN(alu_vec_mode_o[1]) );
  INV_X1 U440 ( .A(n248), .ZN(alu_bmask_a_mux_sel_o) );
  INV_X1 U441 ( .A(csr_access_o), .ZN(imm_a_mux_sel_o[0]) );
  INV_X1 U442 ( .A(n464), .ZN(n472) );
  NOR3_X1 U443 ( .A1(n472), .A2(instr_rdata_i[22]), .A3(n251), .ZN(n261) );
  NOR3_X1 U444 ( .A1(n252), .A2(instr_rdata_i[31]), .A3(n541), .ZN(n260) );
  NOR3_X1 U445 ( .A1(instr_rdata_i[22]), .A2(instr_rdata_i[24]), .A3(
        instr_rdata_i[20]), .ZN(n253) );
  NAND2_X1 U446 ( .A1(n254), .A2(n253), .ZN(n258) );
  NAND3_X1 U447 ( .A1(n256), .A2(n407), .A3(n255), .ZN(n257) );
  AOI21_X1 U448 ( .B1(n258), .B2(n257), .A(instr_rdata_i[21]), .ZN(n259) );
  AOI211_X1 U449 ( .C1(n462), .C2(n261), .A(n260), .B(n259), .ZN(n263) );
  NOR4_X1 U450 ( .A1(n263), .A2(instr_rdata_i[23]), .A3(n262), .A4(
        imm_a_mux_sel_o[0]), .ZN(csr_status_o) );
  AND2_X1 U451 ( .A1(n275), .A2(jump_in_dec_o[0]), .ZN(jump_in_id_o[0]) );
  AND2_X1 U452 ( .A1(jump_in_dec_o[1]), .A2(n275), .ZN(jump_in_id_o[1]) );
  NOR2_X1 U453 ( .A1(n274), .A2(n389), .ZN(data_load_event_o) );
  INV_X1 U454 ( .A(n269), .ZN(n264) );
  OAI22_X1 U455 ( .A1(n264), .A2(n595), .B1(n288), .B2(n274), .ZN(
        data_sign_extension_o[0]) );
  INV_X1 U456 ( .A(n265), .ZN(n272) );
  INV_X1 U457 ( .A(n198), .ZN(n561) );
  NAND4_X1 U458 ( .A1(n269), .A2(n406), .A3(n333), .A4(n414), .ZN(n267) );
  OAI21_X1 U459 ( .B1(n272), .B2(n561), .A(n267), .ZN(data_type_o[0]) );
  NAND3_X1 U460 ( .A1(n269), .A2(n268), .A3(n414), .ZN(n270) );
  OAI21_X1 U461 ( .B1(n272), .B2(n271), .A(n270), .ZN(data_type_o[1]) );
  OR2_X1 U462 ( .A1(data_misaligned_i), .A2(regfile_alu_waddr_sel_o), .ZN(
        prepost_useincr_o) );
  NOR2_X1 U463 ( .A1(n559), .A2(n273), .ZN(data_we_o) );
  NOR2_X1 U464 ( .A1(deassert_we_i), .A2(n274), .ZN(regfile_mem_we_o) );
  AOI21_X1 U465 ( .B1(data_we_o), .B2(n275), .A(regfile_mem_we_o), .ZN(n276)
         );
  INV_X1 U466 ( .A(n276), .ZN(data_req_o) );
  NOR3_X1 U467 ( .A1(deassert_we_i), .A2(n342), .A3(imm_a_mux_sel_o[0]), .ZN(
        csr_op_o[0]) );
  NOR3_X1 U468 ( .A1(deassert_we_i), .A2(n545), .A3(imm_a_mux_sel_o[0]), .ZN(
        csr_op_o[1]) );
  AND2_X1 U469 ( .A1(regfile_alu_we_dec_o), .A2(n275), .ZN(regfile_alu_we_o)
         );
  NAND2_X1 U470 ( .A1(n467), .A2(n463), .ZN(n373) );
  AOI21_X1 U471 ( .B1(n277), .B2(n373), .A(n572), .ZN(mult_dot_signed_o[0]) );
  NAND2_X1 U472 ( .A1(n278), .A2(instr_rdata_i[28]), .ZN(n279) );
  AOI21_X1 U473 ( .B1(n373), .B2(n279), .A(n572), .ZN(mult_dot_signed_o[1]) );
  INV_X1 U474 ( .A(mult_signed_mode_o[1]), .ZN(n281) );
  INV_X1 U475 ( .A(n390), .ZN(n569) );
  NAND3_X1 U476 ( .A1(n516), .A2(n400), .A3(n569), .ZN(n280) );
  NAND2_X1 U477 ( .A1(n281), .A2(n280), .ZN(mult_signed_mode_o[0]) );
  NOR2_X1 U478 ( .A1(n282), .A2(n547), .ZN(mult_sel_subword_o) );
  AOI21_X1 U479 ( .B1(n543), .B2(n299), .A(mult_dot_signed_o[0]), .ZN(n283) );
  NOR2_X1 U480 ( .A1(deassert_we_i), .A2(n283), .ZN(mult_dot_en_o) );
  AOI21_X1 U481 ( .B1(n516), .B2(n338), .A(\mult_imm_mux_o[0] ), .ZN(n284) );
  NOR2_X1 U482 ( .A1(deassert_we_i), .A2(n284), .ZN(mult_int_en_o) );
  INV_X1 U483 ( .A(n347), .ZN(n285) );
  NAND4_X1 U484 ( .A1(n516), .A2(n420), .A3(n285), .A4(instr_rdata_i[25]), 
        .ZN(n287) );
  AOI22_X1 U485 ( .A1(n543), .A2(n342), .B1(\mult_imm_mux_o[0] ), .B2(n157), 
        .ZN(n286) );
  NAND2_X1 U486 ( .A1(n287), .A2(n286), .ZN(mult_operator_o[0]) );
  OR2_X1 U487 ( .A1(n289), .A2(n288), .ZN(n290) );
  OR2_X1 U488 ( .A1(n346), .A2(n290), .ZN(n295) );
  AOI21_X1 U489 ( .B1(n291), .B2(n414), .A(n355), .ZN(n294) );
  OR3_X1 U490 ( .A1(n293), .A2(n292), .A3(n326), .ZN(n536) );
  NOR2_X1 U491 ( .A1(n294), .A2(n536), .ZN(n532) );
  OAI211_X1 U492 ( .C1(n355), .C2(n295), .A(n532), .B(n539), .ZN(
        mult_operator_o[1]) );
  INV_X1 U493 ( .A(n516), .ZN(n564) );
  OR2_X1 U494 ( .A1(n564), .A2(n295), .ZN(n570) );
  NAND2_X1 U495 ( .A1(n570), .A2(n572), .ZN(mult_operator_o[2]) );
  INV_X1 U496 ( .A(n500), .ZN(n431) );
  INV_X1 U497 ( .A(n296), .ZN(n297) );
  OAI21_X1 U498 ( .B1(n572), .B2(n431), .A(n297), .ZN(is_clpx_o) );
  INV_X1 U499 ( .A(n298), .ZN(n305) );
  OAI21_X1 U500 ( .B1(n300), .B2(n299), .A(n543), .ZN(n303) );
  NAND2_X1 U501 ( .A1(n516), .A2(n301), .ZN(n302) );
  NAND4_X1 U502 ( .A1(n305), .A2(n304), .A3(n303), .A4(n302), .ZN(
        imm_b_mux_sel_o[0]) );
  AOI22_X1 U503 ( .A1(n543), .A2(n411), .B1(n306), .B2(n507), .ZN(n307) );
  NAND2_X1 U504 ( .A1(n308), .A2(n307), .ZN(imm_b_mux_sel_o[1]) );
  INV_X1 U505 ( .A(n309), .ZN(n313) );
  INV_X1 U506 ( .A(alu_op_b_mux_sel_o[2]), .ZN(n312) );
  AOI22_X1 U507 ( .A1(n317), .A2(n411), .B1(n310), .B2(alu_operator_o[6]), 
        .ZN(n311) );
  OAI211_X1 U508 ( .C1(n313), .C2(n353), .A(n312), .B(n311), .ZN(
        imm_b_mux_sel_o[2]) );
  OAI22_X1 U509 ( .A1(n518), .A2(n436), .B1(n342), .B2(n572), .ZN(
        alu_vec_mode_o[0]) );
  INV_X1 U510 ( .A(n314), .ZN(n315) );
  NOR2_X1 U511 ( .A1(n315), .A2(n565), .ZN(n327) );
  AOI21_X1 U512 ( .B1(n316), .B2(n288), .A(n327), .ZN(n319) );
  AOI21_X1 U513 ( .B1(n554), .B2(n317), .A(alu_op_a_mux_sel_o[2]), .ZN(n318)
         );
  OAI21_X1 U514 ( .B1(n319), .B2(n328), .A(n318), .ZN(alu_op_b_mux_sel_o[0])
         );
  INV_X1 U515 ( .A(n484), .ZN(n324) );
  INV_X1 U516 ( .A(n320), .ZN(n321) );
  AOI211_X1 U517 ( .C1(n324), .C2(n322), .A(n321), .B(n327), .ZN(n323) );
  OAI22_X1 U518 ( .A1(n328), .A2(n323), .B1(data_misaligned_i), .B2(n596), 
        .ZN(alu_op_a_mux_sel_o[0]) );
  AOI22_X1 U519 ( .A1(n326), .A2(n157), .B1(n325), .B2(n324), .ZN(n330) );
  INV_X1 U520 ( .A(n327), .ZN(n329) );
  AOI21_X1 U521 ( .B1(n330), .B2(n329), .A(n328), .ZN(alu_op_a_mux_sel_o[1])
         );
  INV_X1 U522 ( .A(n331), .ZN(n399) );
  AOI22_X1 U523 ( .A1(n399), .A2(n463), .B1(instr_rdata_i[12]), .B2(n17), .ZN(
        n335) );
  AOI21_X1 U524 ( .B1(n333), .B2(n420), .A(n332), .ZN(n334) );
  OAI21_X1 U525 ( .B1(n335), .B2(n440), .A(n334), .ZN(n340) );
  INV_X1 U526 ( .A(n336), .ZN(n339) );
  OAI22_X1 U527 ( .A1(n346), .A2(n389), .B1(n477), .B2(n378), .ZN(n337) );
  NOR4_X1 U528 ( .A1(n340), .A2(n339), .A3(n338), .A4(n337), .ZN(n403) );
  INV_X1 U529 ( .A(n341), .ZN(n344) );
  OAI21_X1 U530 ( .B1(n342), .B2(n558), .A(n390), .ZN(n343) );
  AOI22_X1 U531 ( .A1(n344), .A2(n569), .B1(n343), .B2(n392), .ZN(n352) );
  NOR2_X1 U532 ( .A1(n451), .A2(n345), .ZN(n401) );
  OAI22_X1 U533 ( .A1(n347), .A2(n393), .B1(n346), .B2(n378), .ZN(n348) );
  AOI21_X1 U534 ( .B1(n401), .B2(n349), .A(n348), .ZN(n351) );
  INV_X1 U535 ( .A(n350), .ZN(n444) );
  AND4_X1 U536 ( .A1(n403), .A2(n352), .A3(n351), .A4(n444), .ZN(n388) );
  OR2_X1 U537 ( .A1(n355), .A2(n353), .ZN(n482) );
  OAI21_X1 U538 ( .B1(n354), .B2(n488), .A(n482), .ZN(n370) );
  OAI21_X1 U539 ( .B1(n355), .B2(n414), .A(n488), .ZN(n413) );
  OAI21_X1 U540 ( .B1(n413), .B2(n379), .A(n356), .ZN(n358) );
  INV_X1 U541 ( .A(n389), .ZN(n419) );
  INV_X1 U542 ( .A(n539), .ZN(n380) );
  AOI22_X1 U543 ( .A1(n379), .A2(n419), .B1(n380), .B2(instr_rdata_i[12]), 
        .ZN(n357) );
  NAND2_X1 U544 ( .A1(n418), .A2(n399), .ZN(n506) );
  NAND3_X1 U545 ( .A1(n358), .A2(n357), .A3(n506), .ZN(n369) );
  INV_X1 U546 ( .A(n359), .ZN(n555) );
  NAND2_X1 U547 ( .A1(n364), .A2(instr_rdata_i[26]), .ZN(n502) );
  INV_X1 U548 ( .A(n554), .ZN(n430) );
  NAND2_X1 U549 ( .A1(n405), .A2(n360), .ZN(n361) );
  NAND4_X1 U550 ( .A1(n502), .A2(n362), .A3(n430), .A4(n361), .ZN(n475) );
  AOI211_X1 U551 ( .C1(n363), .C2(instr_rdata_i[25]), .A(n555), .B(n475), .ZN(
        n367) );
  INV_X1 U552 ( .A(n525), .ZN(n432) );
  NOR2_X1 U553 ( .A1(n364), .A2(n524), .ZN(n365) );
  MUX2_X1 U554 ( .A(n432), .B(n365), .S(n464), .Z(n366) );
  AOI21_X1 U555 ( .B1(n367), .B2(n366), .A(n533), .ZN(n368) );
  AOI211_X1 U556 ( .C1(n454), .C2(n370), .A(n369), .B(n368), .ZN(n387) );
  INV_X1 U557 ( .A(n371), .ZN(n376) );
  NAND3_X1 U558 ( .A1(n374), .A2(n373), .A3(n372), .ZN(n557) );
  OR4_X1 U559 ( .A1(n377), .A2(n376), .A3(n557), .A4(n375), .ZN(n386) );
  INV_X1 U560 ( .A(n378), .ZN(n439) );
  AOI22_X1 U561 ( .A1(n418), .A2(n439), .B1(n379), .B2(n399), .ZN(n383) );
  NAND2_X1 U562 ( .A1(n380), .A2(n545), .ZN(n549) );
  NAND4_X1 U563 ( .A1(n383), .A2(n382), .A3(n381), .A4(n549), .ZN(n385) );
  AOI211_X1 U564 ( .C1(n535), .C2(n386), .A(n385), .B(n384), .ZN(n428) );
  OAI211_X1 U565 ( .C1(n388), .C2(n551), .A(n387), .B(n428), .ZN(
        alu_operator_o[0]) );
  OAI21_X1 U566 ( .B1(n390), .B2(n440), .A(n389), .ZN(n398) );
  INV_X1 U567 ( .A(n391), .ZN(n396) );
  INV_X1 U568 ( .A(n392), .ZN(n394) );
  OAI22_X1 U569 ( .A1(n396), .A2(n558), .B1(n394), .B2(n393), .ZN(n397) );
  AOI211_X1 U570 ( .C1(n400), .C2(n399), .A(n398), .B(n397), .ZN(n402) );
  NAND2_X1 U571 ( .A1(n401), .A2(n464), .ZN(n449) );
  AND4_X1 U572 ( .A1(n403), .A2(n445), .A3(n402), .A4(n449), .ZN(n429) );
  INV_X1 U573 ( .A(n404), .ZN(n412) );
  NAND2_X1 U574 ( .A1(n406), .A2(n405), .ZN(n410) );
  NAND3_X1 U575 ( .A1(n408), .A2(n407), .A3(n501), .ZN(n409) );
  NAND4_X1 U576 ( .A1(n412), .A2(n411), .A3(n410), .A4(n409), .ZN(n426) );
  NAND2_X1 U577 ( .A1(n413), .A2(n17), .ZN(n423) );
  OAI22_X1 U578 ( .A1(n416), .A2(n592), .B1(n539), .B2(n414), .ZN(n417) );
  INV_X1 U579 ( .A(n417), .ZN(n422) );
  OAI21_X1 U580 ( .B1(n420), .B2(n419), .A(n418), .ZN(n421) );
  NAND3_X1 U581 ( .A1(n423), .A2(n422), .A3(n421), .ZN(n425) );
  AOI211_X1 U582 ( .C1(n535), .C2(n426), .A(n425), .B(n424), .ZN(n427) );
  OAI211_X1 U583 ( .C1(n429), .C2(n551), .A(n428), .B(n427), .ZN(
        alu_operator_o[1]) );
  OAI211_X1 U584 ( .C1(n433), .C2(n432), .A(n431), .B(n430), .ZN(n434) );
  OAI21_X1 U585 ( .B1(n435), .B2(n434), .A(n543), .ZN(n460) );
  NOR2_X1 U586 ( .A1(n38), .A2(n288), .ZN(n438) );
  OAI22_X1 U587 ( .A1(n506), .A2(n575), .B1(n436), .B2(n560), .ZN(n437) );
  AOI211_X1 U588 ( .C1(n439), .C2(bmask_a_mux_o[0]), .A(n438), .B(n437), .ZN(
        n459) );
  INV_X1 U589 ( .A(n440), .ZN(n442) );
  NAND3_X1 U590 ( .A1(n442), .A2(n463), .A3(n17), .ZN(n443) );
  NAND4_X1 U591 ( .A1(n31), .A2(n445), .A3(n444), .A4(n443), .ZN(n452) );
  INV_X1 U592 ( .A(n477), .ZN(n447) );
  NAND2_X1 U593 ( .A1(n446), .A2(n480), .ZN(n453) );
  NAND2_X1 U594 ( .A1(n447), .A2(n453), .ZN(n448) );
  OAI211_X1 U595 ( .C1(n451), .C2(n450), .A(n449), .B(n448), .ZN(n517) );
  OAI21_X1 U596 ( .B1(n452), .B2(n517), .A(n516), .ZN(n458) );
  AOI21_X1 U597 ( .B1(n455), .B2(n454), .A(n453), .ZN(n457) );
  OR2_X1 U598 ( .A1(n488), .A2(n575), .ZN(n456) );
  OR2_X1 U599 ( .A1(n457), .A2(n456), .ZN(n521) );
  NAND4_X1 U600 ( .A1(n460), .A2(n459), .A3(n458), .A4(n521), .ZN(
        alu_operator_o[2]) );
  INV_X1 U601 ( .A(n461), .ZN(n466) );
  OAI21_X1 U602 ( .B1(n464), .B2(n463), .A(n462), .ZN(n465) );
  NAND2_X1 U603 ( .A1(n466), .A2(n465), .ZN(n504) );
  INV_X1 U604 ( .A(n467), .ZN(n473) );
  AOI21_X1 U605 ( .B1(n469), .B2(instr_rdata_i[28]), .A(n468), .ZN(n471) );
  OAI22_X1 U606 ( .A1(n473), .A2(n472), .B1(n471), .B2(n470), .ZN(n474) );
  NOR4_X1 U607 ( .A1(n504), .A2(n476), .A3(n475), .A4(n474), .ZN(n530) );
  NOR2_X1 U608 ( .A1(n477), .A2(n480), .ZN(n478) );
  OR2_X1 U609 ( .A1(n479), .A2(n478), .ZN(n495) );
  INV_X1 U610 ( .A(n480), .ZN(n492) );
  OAI22_X1 U611 ( .A1(n482), .A2(n481), .B1(n480), .B2(n488), .ZN(n489) );
  AND3_X1 U612 ( .A1(n485), .A2(n484), .A3(n483), .ZN(n486) );
  OR2_X1 U613 ( .A1(n539), .A2(n545), .ZN(n531) );
  OAI211_X1 U614 ( .C1(n488), .C2(n487), .A(n486), .B(n531), .ZN(n508) );
  OAI21_X1 U615 ( .B1(n489), .B2(n508), .A(n507), .ZN(n490) );
  OAI211_X1 U616 ( .C1(n492), .C2(n38), .A(n490), .B(alu_bmask_a_mux_sel_o), 
        .ZN(n494) );
  AOI211_X1 U617 ( .C1(n516), .C2(n495), .A(n494), .B(n493), .ZN(n496) );
  OAI21_X1 U618 ( .B1(n530), .B2(n572), .A(n496), .ZN(alu_operator_o[3]) );
  INV_X1 U619 ( .A(n497), .ZN(n512) );
  INV_X1 U620 ( .A(n498), .ZN(n499) );
  AOI211_X1 U621 ( .C1(n501), .C2(n541), .A(n500), .B(n499), .ZN(n528) );
  NAND3_X1 U622 ( .A1(n528), .A2(n503), .A3(n502), .ZN(n505) );
  OAI21_X1 U623 ( .B1(n505), .B2(n504), .A(n543), .ZN(n511) );
  INV_X1 U624 ( .A(n506), .ZN(n509) );
  OAI21_X1 U625 ( .B1(n509), .B2(n508), .A(n507), .ZN(n510) );
  OAI211_X1 U626 ( .C1(n512), .C2(n564), .A(n511), .B(n510), .ZN(
        alu_operator_o[4]) );
  INV_X1 U627 ( .A(n513), .ZN(n514) );
  OAI21_X1 U628 ( .B1(n514), .B2(n554), .A(n543), .ZN(n520) );
  AOI22_X1 U629 ( .A1(n517), .A2(n516), .B1(bmask_a_mux_o[0]), .B2(n515), .ZN(
        n519) );
  AND3_X1 U630 ( .A1(n520), .A2(n519), .A3(n518), .ZN(n523) );
  NAND3_X1 U631 ( .A1(n523), .A2(n522), .A3(n521), .ZN(alu_operator_o[5]) );
  NOR3_X1 U632 ( .A1(n526), .A2(n525), .A3(n524), .ZN(n527) );
  AND4_X1 U633 ( .A1(n530), .A2(n529), .A3(n528), .A4(n527), .ZN(n534) );
  OAI211_X1 U634 ( .C1(n534), .C2(n533), .A(n532), .B(n531), .ZN(alu_en_o) );
  NOR3_X1 U635 ( .A1(n536), .A2(n574), .A3(n535), .ZN(n552) );
  NAND2_X1 U636 ( .A1(n548), .A2(n537), .ZN(n538) );
  OAI211_X1 U637 ( .C1(n540), .C2(n539), .A(n552), .B(n538), .ZN(
        alu_bmask_b_mux_sel_o) );
  NAND3_X1 U638 ( .A1(n543), .A2(n542), .A3(n541), .ZN(n544) );
  OAI21_X1 U639 ( .B1(n560), .B2(n545), .A(n544), .ZN(bmask_b_mux_o[0]) );
  NAND3_X1 U640 ( .A1(n548), .A2(n547), .A3(n546), .ZN(n550) );
  NAND4_X1 U641 ( .A1(n552), .A2(n551), .A3(n550), .A4(n549), .ZN(
        bmask_b_mux_o[1]) );
  INV_X1 U642 ( .A(n553), .ZN(n556) );
  NOR4_X1 U643 ( .A1(n557), .A2(n556), .A3(n555), .A4(n554), .ZN(n573) );
  OAI22_X1 U644 ( .A1(n561), .A2(n560), .B1(n559), .B2(n558), .ZN(n562) );
  OR3_X1 U645 ( .A1(alu_operator_o[6]), .A2(n563), .A3(n562), .ZN(n568) );
  AOI21_X1 U646 ( .B1(n566), .B2(n565), .A(n564), .ZN(n567) );
  AOI211_X1 U647 ( .C1(bmask_a_mux_o[0]), .C2(n569), .A(n568), .B(n567), .ZN(
        n571) );
  OAI211_X1 U648 ( .C1(n573), .C2(n572), .A(n571), .B(n570), .ZN(regc_used_o)
         );
  INV_X1 U649 ( .A(n574), .ZN(n577) );
  NOR3_X1 U650 ( .A1(n577), .A2(n576), .A3(n575), .ZN(fencei_insn_o) );
  NOR2_X1 U651 ( .A1(n583), .A2(n578), .ZN(pipe_flush_o) );
  NOR2_X1 U652 ( .A1(n583), .A2(n579), .ZN(dret_dec_o) );
  INV_X1 U653 ( .A(n580), .ZN(n582) );
  NOR3_X1 U654 ( .A1(n583), .A2(n582), .A3(n581), .ZN(uret_insn_o) );
  NOR2_X1 U655 ( .A1(n584), .A2(n583), .ZN(mret_dec_o) );
  INV_X1 U656 ( .A(dret_dec_o), .ZN(n585) );
  NOR2_X1 U657 ( .A1(n585), .A2(n586), .ZN(dret_insn_o) );
  INV_X1 U658 ( .A(mret_dec_o), .ZN(n587) );
  NOR2_X1 U659 ( .A1(n587), .A2(n586), .ZN(mret_insn_o) );
  INV_X2 U136 ( .A(n76), .ZN(n408) );
  NOR2_X2 U26 ( .A1(n35), .A2(n149), .ZN(n336) );
  INV_X1 U10 ( .A(instr_rdata_i[14]), .ZN(n558) );
  CLKBUF_X1 U3 ( .A(instr_rdata_i[5]), .Z(n325) );
  INV_X1 U18 ( .A(n395), .ZN(n288) );
  AND2_X1 U85 ( .A1(n34), .A2(instr_rdata_i[6]), .ZN(n125) );
  OR2_X1 U56 ( .A1(n89), .A2(n56), .ZN(n533) );
  OR2_X1 U8 ( .A1(n89), .A2(n20), .ZN(n488) );
  NOR3_X1 U19 ( .A1(n250), .A2(n574), .A3(n481), .ZN(hwloop_we_o[2]) );
  INV_X1 U142 ( .A(instr_rdata_i[13]), .ZN(n545) );
  MUX2_X1 U11 ( .A(n144), .B(n143), .S(n218), .Z(n149) );
  INV_X1 U12 ( .A(instr_rdata_i[12]), .ZN(n342) );
  AND2_X2 U25 ( .A1(instr_rdata_i[12]), .A2(n591), .ZN(n198) );
  INV_X2 U33 ( .A(instr_rdata_i[13]), .ZN(n591) );
  NAND2_X1 U36 ( .A1(n336), .A2(n46), .ZN(n45) );
  NOR2_X2 U37 ( .A1(n225), .A2(n415), .ZN(hwloop_target_mux_sel_o) );
  OR2_X1 U39 ( .A1(data_misaligned_i), .A2(n575), .ZN(n328) );
  OR2_X1 U43 ( .A1(n446), .A2(n488), .ZN(n598) );
  NOR2_X1 U64 ( .A1(n157), .A2(instr_rdata_i[13]), .ZN(n574) );
  AND2_X1 U79 ( .A1(n163), .A2(n164), .ZN(n597) );
  INV_X1 U100 ( .A(n454), .ZN(n592) );
  CLKBUF_X1 U157 ( .A(instr_rdata_i[6]), .Z(n593) );
  CLKBUF_X1 U312 ( .A(instr_rdata_i[2]), .Z(n594) );
  CLKBUF_X1 U343 ( .A(instr_rdata_i[30]), .Z(n595) );
  CLKBUF_X1 U344 ( .A(jump_target_mux_sel_o[0]), .Z(n596) );
  OAI211_X1 U346 ( .C1(n598), .C2(n254), .A(n165), .B(n597), .ZN(n166) );
  NAND2_X2 U660 ( .A1(n333), .A2(n360), .ZN(n546) );
  NAND3_X1 U661 ( .A1(n168), .A2(n169), .A3(n170), .ZN(illegal_insn_o) );
endmodule


module register_file_test_wrap_ADDR_WIDTH6_FPU0_Zfinx0 ( clk, rst_n, test_en_i, 
        raddr_a_i, rdata_a_o, raddr_b_i, rdata_b_o, raddr_c_i, rdata_c_o, 
        waddr_a_i, wdata_a_i, we_a_i, waddr_b_i, wdata_b_i, we_b_i, BIST, 
        CSN_T, WEN_T, A_T, D_T, Q_T );
  input [5:0] raddr_a_i;
  output [31:0] rdata_a_o;
  input [5:0] raddr_b_i;
  output [31:0] rdata_b_o;
  input [5:0] raddr_c_i;
  output [31:0] rdata_c_o;
  input [5:0] waddr_a_i;
  input [31:0] wdata_a_i;
  input [5:0] waddr_b_i;
  input [31:0] wdata_b_i;
  input [5:0] A_T;
  input [31:0] D_T;
  output [31:0] Q_T;
  input clk, rst_n, test_en_i, we_a_i, we_b_i, BIST, CSN_T, WEN_T;


  riscv_register_file_ADDR_WIDTH6_DATA_WIDTH32_FPU0_Zfinx0 riscv_register_file_i ( 
        .clk(clk), .rst_n(rst_n), .test_en_i(1'b0), .raddr_a_i({1'b0, 
        raddr_a_i[4:0]}), .rdata_a_o(rdata_a_o), .raddr_b_i({1'b0, 
        raddr_b_i[4:0]}), .rdata_b_o(rdata_b_o), .raddr_c_i({1'b0, 
        raddr_c_i[4:0]}), .rdata_c_o(rdata_c_o), .waddr_a_i({1'b0, 
        waddr_a_i[4:0]}), .wdata_a_i(wdata_a_i), .we_a_i(we_a_i), .waddr_b_i({
        1'b0, waddr_b_i[4:0]}), .wdata_b_i(wdata_b_i), .we_b_i(we_b_i) );
endmodule


module SNPS_CLOCK_GATE_HIGH_riscv_if_stage_2_128_0_1a110800_0 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net1, net4;
  assign net1 = EN;
  assign net4 = TE;

  CLKGATETST_X1 latch ( .CK(CLK), .E(net1), .SE(net4), .GCK(ENCLK) );
endmodule


module riscv_compressed_decoder_FPU0 ( instr_i, instr_o, is_compressed_o, 
        illegal_instr_o );
  input [31:0] instr_i;
  output [31:0] instr_o;
  output is_compressed_o, illegal_instr_o;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193;

  NAND2_X1 U3 ( .A1(instr_i[1]), .A2(instr_i[0]), .ZN(is_compressed_o) );
  INV_X1 U4 ( .A(instr_i[3]), .ZN(n109) );
  INV_X1 U5 ( .A(instr_i[13]), .ZN(n142) );
  INV_X1 U6 ( .A(instr_i[0]), .ZN(n64) );
  NOR2_X1 U7 ( .A1(instr_i[1]), .A2(n64), .ZN(n105) );
  INV_X1 U8 ( .A(n105), .ZN(n178) );
  NOR3_X1 U9 ( .A1(instr_i[14]), .A2(n142), .A3(n178), .ZN(n59) );
  INV_X1 U10 ( .A(n59), .ZN(n189) );
  OAI21_X1 U11 ( .B1(n109), .B2(is_compressed_o), .A(n189), .ZN(instr_o[3]) );
  INV_X1 U12 ( .A(instr_i[14]), .ZN(n42) );
  NOR2_X1 U13 ( .A1(instr_i[15]), .A2(n42), .ZN(n143) );
  INV_X1 U14 ( .A(instr_i[1]), .ZN(n32) );
  NOR2_X1 U15 ( .A1(instr_i[0]), .A2(n32), .ZN(n52) );
  NOR2_X1 U16 ( .A1(n52), .A2(n105), .ZN(n76) );
  INV_X1 U17 ( .A(n76), .ZN(n19) );
  INV_X1 U18 ( .A(n52), .ZN(n145) );
  INV_X1 U19 ( .A(instr_i[15]), .ZN(n81) );
  NAND2_X1 U20 ( .A1(n81), .A2(n142), .ZN(n111) );
  INV_X1 U21 ( .A(n111), .ZN(n36) );
  NAND2_X1 U22 ( .A1(n36), .A2(n42), .ZN(n75) );
  NOR2_X1 U23 ( .A1(n145), .A2(n75), .ZN(n106) );
  AOI21_X1 U24 ( .B1(n143), .B2(n19), .A(n106), .ZN(n28) );
  NOR3_X1 U25 ( .A1(instr_i[10]), .A2(instr_i[11]), .A3(instr_i[7]), .ZN(n20)
         );
  INV_X1 U26 ( .A(instr_i[9]), .ZN(n56) );
  NAND2_X1 U27 ( .A1(n20), .A2(n56), .ZN(n34) );
  NOR2_X1 U28 ( .A1(instr_i[8]), .A2(n34), .ZN(n37) );
  INV_X1 U29 ( .A(n37), .ZN(n96) );
  NAND3_X1 U30 ( .A1(n42), .A2(n142), .A3(instr_i[15]), .ZN(n172) );
  NOR2_X1 U31 ( .A1(n178), .A2(n172), .ZN(n22) );
  INV_X1 U32 ( .A(instr_i[12]), .ZN(n182) );
  NAND2_X1 U33 ( .A1(instr_i[10]), .A2(instr_i[11]), .ZN(n175) );
  NOR2_X1 U34 ( .A1(n182), .A2(n175), .ZN(n173) );
  AOI22_X1 U35 ( .A1(n52), .A2(instr_i[13]), .B1(n22), .B2(n173), .ZN(n27) );
  NOR2_X1 U36 ( .A1(instr_i[1]), .A2(instr_i[0]), .ZN(n118) );
  NOR2_X1 U37 ( .A1(instr_i[6]), .A2(instr_i[5]), .ZN(n176) );
  INV_X1 U38 ( .A(n75), .ZN(n83) );
  NAND4_X1 U39 ( .A1(n176), .A2(n83), .A3(n37), .A4(n182), .ZN(n21) );
  NAND3_X1 U40 ( .A1(n142), .A2(n172), .A3(n21), .ZN(n25) );
  NOR2_X1 U41 ( .A1(n145), .A2(n172), .ZN(n38) );
  INV_X1 U42 ( .A(instr_i[4]), .ZN(n41) );
  INV_X1 U43 ( .A(instr_i[2]), .ZN(n134) );
  NAND4_X1 U44 ( .A1(n176), .A2(n109), .A3(n41), .A4(n134), .ZN(n33) );
  NAND2_X1 U45 ( .A1(n38), .A2(n33), .ZN(n73) );
  INV_X1 U46 ( .A(n22), .ZN(n66) );
  NOR2_X1 U47 ( .A1(instr_i[11]), .A2(n66), .ZN(n124) );
  NOR2_X1 U48 ( .A1(n106), .A2(n124), .ZN(n63) );
  AOI221_X1 U49 ( .B1(n73), .B2(n63), .C1(n96), .C2(n63), .A(n182), .ZN(n24)
         );
  NAND3_X1 U50 ( .A1(instr_i[13]), .A2(n105), .A3(n143), .ZN(n184) );
  AOI211_X1 U51 ( .C1(n63), .C2(n184), .A(instr_i[12]), .B(n33), .ZN(n23) );
  AOI211_X1 U52 ( .C1(n118), .C2(n25), .A(n24), .B(n23), .ZN(n26) );
  OAI211_X1 U53 ( .C1(n28), .C2(n96), .A(n27), .B(n26), .ZN(illegal_instr_o)
         );
  NOR2_X1 U54 ( .A1(n42), .A2(instr_i[13]), .ZN(n65) );
  NAND2_X1 U55 ( .A1(n65), .A2(n118), .ZN(n89) );
  NOR2_X1 U56 ( .A1(n81), .A2(n89), .ZN(n132) );
  NAND2_X1 U57 ( .A1(n36), .A2(n118), .ZN(n129) );
  INV_X1 U58 ( .A(n129), .ZN(n131) );
  NOR2_X1 U59 ( .A1(n132), .A2(n131), .ZN(n31) );
  NAND2_X1 U60 ( .A1(instr_i[13]), .A2(n42), .ZN(n29) );
  OAI211_X1 U61 ( .C1(n173), .C2(n172), .A(n111), .B(n29), .ZN(n104) );
  OAI21_X1 U62 ( .B1(instr_i[14]), .B2(n104), .A(instr_i[0]), .ZN(n30) );
  OAI211_X1 U63 ( .C1(instr_i[13]), .C2(n32), .A(n31), .B(n30), .ZN(instr_o[1]) );
  INV_X1 U64 ( .A(n38), .ZN(n43) );
  NOR2_X1 U65 ( .A1(n33), .A2(n43), .ZN(n98) );
  INV_X1 U66 ( .A(n98), .ZN(n45) );
  NOR2_X1 U68 ( .A1(n37), .A2(n45), .ZN(n46) );
  AOI211_X1 U69 ( .C1(instr_i[2]), .C2(n190), .A(n59), .B(n46), .ZN(n35) );
  INV_X1 U70 ( .A(instr_i[8]), .ZN(n188) );
  NOR2_X1 U71 ( .A1(n188), .A2(n34), .ZN(n82) );
  NOR2_X1 U72 ( .A1(n82), .A2(n184), .ZN(n79) );
  INV_X1 U73 ( .A(n79), .ZN(n138) );
  OAI211_X1 U74 ( .C1(instr_i[12]), .C2(n45), .A(n35), .B(n138), .ZN(
        instr_o[2]) );
  INV_X1 U75 ( .A(n184), .ZN(n169) );
  NOR2_X1 U76 ( .A1(n173), .A2(n66), .ZN(n90) );
  INV_X1 U77 ( .A(n90), .ZN(n78) );
  NAND2_X1 U78 ( .A1(n105), .A2(n36), .ZN(n136) );
  NAND3_X1 U79 ( .A1(n38), .A2(instr_i[12]), .A3(n37), .ZN(n39) );
  NAND4_X1 U80 ( .A1(n73), .A2(n78), .A3(n136), .A4(n39), .ZN(n95) );
  AOI211_X1 U81 ( .C1(n83), .C2(n64), .A(n169), .B(n95), .ZN(n40) );
  OAI21_X1 U82 ( .B1(is_compressed_o), .B2(n41), .A(n40), .ZN(instr_o[4]) );
  NAND3_X1 U83 ( .A1(instr_i[15]), .A2(instr_i[14]), .A3(n105), .ZN(n163) );
  INV_X1 U84 ( .A(n163), .ZN(n179) );
  NOR2_X1 U85 ( .A1(n179), .A2(n59), .ZN(n152) );
  NOR4_X1 U86 ( .A1(instr_i[0]), .A2(instr_i[13]), .A3(n81), .A4(n42), .ZN(
        n103) );
  AOI211_X1 U87 ( .C1(n190), .C2(instr_i[5]), .A(n79), .B(n103), .ZN(n44) );
  OR3_X1 U88 ( .A1(n66), .A2(n175), .A3(instr_i[12]), .ZN(n120) );
  NAND4_X1 U89 ( .A1(n152), .A2(n44), .A3(n43), .A4(n120), .ZN(instr_o[5]) );
  INV_X1 U90 ( .A(instr_i[6]), .ZN(n125) );
  OAI211_X1 U91 ( .C1(n125), .C2(is_compressed_o), .A(n152), .B(n45), .ZN(
        instr_o[6]) );
  OAI21_X1 U92 ( .B1(n76), .B2(n111), .A(n73), .ZN(n123) );
  NOR2_X1 U93 ( .A1(n90), .A2(n123), .ZN(n116) );
  NAND2_X1 U94 ( .A1(n116), .A2(is_compressed_o), .ZN(n49) );
  NOR2_X1 U95 ( .A1(n79), .A2(n49), .ZN(n55) );
  INV_X1 U96 ( .A(instr_i[7]), .ZN(n149) );
  AOI22_X1 U97 ( .A1(n131), .A2(instr_i[2]), .B1(n59), .B2(n81), .ZN(n48) );
  OAI21_X1 U98 ( .B1(n179), .B2(n46), .A(instr_i[12]), .ZN(n47) );
  OAI211_X1 U99 ( .C1(n55), .C2(n149), .A(n48), .B(n47), .ZN(instr_o[7]) );
  NAND2_X1 U100 ( .A1(n163), .A2(n129), .ZN(n53) );
  INV_X1 U101 ( .A(n53), .ZN(n51) );
  OAI21_X1 U102 ( .B1(n169), .B2(n49), .A(instr_i[8]), .ZN(n50) );
  OAI21_X1 U103 ( .B1(n51), .B2(n109), .A(n50), .ZN(instr_o[8]) );
  AND2_X1 U104 ( .A1(n52), .A2(n65), .ZN(n133) );
  NAND2_X1 U105 ( .A1(instr_i[15]), .A2(n133), .ZN(n114) );
  AOI22_X1 U106 ( .A1(instr_i[6]), .A2(n132), .B1(instr_i[4]), .B2(n53), .ZN(
        n54) );
  OAI221_X1 U107 ( .B1(n56), .B2(n55), .C1(n56), .C2(n114), .A(n54), .ZN(
        instr_o[9]) );
  NAND3_X1 U108 ( .A1(n138), .A2(is_compressed_o), .A3(n163), .ZN(n57) );
  NOR3_X1 U109 ( .A1(n103), .A2(n123), .A3(n57), .ZN(n58) );
  INV_X1 U110 ( .A(instr_i[10]), .ZN(n92) );
  OAI211_X1 U111 ( .C1(n58), .C2(n92), .A(n129), .B(n78), .ZN(instr_o[10]) );
  INV_X1 U112 ( .A(instr_i[11]), .ZN(n130) );
  NOR2_X1 U113 ( .A1(n58), .A2(n130), .ZN(instr_o[11]) );
  NOR2_X1 U114 ( .A1(instr_i[10]), .A2(n66), .ZN(n137) );
  INV_X1 U115 ( .A(instr_i[5]), .ZN(n115) );
  NOR3_X1 U116 ( .A1(instr_i[12]), .A2(n66), .A3(n115), .ZN(n69) );
  AOI22_X1 U117 ( .A1(n190), .A2(instr_i[12]), .B1(instr_i[6]), .B2(n69), .ZN(
        n60) );
  NAND2_X1 U118 ( .A1(instr_i[12]), .A2(n59), .ZN(n192) );
  OAI211_X1 U119 ( .C1(n134), .C2(n138), .A(n60), .B(n192), .ZN(n61) );
  AOI211_X1 U120 ( .C1(n179), .C2(instr_i[13]), .A(n137), .B(n61), .ZN(n62) );
  NAND2_X1 U121 ( .A1(n63), .A2(n62), .ZN(instr_o[12]) );
  AOI22_X1 U122 ( .A1(n190), .A2(instr_i[13]), .B1(n65), .B2(n64), .ZN(n68) );
  AOI221_X1 U123 ( .B1(instr_i[12]), .B2(instr_i[10]), .C1(n125), .C2(
        instr_i[10]), .A(n66), .ZN(n70) );
  AOI22_X1 U124 ( .A1(instr_i[11]), .A2(n70), .B1(n79), .B2(instr_i[3]), .ZN(
        n67) );
  NAND3_X1 U125 ( .A1(n68), .A2(n67), .A3(n192), .ZN(instr_o[13]) );
  AOI211_X1 U126 ( .C1(instr_i[4]), .C2(n79), .A(n124), .B(n69), .ZN(n72) );
  INV_X1 U127 ( .A(n192), .ZN(n86) );
  AOI211_X1 U128 ( .C1(n190), .C2(instr_i[14]), .A(n86), .B(n70), .ZN(n71) );
  NAND2_X1 U129 ( .A1(n72), .A2(n71), .ZN(instr_o[14]) );
  INV_X1 U130 ( .A(n73), .ZN(n102) );
  AOI21_X1 U131 ( .B1(n102), .B2(instr_i[12]), .A(n98), .ZN(n74) );
  OAI21_X1 U132 ( .B1(n76), .B2(n75), .A(n74), .ZN(n77) );
  INV_X1 U133 ( .A(n77), .ZN(n94) );
  NAND4_X1 U134 ( .A1(n94), .A2(n78), .A3(n89), .A4(n163), .ZN(n87) );
  AOI22_X1 U135 ( .A1(instr_i[7]), .A2(n87), .B1(n79), .B2(instr_i[5]), .ZN(
        n80) );
  OAI211_X1 U136 ( .C1(is_compressed_o), .C2(n81), .A(n80), .B(n192), .ZN(
        instr_o[15]) );
  NAND2_X1 U137 ( .A1(n169), .A2(n82), .ZN(n135) );
  INV_X1 U138 ( .A(n135), .ZN(n162) );
  AOI211_X1 U139 ( .C1(n190), .C2(instr_i[16]), .A(n133), .B(n162), .ZN(n85)
         );
  AOI22_X1 U140 ( .A1(n169), .A2(instr_i[6]), .B1(instr_i[8]), .B2(n87), .ZN(
        n84) );
  NAND2_X1 U141 ( .A1(n118), .A2(n83), .ZN(n154) );
  NAND4_X1 U142 ( .A1(n85), .A2(n84), .A3(n192), .A4(n154), .ZN(instr_o[16])
         );
  NOR2_X1 U143 ( .A1(n138), .A2(n182), .ZN(n165) );
  NOR2_X1 U144 ( .A1(n86), .A2(n165), .ZN(n100) );
  AOI22_X1 U145 ( .A1(instr_i[9]), .A2(n87), .B1(n190), .B2(instr_i[17]), .ZN(
        n88) );
  NAND2_X1 U146 ( .A1(n100), .A2(n88), .ZN(instr_o[17]) );
  NAND2_X1 U147 ( .A1(n89), .A2(n163), .ZN(n146) );
  AOI211_X1 U148 ( .C1(n190), .C2(instr_i[18]), .A(n90), .B(n146), .ZN(n91) );
  OAI211_X1 U149 ( .C1(n94), .C2(n92), .A(n100), .B(n91), .ZN(instr_o[18]) );
  NAND2_X1 U150 ( .A1(n190), .A2(instr_i[19]), .ZN(n93) );
  OAI211_X1 U151 ( .C1(n94), .C2(n130), .A(n100), .B(n93), .ZN(instr_o[19]) );
  NOR3_X1 U152 ( .A1(n103), .A2(n106), .A3(n95), .ZN(n101) );
  NOR2_X1 U153 ( .A1(n182), .A2(n96), .ZN(n97) );
  AOI22_X1 U154 ( .A1(n190), .A2(instr_i[20]), .B1(n98), .B2(n97), .ZN(n99) );
  OAI211_X1 U155 ( .C1(n101), .C2(n134), .A(n100), .B(n99), .ZN(instr_o[20])
         );
  AOI211_X1 U156 ( .C1(n105), .C2(n104), .A(n103), .B(n102), .ZN(n110) );
  INV_X1 U157 ( .A(n106), .ZN(n108) );
  AOI21_X1 U158 ( .B1(n190), .B2(instr_i[21]), .A(n165), .ZN(n107) );
  OAI221_X1 U159 ( .B1(n109), .B2(n110), .C1(n109), .C2(n108), .A(n107), .ZN(
        instr_o[21]) );
  OAI21_X1 U160 ( .B1(n145), .B2(n111), .A(n110), .ZN(n112) );
  AOI22_X1 U161 ( .A1(n190), .A2(instr_i[22]), .B1(instr_i[4]), .B2(n112), 
        .ZN(n113) );
  INV_X1 U162 ( .A(n165), .ZN(n121) );
  OAI211_X1 U163 ( .C1(n129), .C2(n125), .A(n113), .B(n121), .ZN(instr_o[22])
         );
  INV_X1 U164 ( .A(n114), .ZN(n156) );
  NAND2_X1 U165 ( .A1(n189), .A2(n154), .ZN(n170) );
  NOR2_X1 U166 ( .A1(n156), .A2(n170), .ZN(n150) );
  AOI21_X1 U167 ( .B1(n116), .B2(n150), .A(n115), .ZN(n117) );
  AOI211_X1 U168 ( .C1(n190), .C2(instr_i[23]), .A(n117), .B(n132), .ZN(n122)
         );
  NAND4_X1 U169 ( .A1(n143), .A2(instr_i[10]), .A3(n118), .A4(n142), .ZN(n119)
         );
  NAND4_X1 U170 ( .A1(n122), .A2(n121), .A3(n120), .A4(n119), .ZN(instr_o[23])
         );
  NOR4_X1 U171 ( .A1(n156), .A2(n137), .A3(n124), .A4(n123), .ZN(n126) );
  AOI21_X1 U172 ( .B1(n126), .B2(n135), .A(n125), .ZN(n127) );
  AOI211_X1 U173 ( .C1(n190), .C2(instr_i[24]), .A(n127), .B(n165), .ZN(n128)
         );
  OAI221_X1 U174 ( .B1(n130), .B2(n129), .C1(n130), .C2(n189), .A(n128), .ZN(
        instr_o[24]) );
  NOR3_X1 U175 ( .A1(n133), .A2(n132), .A3(n131), .ZN(n141) );
  AOI21_X1 U176 ( .B1(n152), .B2(n135), .A(n134), .ZN(n139) );
  INV_X1 U177 ( .A(n136), .ZN(n180) );
  AOI21_X1 U178 ( .B1(instr_i[11]), .B2(n137), .A(n180), .ZN(n164) );
  AOI21_X1 U179 ( .B1(n164), .B2(n138), .A(n182), .ZN(n151) );
  AOI211_X1 U180 ( .C1(n190), .C2(instr_i[25]), .A(n139), .B(n151), .ZN(n140)
         );
  OAI21_X1 U181 ( .B1(n141), .B2(n182), .A(n140), .ZN(instr_o[25]) );
  NAND2_X1 U182 ( .A1(n143), .A2(n142), .ZN(n144) );
  NOR2_X1 U183 ( .A1(n145), .A2(n144), .ZN(n157) );
  AOI22_X1 U184 ( .A1(n190), .A2(instr_i[26]), .B1(instr_i[2]), .B2(n157), 
        .ZN(n148) );
  AOI221_X1 U185 ( .B1(n162), .B2(instr_i[5]), .C1(n146), .C2(instr_i[5]), .A(
        n151), .ZN(n147) );
  OAI211_X1 U186 ( .C1(n150), .C2(n149), .A(n148), .B(n147), .ZN(instr_o[26])
         );
  INV_X1 U187 ( .A(n151), .ZN(n161) );
  INV_X1 U188 ( .A(n152), .ZN(n153) );
  AOI22_X1 U189 ( .A1(n190), .A2(instr_i[27]), .B1(instr_i[6]), .B2(n153), 
        .ZN(n160) );
  INV_X1 U190 ( .A(n154), .ZN(n155) );
  OAI21_X1 U191 ( .B1(n156), .B2(n155), .A(instr_i[8]), .ZN(n159) );
  OAI21_X1 U192 ( .B1(n162), .B2(n157), .A(instr_i[3]), .ZN(n158) );
  NAND4_X1 U193 ( .A1(n161), .A2(n160), .A3(n159), .A4(n158), .ZN(instr_o[27])
         );
  AOI22_X1 U194 ( .A1(n190), .A2(instr_i[28]), .B1(instr_i[4]), .B2(n162), 
        .ZN(n167) );
  AOI21_X1 U195 ( .B1(n164), .B2(n163), .A(n182), .ZN(n168) );
  AOI211_X1 U196 ( .C1(instr_i[9]), .C2(n170), .A(n168), .B(n165), .ZN(n166)
         );
  NAND2_X1 U197 ( .A1(n167), .A2(n166), .ZN(instr_o[28]) );
  AOI21_X1 U198 ( .B1(instr_i[12]), .B2(n169), .A(n168), .ZN(n191) );
  AOI22_X1 U199 ( .A1(instr_i[10]), .A2(n170), .B1(n190), .B2(instr_i[29]), 
        .ZN(n171) );
  NAND2_X1 U200 ( .A1(n191), .A2(n171), .ZN(instr_o[29]) );
  NOR2_X1 U201 ( .A1(n173), .A2(n172), .ZN(n174) );
  OAI21_X1 U202 ( .B1(n176), .B2(n175), .A(n174), .ZN(n177) );
  NOR2_X1 U203 ( .A1(n178), .A2(n177), .ZN(n181) );
  AOI22_X1 U204 ( .A1(instr_i[10]), .A2(n181), .B1(n190), .B2(instr_i[30]), 
        .ZN(n187) );
  AOI211_X1 U205 ( .C1(instr_i[11]), .C2(n181), .A(n180), .B(n179), .ZN(n183)
         );
  AOI21_X1 U206 ( .B1(n184), .B2(n183), .A(n182), .ZN(n185) );
  INV_X1 U207 ( .A(n185), .ZN(n186) );
  OAI211_X1 U208 ( .C1(n189), .C2(n188), .A(n187), .B(n186), .ZN(instr_o[30])
         );
  NAND2_X1 U209 ( .A1(n190), .A2(instr_i[31]), .ZN(n193) );
  NAND3_X1 U210 ( .A1(n193), .A2(n192), .A3(n191), .ZN(instr_o[31]) );
  INV_X1 U67 ( .A(is_compressed_o), .ZN(n190) );
endmodule


module riscv_hwloop_controller_N_REGS2 ( current_pc_i, hwlp_start_addr_i, 
        hwlp_end_addr_i, hwlp_counter_i, hwlp_dec_cnt_id_i, hwlp_jump_o, 
        hwlp_targ_addr_o, hwlp_dec_cnt_o_1_, hwlp_dec_cnt_o_0_ );
  input [31:0] current_pc_i;
  input [63:0] hwlp_start_addr_i;
  input [63:0] hwlp_end_addr_i;
  input [63:0] hwlp_counter_i;
  input [1:0] hwlp_dec_cnt_id_i;
  output [31:0] hwlp_targ_addr_o;
  output hwlp_jump_o, hwlp_dec_cnt_o_1_, hwlp_dec_cnt_o_0_;
  wire   n165, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n166,
         n167, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201;

  BUF_X2 U3 ( .A(n173), .Z(hwlp_dec_cnt_o_1_) );
  INV_X2 U4 ( .A(n165), .ZN(hwlp_dec_cnt_o_0_) );
  XNOR2_X1 U5 ( .A(current_pc_i[9]), .B(hwlp_end_addr_i[9]), .ZN(n5) );
  XNOR2_X1 U6 ( .A(current_pc_i[12]), .B(hwlp_end_addr_i[12]), .ZN(n4) );
  XNOR2_X1 U7 ( .A(current_pc_i[8]), .B(hwlp_end_addr_i[8]), .ZN(n3) );
  XNOR2_X1 U8 ( .A(current_pc_i[5]), .B(hwlp_end_addr_i[5]), .ZN(n2) );
  NAND4_X1 U9 ( .A1(n5), .A2(n4), .A3(n3), .A4(n2), .ZN(n11) );
  XNOR2_X1 U10 ( .A(current_pc_i[6]), .B(hwlp_end_addr_i[6]), .ZN(n9) );
  XNOR2_X1 U11 ( .A(current_pc_i[4]), .B(hwlp_end_addr_i[4]), .ZN(n8) );
  XNOR2_X1 U12 ( .A(current_pc_i[3]), .B(hwlp_end_addr_i[3]), .ZN(n7) );
  XNOR2_X1 U13 ( .A(current_pc_i[10]), .B(hwlp_end_addr_i[10]), .ZN(n6) );
  NAND4_X1 U14 ( .A1(n9), .A2(n8), .A3(n7), .A4(n6), .ZN(n10) );
  OR2_X1 U15 ( .A1(n11), .A2(n10), .ZN(n22) );
  XNOR2_X1 U16 ( .A(current_pc_i[22]), .B(hwlp_end_addr_i[22]), .ZN(n15) );
  XNOR2_X1 U17 ( .A(current_pc_i[0]), .B(hwlp_end_addr_i[0]), .ZN(n14) );
  XNOR2_X1 U18 ( .A(current_pc_i[19]), .B(hwlp_end_addr_i[19]), .ZN(n13) );
  XNOR2_X1 U19 ( .A(current_pc_i[17]), .B(hwlp_end_addr_i[17]), .ZN(n12) );
  NAND4_X1 U20 ( .A1(n15), .A2(n14), .A3(n13), .A4(n12), .ZN(n21) );
  XNOR2_X1 U21 ( .A(current_pc_i[18]), .B(hwlp_end_addr_i[18]), .ZN(n19) );
  XNOR2_X1 U22 ( .A(current_pc_i[16]), .B(hwlp_end_addr_i[16]), .ZN(n18) );
  XNOR2_X1 U23 ( .A(current_pc_i[7]), .B(hwlp_end_addr_i[7]), .ZN(n17) );
  XNOR2_X1 U24 ( .A(current_pc_i[11]), .B(hwlp_end_addr_i[11]), .ZN(n16) );
  NAND4_X1 U25 ( .A1(n19), .A2(n18), .A3(n17), .A4(n16), .ZN(n20) );
  NOR3_X1 U26 ( .A1(n22), .A2(n21), .A3(n20), .ZN(n76) );
  OR2_X1 U27 ( .A1(hwlp_counter_i[30]), .A2(hwlp_counter_i[3]), .ZN(n23) );
  NOR3_X1 U28 ( .A1(n23), .A2(hwlp_counter_i[29]), .A3(hwlp_counter_i[28]), 
        .ZN(n29) );
  OR2_X1 U29 ( .A1(hwlp_counter_i[22]), .A2(hwlp_counter_i[20]), .ZN(n24) );
  NOR3_X1 U30 ( .A1(n24), .A2(hwlp_counter_i[26]), .A3(hwlp_counter_i[24]), 
        .ZN(n28) );
  OR2_X1 U31 ( .A1(hwlp_counter_i[14]), .A2(hwlp_counter_i[12]), .ZN(n25) );
  NOR3_X1 U32 ( .A1(n25), .A2(hwlp_counter_i[18]), .A3(hwlp_counter_i[16]), 
        .ZN(n27) );
  NOR2_X1 U33 ( .A1(hwlp_counter_i[31]), .A2(hwlp_counter_i[5]), .ZN(n26) );
  NAND4_X1 U34 ( .A1(n29), .A2(n28), .A3(n27), .A4(n26), .ZN(n40) );
  NOR2_X1 U35 ( .A1(hwlp_counter_i[10]), .A2(hwlp_counter_i[8]), .ZN(n33) );
  NOR2_X1 U36 ( .A1(hwlp_counter_i[6]), .A2(hwlp_counter_i[4]), .ZN(n32) );
  NOR2_X1 U37 ( .A1(hwlp_counter_i[25]), .A2(hwlp_counter_i[23]), .ZN(n31) );
  NOR2_X1 U38 ( .A1(hwlp_counter_i[27]), .A2(hwlp_counter_i[2]), .ZN(n30) );
  NAND4_X1 U39 ( .A1(n33), .A2(n32), .A3(n31), .A4(n30), .ZN(n39) );
  NOR2_X1 U40 ( .A1(hwlp_counter_i[21]), .A2(hwlp_counter_i[19]), .ZN(n37) );
  NOR2_X1 U41 ( .A1(hwlp_counter_i[17]), .A2(hwlp_counter_i[15]), .ZN(n36) );
  NOR2_X1 U42 ( .A1(hwlp_counter_i[13]), .A2(hwlp_counter_i[11]), .ZN(n35) );
  NOR2_X1 U43 ( .A1(hwlp_counter_i[9]), .A2(hwlp_counter_i[7]), .ZN(n34) );
  NAND4_X1 U44 ( .A1(n37), .A2(n36), .A3(n35), .A4(n34), .ZN(n38) );
  NOR3_X1 U45 ( .A1(n40), .A2(n39), .A3(n38), .ZN(n44) );
  INV_X1 U46 ( .A(hwlp_counter_i[0]), .ZN(n41) );
  NAND2_X1 U47 ( .A1(hwlp_dec_cnt_id_i[0]), .A2(n41), .ZN(n42) );
  NAND2_X1 U48 ( .A1(n42), .A2(hwlp_counter_i[1]), .ZN(n43) );
  NAND2_X1 U49 ( .A1(n44), .A2(n43), .ZN(n75) );
  INV_X1 U50 ( .A(hwlp_end_addr_i[13]), .ZN(n46) );
  INV_X1 U51 ( .A(hwlp_end_addr_i[20]), .ZN(n45) );
  AOI22_X1 U52 ( .A1(current_pc_i[13]), .A2(n46), .B1(n45), .B2(
        current_pc_i[20]), .ZN(n50) );
  XNOR2_X1 U53 ( .A(current_pc_i[29]), .B(hwlp_end_addr_i[29]), .ZN(n49) );
  XNOR2_X1 U54 ( .A(current_pc_i[30]), .B(hwlp_end_addr_i[30]), .ZN(n48) );
  XNOR2_X1 U55 ( .A(current_pc_i[27]), .B(hwlp_end_addr_i[27]), .ZN(n47) );
  NAND4_X1 U56 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .ZN(n62) );
  INV_X1 U57 ( .A(current_pc_i[14]), .ZN(n60) );
  INV_X1 U58 ( .A(hwlp_end_addr_i[15]), .ZN(n57) );
  INV_X1 U59 ( .A(current_pc_i[15]), .ZN(n52) );
  INV_X1 U60 ( .A(current_pc_i[20]), .ZN(n51) );
  AOI22_X1 U61 ( .A1(n52), .A2(hwlp_end_addr_i[15]), .B1(hwlp_end_addr_i[20]), 
        .B2(n51), .ZN(n55) );
  INV_X1 U62 ( .A(current_pc_i[13]), .ZN(n53) );
  AOI22_X1 U63 ( .A1(n53), .A2(hwlp_end_addr_i[13]), .B1(hwlp_end_addr_i[14]), 
        .B2(n60), .ZN(n54) );
  NAND2_X1 U64 ( .A1(n55), .A2(n54), .ZN(n56) );
  AOI21_X1 U65 ( .B1(n57), .B2(current_pc_i[15]), .A(n56), .ZN(n59) );
  XNOR2_X1 U66 ( .A(current_pc_i[2]), .B(hwlp_end_addr_i[2]), .ZN(n58) );
  OAI211_X1 U67 ( .C1(hwlp_end_addr_i[14]), .C2(n60), .A(n59), .B(n58), .ZN(
        n61) );
  NOR2_X1 U68 ( .A1(n62), .A2(n61), .ZN(n74) );
  XNOR2_X1 U69 ( .A(current_pc_i[28]), .B(hwlp_end_addr_i[28]), .ZN(n66) );
  XNOR2_X1 U70 ( .A(current_pc_i[25]), .B(hwlp_end_addr_i[25]), .ZN(n65) );
  XNOR2_X1 U71 ( .A(current_pc_i[26]), .B(hwlp_end_addr_i[26]), .ZN(n64) );
  XNOR2_X1 U72 ( .A(current_pc_i[23]), .B(hwlp_end_addr_i[23]), .ZN(n63) );
  NAND4_X1 U73 ( .A1(n66), .A2(n65), .A3(n64), .A4(n63), .ZN(n72) );
  XNOR2_X1 U74 ( .A(current_pc_i[31]), .B(hwlp_end_addr_i[31]), .ZN(n70) );
  XNOR2_X1 U75 ( .A(current_pc_i[21]), .B(hwlp_end_addr_i[21]), .ZN(n69) );
  XNOR2_X1 U76 ( .A(current_pc_i[1]), .B(hwlp_end_addr_i[1]), .ZN(n68) );
  XNOR2_X1 U77 ( .A(current_pc_i[24]), .B(hwlp_end_addr_i[24]), .ZN(n67) );
  NAND4_X1 U78 ( .A1(n70), .A2(n69), .A3(n68), .A4(n67), .ZN(n71) );
  NOR2_X1 U79 ( .A1(n72), .A2(n71), .ZN(n73) );
  NAND4_X1 U80 ( .A1(n76), .A2(n75), .A3(n74), .A4(n73), .ZN(n165) );
  INV_X1 U81 ( .A(current_pc_i[4]), .ZN(n89) );
  INV_X1 U82 ( .A(current_pc_i[7]), .ZN(n80) );
  OAI22_X1 U83 ( .A1(hwlp_end_addr_i[36]), .A2(n89), .B1(n80), .B2(
        hwlp_end_addr_i[39]), .ZN(n78) );
  INV_X1 U84 ( .A(current_pc_i[3]), .ZN(n88) );
  INV_X1 U85 ( .A(current_pc_i[5]), .ZN(n91) );
  OAI22_X1 U86 ( .A1(hwlp_end_addr_i[35]), .A2(n88), .B1(n91), .B2(
        hwlp_end_addr_i[37]), .ZN(n77) );
  NOR2_X1 U87 ( .A1(n78), .A2(n77), .ZN(n105) );
  INV_X1 U88 ( .A(current_pc_i[9]), .ZN(n98) );
  INV_X1 U89 ( .A(current_pc_i[2]), .ZN(n79) );
  AOI22_X1 U90 ( .A1(n80), .A2(hwlp_end_addr_i[39]), .B1(n79), .B2(
        hwlp_end_addr_i[34]), .ZN(n81) );
  INV_X1 U91 ( .A(n81), .ZN(n84) );
  INV_X1 U92 ( .A(current_pc_i[31]), .ZN(n124) );
  INV_X1 U93 ( .A(current_pc_i[24]), .ZN(n129) );
  OAI22_X1 U94 ( .A1(n124), .A2(hwlp_end_addr_i[63]), .B1(n129), .B2(
        hwlp_end_addr_i[56]), .ZN(n83) );
  INV_X1 U95 ( .A(current_pc_i[25]), .ZN(n127) );
  INV_X1 U96 ( .A(current_pc_i[26]), .ZN(n128) );
  OAI22_X1 U97 ( .A1(n127), .A2(hwlp_end_addr_i[57]), .B1(n128), .B2(
        hwlp_end_addr_i[58]), .ZN(n82) );
  NOR3_X1 U98 ( .A1(n84), .A2(n83), .A3(n82), .ZN(n97) );
  INV_X1 U99 ( .A(current_pc_i[27]), .ZN(n126) );
  INV_X1 U100 ( .A(current_pc_i[8]), .ZN(n85) );
  OAI22_X1 U101 ( .A1(n126), .A2(hwlp_end_addr_i[59]), .B1(n85), .B2(
        hwlp_end_addr_i[40]), .ZN(n86) );
  INV_X1 U102 ( .A(n86), .ZN(n95) );
  INV_X1 U103 ( .A(current_pc_i[1]), .ZN(n87) );
  AOI22_X1 U104 ( .A1(n88), .A2(hwlp_end_addr_i[35]), .B1(n87), .B2(
        hwlp_end_addr_i[33]), .ZN(n94) );
  AOI22_X1 U105 ( .A1(n98), .A2(hwlp_end_addr_i[41]), .B1(n89), .B2(
        hwlp_end_addr_i[36]), .ZN(n93) );
  INV_X1 U106 ( .A(current_pc_i[6]), .ZN(n90) );
  AOI22_X1 U107 ( .A1(n91), .A2(hwlp_end_addr_i[37]), .B1(hwlp_end_addr_i[38]), 
        .B2(n90), .ZN(n92) );
  AND4_X1 U108 ( .A1(n95), .A2(n94), .A3(n93), .A4(n92), .ZN(n96) );
  OAI211_X1 U109 ( .C1(n98), .C2(hwlp_end_addr_i[41]), .A(n97), .B(n96), .ZN(
        n101) );
  INV_X1 U110 ( .A(hwlp_end_addr_i[40]), .ZN(n99) );
  NOR2_X1 U111 ( .A1(n99), .A2(current_pc_i[8]), .ZN(n100) );
  NOR2_X1 U112 ( .A1(n101), .A2(n100), .ZN(n104) );
  XNOR2_X1 U113 ( .A(current_pc_i[12]), .B(hwlp_end_addr_i[44]), .ZN(n103) );
  XNOR2_X1 U114 ( .A(current_pc_i[10]), .B(hwlp_end_addr_i[42]), .ZN(n102) );
  NAND4_X1 U115 ( .A1(n105), .A2(n104), .A3(n103), .A4(n102), .ZN(n111) );
  XNOR2_X1 U116 ( .A(current_pc_i[20]), .B(hwlp_end_addr_i[52]), .ZN(n109) );
  XNOR2_X1 U117 ( .A(current_pc_i[15]), .B(hwlp_end_addr_i[47]), .ZN(n108) );
  XNOR2_X1 U118 ( .A(current_pc_i[13]), .B(hwlp_end_addr_i[45]), .ZN(n107) );
  XNOR2_X1 U119 ( .A(current_pc_i[14]), .B(hwlp_end_addr_i[46]), .ZN(n106) );
  NAND4_X1 U120 ( .A1(n109), .A2(n108), .A3(n107), .A4(n106), .ZN(n110) );
  NOR2_X1 U121 ( .A1(n111), .A2(n110), .ZN(n166) );
  XNOR2_X1 U122 ( .A(current_pc_i[21]), .B(hwlp_end_addr_i[53]), .ZN(n115) );
  XNOR2_X1 U123 ( .A(current_pc_i[0]), .B(hwlp_end_addr_i[32]), .ZN(n114) );
  XNOR2_X1 U124 ( .A(current_pc_i[22]), .B(hwlp_end_addr_i[54]), .ZN(n113) );
  XNOR2_X1 U125 ( .A(current_pc_i[18]), .B(hwlp_end_addr_i[50]), .ZN(n112) );
  NAND4_X1 U126 ( .A1(n115), .A2(n114), .A3(n113), .A4(n112), .ZN(n121) );
  XNOR2_X1 U127 ( .A(current_pc_i[19]), .B(hwlp_end_addr_i[51]), .ZN(n119) );
  XNOR2_X1 U128 ( .A(current_pc_i[17]), .B(hwlp_end_addr_i[49]), .ZN(n118) );
  XNOR2_X1 U129 ( .A(current_pc_i[16]), .B(hwlp_end_addr_i[48]), .ZN(n117) );
  XNOR2_X1 U130 ( .A(current_pc_i[11]), .B(hwlp_end_addr_i[43]), .ZN(n116) );
  NAND4_X1 U131 ( .A1(n119), .A2(n118), .A3(n117), .A4(n116), .ZN(n120) );
  NOR2_X1 U132 ( .A1(n121), .A2(n120), .ZN(n164) );
  INV_X1 U133 ( .A(hwlp_end_addr_i[34]), .ZN(n123) );
  INV_X1 U134 ( .A(hwlp_end_addr_i[33]), .ZN(n122) );
  AOI22_X1 U135 ( .A1(current_pc_i[2]), .A2(n123), .B1(n122), .B2(
        current_pc_i[1]), .ZN(n133) );
  INV_X1 U136 ( .A(hwlp_end_addr_i[38]), .ZN(n125) );
  AOI22_X1 U137 ( .A1(current_pc_i[6]), .A2(n125), .B1(n124), .B2(
        hwlp_end_addr_i[63]), .ZN(n132) );
  AOI22_X1 U138 ( .A1(hwlp_end_addr_i[57]), .A2(n127), .B1(n126), .B2(
        hwlp_end_addr_i[59]), .ZN(n131) );
  AOI22_X1 U139 ( .A1(hwlp_end_addr_i[56]), .A2(n129), .B1(n128), .B2(
        hwlp_end_addr_i[58]), .ZN(n130) );
  NAND4_X1 U140 ( .A1(n133), .A2(n132), .A3(n131), .A4(n130), .ZN(n139) );
  XNOR2_X1 U141 ( .A(current_pc_i[29]), .B(hwlp_end_addr_i[61]), .ZN(n137) );
  XNOR2_X1 U142 ( .A(current_pc_i[30]), .B(hwlp_end_addr_i[62]), .ZN(n136) );
  XNOR2_X1 U143 ( .A(current_pc_i[23]), .B(hwlp_end_addr_i[55]), .ZN(n135) );
  XNOR2_X1 U144 ( .A(current_pc_i[28]), .B(hwlp_end_addr_i[60]), .ZN(n134) );
  NAND4_X1 U145 ( .A1(n137), .A2(n136), .A3(n135), .A4(n134), .ZN(n138) );
  NOR2_X1 U146 ( .A1(n139), .A2(n138), .ZN(n163) );
  OR2_X1 U147 ( .A1(hwlp_counter_i[62]), .A2(hwlp_counter_i[35]), .ZN(n140) );
  NOR3_X1 U148 ( .A1(n140), .A2(hwlp_counter_i[61]), .A3(hwlp_counter_i[60]), 
        .ZN(n146) );
  OR2_X1 U149 ( .A1(hwlp_counter_i[54]), .A2(hwlp_counter_i[52]), .ZN(n141) );
  NOR3_X1 U150 ( .A1(n141), .A2(hwlp_counter_i[58]), .A3(hwlp_counter_i[56]), 
        .ZN(n145) );
  OR2_X1 U151 ( .A1(hwlp_counter_i[46]), .A2(hwlp_counter_i[44]), .ZN(n142) );
  NOR3_X1 U152 ( .A1(n142), .A2(hwlp_counter_i[50]), .A3(hwlp_counter_i[48]), 
        .ZN(n144) );
  NOR2_X1 U153 ( .A1(hwlp_counter_i[63]), .A2(hwlp_counter_i[37]), .ZN(n143)
         );
  NAND4_X1 U154 ( .A1(n146), .A2(n145), .A3(n144), .A4(n143), .ZN(n157) );
  NOR2_X1 U155 ( .A1(hwlp_counter_i[42]), .A2(hwlp_counter_i[40]), .ZN(n150)
         );
  NOR2_X1 U156 ( .A1(hwlp_counter_i[38]), .A2(hwlp_counter_i[36]), .ZN(n149)
         );
  NOR2_X1 U157 ( .A1(hwlp_counter_i[57]), .A2(hwlp_counter_i[55]), .ZN(n148)
         );
  NOR2_X1 U158 ( .A1(hwlp_counter_i[59]), .A2(hwlp_counter_i[34]), .ZN(n147)
         );
  NAND4_X1 U159 ( .A1(n150), .A2(n149), .A3(n148), .A4(n147), .ZN(n156) );
  NOR2_X1 U160 ( .A1(hwlp_counter_i[53]), .A2(hwlp_counter_i[51]), .ZN(n154)
         );
  NOR2_X1 U161 ( .A1(hwlp_counter_i[49]), .A2(hwlp_counter_i[47]), .ZN(n153)
         );
  NOR2_X1 U162 ( .A1(hwlp_counter_i[45]), .A2(hwlp_counter_i[43]), .ZN(n152)
         );
  NOR2_X1 U163 ( .A1(hwlp_counter_i[41]), .A2(hwlp_counter_i[39]), .ZN(n151)
         );
  NAND4_X1 U164 ( .A1(n154), .A2(n153), .A3(n152), .A4(n151), .ZN(n155) );
  NOR3_X1 U165 ( .A1(n157), .A2(n156), .A3(n155), .ZN(n161) );
  INV_X1 U166 ( .A(hwlp_counter_i[32]), .ZN(n158) );
  NAND2_X1 U167 ( .A1(hwlp_dec_cnt_id_i[1]), .A2(n158), .ZN(n159) );
  NAND2_X1 U168 ( .A1(n159), .A2(hwlp_counter_i[33]), .ZN(n160) );
  NAND2_X1 U169 ( .A1(n161), .A2(n160), .ZN(n162) );
  NAND4_X1 U170 ( .A1(n166), .A2(n164), .A3(n163), .A4(n162), .ZN(n201) );
  NOR2_X1 U171 ( .A1(hwlp_dec_cnt_o_0_), .A2(n201), .ZN(n173) );
  AOI22_X1 U172 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[33]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[1]), .ZN(n167) );
  INV_X1 U173 ( .A(n167), .ZN(hwlp_targ_addr_o[1]) );
  AOI22_X1 U174 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[32]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[0]), .ZN(n169) );
  INV_X1 U175 ( .A(n169), .ZN(hwlp_targ_addr_o[0]) );
  AOI22_X1 U176 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[34]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[2]), .ZN(n170) );
  INV_X1 U177 ( .A(n170), .ZN(hwlp_targ_addr_o[2]) );
  AOI22_X1 U178 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[35]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[3]), .ZN(n171) );
  INV_X1 U179 ( .A(n171), .ZN(hwlp_targ_addr_o[3]) );
  AOI22_X1 U180 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[51]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[19]), .ZN(n172) );
  INV_X1 U181 ( .A(n172), .ZN(hwlp_targ_addr_o[19]) );
  AOI22_X1 U182 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[52]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[20]), .ZN(n174) );
  INV_X1 U183 ( .A(n174), .ZN(hwlp_targ_addr_o[20]) );
  AOI22_X1 U184 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[53]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[21]), .ZN(n175) );
  INV_X1 U185 ( .A(n175), .ZN(hwlp_targ_addr_o[21]) );
  AOI22_X1 U186 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[54]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[22]), .ZN(n176) );
  INV_X1 U187 ( .A(n176), .ZN(hwlp_targ_addr_o[22]) );
  AOI22_X1 U188 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[56]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[24]), .ZN(n177) );
  INV_X1 U189 ( .A(n177), .ZN(hwlp_targ_addr_o[24]) );
  AOI22_X1 U190 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[55]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[23]), .ZN(n178) );
  INV_X1 U191 ( .A(n178), .ZN(hwlp_targ_addr_o[23]) );
  AOI22_X1 U192 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[57]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[25]), .ZN(n179) );
  INV_X1 U193 ( .A(n179), .ZN(hwlp_targ_addr_o[25]) );
  AOI22_X1 U194 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[58]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[26]), .ZN(n180) );
  INV_X1 U195 ( .A(n180), .ZN(hwlp_targ_addr_o[26]) );
  AOI22_X1 U196 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[44]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[12]), .ZN(n181) );
  INV_X1 U197 ( .A(n181), .ZN(hwlp_targ_addr_o[12]) );
  AOI22_X1 U198 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[43]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[11]), .ZN(n182) );
  INV_X1 U199 ( .A(n182), .ZN(hwlp_targ_addr_o[11]) );
  AOI22_X1 U200 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[46]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[14]), .ZN(n183) );
  INV_X1 U201 ( .A(n183), .ZN(hwlp_targ_addr_o[14]) );
  AOI22_X1 U202 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[45]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[13]), .ZN(n184) );
  INV_X1 U203 ( .A(n184), .ZN(hwlp_targ_addr_o[13]) );
  AOI22_X1 U204 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[48]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[16]), .ZN(n185) );
  INV_X1 U205 ( .A(n185), .ZN(hwlp_targ_addr_o[16]) );
  AOI22_X1 U206 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[47]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[15]), .ZN(n186) );
  INV_X1 U207 ( .A(n186), .ZN(hwlp_targ_addr_o[15]) );
  AOI22_X1 U208 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[49]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[17]), .ZN(n187) );
  INV_X1 U209 ( .A(n187), .ZN(hwlp_targ_addr_o[17]) );
  AOI22_X1 U210 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[50]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[18]), .ZN(n188) );
  INV_X1 U211 ( .A(n188), .ZN(hwlp_targ_addr_o[18]) );
  AOI22_X1 U212 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[40]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[8]), .ZN(n189) );
  INV_X1 U213 ( .A(n189), .ZN(hwlp_targ_addr_o[8]) );
  AOI22_X1 U214 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[39]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[7]), .ZN(n190) );
  INV_X1 U215 ( .A(n190), .ZN(hwlp_targ_addr_o[7]) );
  AOI22_X1 U216 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[42]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[10]), .ZN(n191) );
  INV_X1 U217 ( .A(n191), .ZN(hwlp_targ_addr_o[10]) );
  AOI22_X1 U218 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[41]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[9]), .ZN(n192) );
  INV_X1 U219 ( .A(n192), .ZN(hwlp_targ_addr_o[9]) );
  AOI22_X1 U220 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[36]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[4]), .ZN(n193) );
  INV_X1 U221 ( .A(n193), .ZN(hwlp_targ_addr_o[4]) );
  AOI22_X1 U222 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[37]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[5]), .ZN(n194) );
  INV_X1 U223 ( .A(n194), .ZN(hwlp_targ_addr_o[5]) );
  AOI22_X1 U224 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[38]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[6]), .ZN(n195) );
  INV_X1 U225 ( .A(n195), .ZN(hwlp_targ_addr_o[6]) );
  AOI22_X1 U226 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[63]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[31]), .ZN(n196) );
  INV_X1 U227 ( .A(n196), .ZN(hwlp_targ_addr_o[31]) );
  AOI22_X1 U228 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[59]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[27]), .ZN(n197) );
  INV_X1 U229 ( .A(n197), .ZN(hwlp_targ_addr_o[27]) );
  AOI22_X1 U230 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[60]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[28]), .ZN(n198) );
  INV_X1 U231 ( .A(n198), .ZN(hwlp_targ_addr_o[28]) );
  AOI22_X1 U232 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[61]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[29]), .ZN(n199) );
  INV_X1 U233 ( .A(n199), .ZN(hwlp_targ_addr_o[29]) );
  AOI22_X1 U234 ( .A1(hwlp_dec_cnt_o_1_), .A2(hwlp_start_addr_i[62]), .B1(
        hwlp_dec_cnt_o_0_), .B2(hwlp_start_addr_i[30]), .ZN(n200) );
  INV_X1 U235 ( .A(n200), .ZN(hwlp_targ_addr_o[30]) );
  NAND2_X1 U236 ( .A1(n201), .A2(n165), .ZN(hwlp_jump_o) );
endmodule


module riscv_prefetch_L0_buffer ( clk, rst_n, req_i, branch_i, addr_i, 
        hwloop_i, hwloop_target_i, ready_i, valid_o, rdata_o, addr_o, 
        is_hwlp_o, instr_req_o, instr_addr_o, instr_gnt_i, instr_rvalid_i, 
        instr_rdata_i, busy_o );
  input [31:0] addr_i;
  input [31:0] hwloop_target_i;
  output [31:0] rdata_o;
  output [31:0] addr_o;
  output [31:0] instr_addr_o;
  input [127:0] instr_rdata_i;
  input clk, rst_n, req_i, branch_i, hwloop_i, ready_i, instr_gnt_i,
         instr_rvalid_i;
  output valid_o, is_hwlp_o, instr_req_o, busy_o;
  wire   n_0_net_, fetch_gnt, fetch_valid, is_hwlp_n, is_hwlp_q, n792, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n7, n8, n9, n10, n12, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n528, n529, n530, n531, n532,
         n533, n537, n538, n539, n540, n541, n542, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n560, n561,
         n562, n563, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n578, n579, n580, n581, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n594, n597, n598, n599, n600, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n615, n616, n617,
         n618, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n633, n634, n635, n636, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n651, n652, n653, n654, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n669, n670, n671, n672, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n687, n688,
         n689, n690, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n705, n706, n707, n708, n710, n711, n712, n713, n714, n715,
         n720, n721, n722, n723, n724, n725, n730, n731, n732, n733, n735,
         n736, n737, n738, n739, n740, n744, n745, n746, n747, n748, n750,
         n751, n752, n753, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n793, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n863, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1203, n1204, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1224, n1225;
  wire   [31:2] addr_real_next;
  wire   [126:0] rdata_L0;
  wire   [3:1] addr_L0;
  wire   [31:0] rdata_last_q;
  wire   [3:0] NS;
  wire   [3:0] CS;
  wire   [31:0] addr_n;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32;

  INV_X1 U11 ( .A(n29), .ZN(n30) );
  OR2_X1 U12 ( .A1(n28), .A2(n9), .ZN(n24) );
  XOR2_X1 U13 ( .A(n445), .B(n834), .Z(n8) );
  XOR2_X1 U14 ( .A(n420), .B(n844), .Z(n9) );
  XOR2_X1 U15 ( .A(n424), .B(n831), .Z(n10) );
  INV_X2 U17 ( .A(n314), .ZN(n265) );
  NOR2_X2 U21 ( .A1(n537), .A2(n306), .ZN(n31) );
  INV_X1 U22 ( .A(n484), .ZN(n23) );
  INV_X1 U23 ( .A(n455), .ZN(n21) );
  NOR2_X2 U24 ( .A1(n871), .A2(n306), .ZN(n755) );
  INV_X1 U25 ( .A(n421), .ZN(n25) );
  AND2_X1 U27 ( .A1(n50), .A2(n49), .ZN(n48) );
  INV_X1 U28 ( .A(n412), .ZN(n27) );
  OR2_X1 U29 ( .A1(n381), .A2(n8), .ZN(n44) );
  NAND2_X1 U30 ( .A1(n19), .A2(n48), .ZN(n825) );
  NAND2_X1 U31 ( .A1(ready_i), .A2(n37), .ZN(n19) );
  OAI21_X1 U32 ( .B1(n509), .B2(n21), .A(n20), .ZN(addr_real_next[18]) );
  NAND2_X1 U33 ( .A1(n30), .A2(n454), .ZN(n20) );
  INV_X2 U34 ( .A(n28), .ZN(n854) );
  MUX2_X1 U35 ( .A(n828), .B(n410), .S(n381), .Z(addr_real_next[4]) );
  OAI21_X1 U36 ( .B1(n854), .B2(n23), .A(n22), .ZN(addr_real_next[24]) );
  NAND2_X1 U37 ( .A1(n854), .A2(n483), .ZN(n22) );
  OAI21_X1 U38 ( .B1(n854), .B2(n25), .A(n24), .ZN(addr_real_next[9]) );
  OAI21_X1 U39 ( .B1(n854), .B2(n27), .A(n26), .ZN(addr_real_next[5]) );
  NAND2_X1 U40 ( .A1(n854), .A2(n411), .ZN(n26) );
  OR2_X1 U41 ( .A1(n381), .A2(n10), .ZN(n58) );
  AND2_X1 U42 ( .A1(n39), .A2(n124), .ZN(n29) );
  INV_X1 U43 ( .A(n432), .ZN(n45) );
  INV_X1 U44 ( .A(n423), .ZN(n59) );
  INV_X1 U45 ( .A(n358), .ZN(n55) );
  NOR2_X1 U46 ( .A1(n33), .A2(n51), .ZN(n50) );
  INV_X1 U47 ( .A(n130), .ZN(n51) );
  NOR2_X1 U48 ( .A1(n358), .A2(n56), .ZN(n359) );
  NOR2_X2 U49 ( .A1(n546), .A2(n769), .ZN(n782) );
  CLKBUF_X1 U50 ( .A(addr_i[28]), .Z(n209) );
  CLKBUF_X1 U52 ( .A(addr_i[31]), .Z(n192) );
  CLKBUF_X1 U53 ( .A(addr_i[26]), .Z(n216) );
  CLKBUF_X1 U54 ( .A(addr_i[25]), .Z(n40) );
  CLKBUF_X1 U55 ( .A(addr_i[22]), .Z(n231) );
  CLKBUF_X1 U56 ( .A(addr_i[20]), .Z(n241) );
  CLKBUF_X1 U57 ( .A(addr_i[19]), .Z(n245) );
  CLKBUF_X1 U59 ( .A(addr_i[17]), .Z(n253) );
  CLKBUF_X1 U60 ( .A(addr_i[16]), .Z(n260) );
  CLKBUF_X1 U61 ( .A(addr_i[14]), .Z(n270) );
  CLKBUF_X1 U62 ( .A(addr_i[10]), .Z(n285) );
  CLKBUF_X1 U63 ( .A(addr_i[9]), .Z(n289) );
  CLKBUF_X1 U64 ( .A(addr_i[8]), .Z(n295) );
  CLKBUF_X1 U66 ( .A(rdata_L0[112]), .Z(n41) );
  INV_X2 U67 ( .A(n765), .ZN(n537) );
  NOR2_X2 U68 ( .A1(n82), .A2(n765), .ZN(n32) );
  AND3_X1 U69 ( .A1(n339), .A2(n123), .A3(n787), .ZN(n33) );
  NOR2_X2 U70 ( .A1(n537), .A2(n167), .ZN(n34) );
  OR2_X1 U71 ( .A1(n57), .A2(n52), .ZN(n35) );
  OR2_X1 U72 ( .A1(n57), .A2(n54), .ZN(n36) );
  AND2_X1 U73 ( .A1(n43), .A2(n383), .ZN(n37) );
  NAND2_X1 U75 ( .A1(n39), .A2(addr_o[2]), .ZN(addr_real_next[2]) );
  OAI21_X2 U76 ( .B1(n885), .B2(n537), .A(n83), .ZN(rdata_o[12]) );
  NOR2_X2 U77 ( .A1(n537), .A2(n166), .ZN(n762) );
  OR3_X1 U78 ( .A1(n537), .A2(addr_o[2]), .A3(n60), .ZN(n761) );
  INV_X1 U79 ( .A(n761), .ZN(n42) );
  OAI21_X1 U80 ( .B1(n509), .B2(n45), .A(n44), .ZN(addr_real_next[12]) );
  MUX2_X1 U81 ( .A(n418), .B(n419), .S(n381), .Z(addr_real_next[7]) );
  INV_X2 U83 ( .A(n29), .ZN(n509) );
  NAND2_X1 U85 ( .A1(rdata_L0[95]), .A2(n755), .ZN(n105) );
  MUX2_X1 U86 ( .A(n437), .B(n438), .S(n28), .Z(addr_real_next[14]) );
  NAND2_X1 U87 ( .A1(n383), .A2(n123), .ZN(n49) );
  NAND2_X1 U88 ( .A1(n893), .A2(n41), .ZN(n57) );
  NAND2_X1 U89 ( .A1(n123), .A2(addr_o[1]), .ZN(n52) );
  NOR2_X1 U90 ( .A1(n57), .A2(n53), .ZN(n365) );
  NAND3_X1 U91 ( .A1(addr_L0[2]), .A2(addr_L0[1]), .A3(addr_L0[3]), .ZN(n53)
         );
  NAND3_X1 U92 ( .A1(hwloop_target_i[2]), .A2(hwloop_target_i[1]), .A3(
        hwloop_target_i[3]), .ZN(n54) );
  NAND2_X1 U93 ( .A1(n55), .A2(n57), .ZN(n176) );
  NOR2_X1 U94 ( .A1(n57), .A2(n400), .ZN(n56) );
  OAI21_X1 U95 ( .B1(n509), .B2(n59), .A(n58), .ZN(addr_real_next[10]) );
  OR2_X1 U96 ( .A1(n788), .A2(CS[2]), .ZN(n149) );
  INV_X1 U97 ( .A(n149), .ZN(n142) );
  NAND2_X1 U98 ( .A1(n142), .A2(CS[1]), .ZN(n87) );
  OR2_X1 U99 ( .A1(n87), .A2(CS[3]), .ZN(n141) );
  OR2_X1 U100 ( .A1(n829), .A2(CS[1]), .ZN(n392) );
  OAI211_X1 U101 ( .C1(n149), .C2(n787), .A(n141), .B(n392), .ZN(n538) );
  NAND2_X1 U102 ( .A1(addr_o[3]), .A2(addr_o[2]), .ZN(n306) );
  INV_X1 U103 ( .A(n872), .ZN(n64) );
  NAND2_X1 U104 ( .A1(n871), .A2(rdata_last_q[0]), .ZN(n103) );
  INV_X1 U105 ( .A(n103), .ZN(n62) );
  NAND3_X1 U106 ( .A1(n827), .A2(addr_o[3]), .A3(addr_o[2]), .ZN(n61) );
  AOI21_X1 U107 ( .B1(n62), .B2(rdata_last_q[1]), .A(n61), .ZN(n63) );
  AND2_X1 U108 ( .A1(n871), .A2(rdata_last_q[17]), .ZN(n116) );
  NOR2_X1 U109 ( .A1(n871), .A2(n60), .ZN(n66) );
  INV_X1 U110 ( .A(n66), .ZN(n65) );
  OAI22_X1 U111 ( .A1(n116), .A2(n855), .B1(rdata_L0[80]), .B2(n65), .ZN(n71)
         );
  INV_X1 U113 ( .A(n756), .ZN(n777) );
  INV_X1 U114 ( .A(n116), .ZN(n69) );
  NAND2_X1 U115 ( .A1(n871), .A2(n830), .ZN(n67) );
  NAND4_X1 U116 ( .A1(n67), .A2(addr_o[3]), .A3(addr_o[1]), .A4(n826), .ZN(n68) );
  AOI21_X1 U117 ( .B1(n777), .B2(n69), .A(n68), .ZN(n70) );
  NAND2_X1 U118 ( .A1(addr_o[6]), .A2(addr_o[7]), .ZN(n194) );
  NAND2_X1 U119 ( .A1(addr_o[5]), .A2(addr_o[4]), .ZN(n413) );
  NOR2_X1 U120 ( .A1(n194), .A2(n413), .ZN(n430) );
  INV_X1 U121 ( .A(n430), .ZN(n422) );
  XOR2_X1 U122 ( .A(n422), .B(n832), .Z(n72) );
  NOR2_X1 U123 ( .A1(n306), .A2(n413), .ZN(n195) );
  INV_X1 U124 ( .A(n195), .ZN(n302) );
  NOR2_X1 U125 ( .A1(n302), .A2(n194), .ZN(n291) );
  XNOR2_X1 U126 ( .A(n291), .B(n832), .ZN(n296) );
  MUX2_X1 U127 ( .A(n72), .B(n296), .S(n381), .Z(addr_real_next[8]) );
  AOI22_X1 U129 ( .A1(rdata_L0[123]), .A2(n755), .B1(rdata_last_q[28]), .B2(
        n871), .ZN(n76) );
  OR2_X1 U130 ( .A1(addr_o[2]), .A2(addr_o[3]), .ZN(n166) );
  NOR2_X1 U131 ( .A1(n871), .A2(n166), .ZN(n774) );
  NAND2_X1 U133 ( .A1(rdata_L0[28]), .A2(n774), .ZN(n75) );
  NAND2_X1 U134 ( .A1(rdata_L0[91]), .A2(n756), .ZN(n74) );
  OR2_X1 U135 ( .A1(n826), .A2(addr_o[3]), .ZN(n167) );
  NOR2_X1 U136 ( .A1(n871), .A2(n167), .ZN(n773) );
  NAND2_X1 U137 ( .A1(rdata_L0[60]), .A2(n773), .ZN(n73) );
  OAI21_X1 U140 ( .B1(n392), .B2(CS[3]), .A(addr_o[1]), .ZN(n77) );
  INV_X1 U141 ( .A(n77), .ZN(n78) );
  AND2_X1 U142 ( .A1(n141), .A2(n78), .ZN(n765) );
  INV_X1 U143 ( .A(rdata_L0[76]), .ZN(n81) );
  NAND2_X1 U145 ( .A1(rdata_L0[44]), .A2(n744), .ZN(n80) );
  AOI22_X1 U146 ( .A1(rdata_L0[12]), .A2(n892), .B1(rdata_last_q[12]), .B2(
        n871), .ZN(n79) );
  OAI211_X1 U147 ( .C1(n81), .C2(n777), .A(n80), .B(n79), .ZN(n720) );
  INV_X1 U148 ( .A(n755), .ZN(n82) );
  AOI22_X1 U149 ( .A1(n720), .A2(n537), .B1(rdata_L0[107]), .B2(n32), .ZN(n83)
         );
  INV_X1 U150 ( .A(n306), .ZN(n123) );
  OR2_X1 U151 ( .A1(CS[2]), .A2(CS[0]), .ZN(n84) );
  NOR2_X1 U152 ( .A1(n84), .A2(n787), .ZN(n383) );
  INV_X1 U153 ( .A(n383), .ZN(n342) );
  NAND2_X1 U154 ( .A1(CS[1]), .A2(CS[2]), .ZN(n393) );
  INV_X1 U155 ( .A(n393), .ZN(n345) );
  NOR2_X1 U156 ( .A1(CS[3]), .A2(CS[0]), .ZN(n85) );
  AOI22_X1 U157 ( .A1(n383), .A2(n793), .B1(n345), .B2(n85), .ZN(n130) );
  NOR2_X1 U158 ( .A1(n149), .A2(CS[1]), .ZN(n339) );
  OR2_X1 U159 ( .A1(CS[3]), .A2(CS[1]), .ZN(n86) );
  AND2_X1 U160 ( .A1(fetch_valid), .A2(CS[0]), .ZN(n346) );
  NAND2_X1 U161 ( .A1(CS[1]), .A2(CS[3]), .ZN(n90) );
  OAI211_X1 U162 ( .C1(n35), .C2(n86), .A(n346), .B(n90), .ZN(n89) );
  INV_X1 U163 ( .A(n87), .ZN(n88) );
  NOR2_X1 U164 ( .A1(n392), .A2(n788), .ZN(n390) );
  NOR2_X1 U165 ( .A1(n88), .A2(n390), .ZN(n337) );
  OAI211_X1 U166 ( .C1(CS[1]), .C2(CS[2]), .A(n393), .B(CS[3]), .ZN(n91) );
  NAND3_X1 U167 ( .A1(n89), .A2(n337), .A3(n91), .ZN(n125) );
  INV_X1 U168 ( .A(branch_i), .ZN(n172) );
  AND2_X1 U169 ( .A1(n125), .A2(n172), .ZN(valid_o) );
  OAI211_X1 U170 ( .C1(n345), .C2(CS[3]), .A(CS[0]), .B(n90), .ZN(n92) );
  NAND2_X1 U171 ( .A1(n92), .A2(n91), .ZN(n93) );
  AND2_X1 U172 ( .A1(hwloop_i), .A2(n93), .ZN(n171) );
  INV_X1 U173 ( .A(n171), .ZN(n94) );
  NAND4_X1 U174 ( .A1(n787), .A2(n829), .A3(n788), .A4(CS[1]), .ZN(n158) );
  NAND2_X1 U175 ( .A1(n94), .A2(n158), .ZN(n_0_net_) );
  INV_X1 U176 ( .A(n854), .ZN(n174) );
  XNOR2_X1 U177 ( .A(n60), .B(addr_o[2]), .ZN(n315) );
  AND2_X1 U178 ( .A1(n174), .A2(n315), .ZN(addr_real_next[3]) );
  AOI22_X1 U179 ( .A1(rdata_L0[124]), .A2(n755), .B1(rdata_last_q[29]), .B2(
        n871), .ZN(n98) );
  NAND2_X1 U180 ( .A1(rdata_L0[29]), .A2(n774), .ZN(n97) );
  NAND2_X1 U181 ( .A1(rdata_L0[92]), .A2(n756), .ZN(n96) );
  NAND2_X1 U182 ( .A1(rdata_L0[61]), .A2(n773), .ZN(n95) );
  INV_X1 U185 ( .A(rdata_L0[77]), .ZN(n101) );
  NAND2_X1 U186 ( .A1(rdata_L0[45]), .A2(n744), .ZN(n100) );
  AOI22_X1 U187 ( .A1(rdata_L0[13]), .A2(n892), .B1(rdata_last_q[13]), .B2(
        n871), .ZN(n99) );
  OAI211_X1 U188 ( .C1(n101), .C2(n777), .A(n100), .B(n99), .ZN(n730) );
  AOI22_X1 U189 ( .A1(n730), .A2(n537), .B1(rdata_L0[108]), .B2(n32), .ZN(n102) );
  OAI21_X1 U190 ( .B1(n884), .B2(n537), .A(n102), .ZN(rdata_o[13]) );
  INV_X1 U191 ( .A(fetch_gnt), .ZN(n357) );
  NAND2_X1 U192 ( .A1(n521), .A2(CS[1]), .ZN(n175) );
  NAND2_X1 U193 ( .A1(n521), .A2(n339), .ZN(n352) );
  NOR2_X1 U194 ( .A1(n352), .A2(CS[3]), .ZN(n382) );
  INV_X1 U195 ( .A(hwloop_i), .ZN(n380) );
  NAND2_X1 U196 ( .A1(n382), .A2(n380), .ZN(n151) );
  OAI21_X1 U197 ( .B1(n342), .B2(n175), .A(n151), .ZN(n128) );
  AOI22_X1 U198 ( .A1(n774), .A2(rdata_L0[0]), .B1(rdata_L0[64]), .B2(n756), 
        .ZN(n106) );
  NAND2_X1 U199 ( .A1(rdata_L0[32]), .A2(n744), .ZN(n104) );
  NAND4_X1 U200 ( .A1(n106), .A2(n105), .A3(n104), .A4(n103), .ZN(n186) );
  AOI22_X1 U201 ( .A1(n863), .A2(n755), .B1(rdata_last_q[1]), .B2(n871), .ZN(
        n110) );
  NAND2_X1 U202 ( .A1(rdata_L0[1]), .A2(n774), .ZN(n109) );
  NAND2_X1 U203 ( .A1(rdata_L0[65]), .A2(n756), .ZN(n108) );
  NAND2_X1 U204 ( .A1(rdata_L0[33]), .A2(n744), .ZN(n107) );
  NAND4_X1 U205 ( .A1(n110), .A2(n109), .A3(n108), .A4(n107), .ZN(n189) );
  NAND2_X1 U206 ( .A1(n186), .A2(n189), .ZN(n111) );
  NAND2_X1 U207 ( .A1(n111), .A2(n827), .ZN(n322) );
  NAND2_X1 U208 ( .A1(n322), .A2(addr_o[2]), .ZN(n122) );
  NAND2_X1 U209 ( .A1(rdata_L0[48]), .A2(n744), .ZN(n115) );
  NAND2_X1 U210 ( .A1(rdata_L0[80]), .A2(n756), .ZN(n114) );
  AOI22_X1 U211 ( .A1(n893), .A2(n755), .B1(rdata_last_q[16]), .B2(n871), .ZN(
        n113) );
  NAND2_X1 U212 ( .A1(rdata_L0[16]), .A2(n774), .ZN(n112) );
  NAND4_X1 U213 ( .A1(n115), .A2(n114), .A3(n113), .A4(n112), .ZN(n185) );
  NAND2_X1 U214 ( .A1(n855), .A2(n756), .ZN(n120) );
  AOI21_X1 U215 ( .B1(n41), .B2(n755), .A(n116), .ZN(n119) );
  NAND2_X1 U216 ( .A1(rdata_L0[17]), .A2(n774), .ZN(n118) );
  NAND2_X1 U217 ( .A1(rdata_L0[49]), .A2(n744), .ZN(n117) );
  NAND4_X1 U218 ( .A1(n120), .A2(n119), .A3(n118), .A4(n117), .ZN(n334) );
  NAND3_X1 U219 ( .A1(n185), .A2(addr_o[1]), .A3(n334), .ZN(n321) );
  AOI21_X1 U220 ( .B1(n321), .B2(n826), .A(n60), .ZN(n121) );
  NAND2_X1 U221 ( .A1(n122), .A2(n121), .ZN(n358) );
  NAND2_X1 U222 ( .A1(n176), .A2(n123), .ZN(n127) );
  AND2_X1 U223 ( .A1(n125), .A2(n124), .ZN(n126) );
  NAND2_X1 U224 ( .A1(n127), .A2(n126), .ZN(n343) );
  NAND2_X1 U225 ( .A1(n128), .A2(n343), .ZN(n405) );
  INV_X1 U226 ( .A(n405), .ZN(n132) );
  NAND2_X1 U227 ( .A1(fetch_valid), .A2(n339), .ZN(n362) );
  NOR2_X1 U228 ( .A1(n521), .A2(n362), .ZN(n344) );
  NAND2_X1 U229 ( .A1(n344), .A2(n787), .ZN(n387) );
  INV_X1 U230 ( .A(n387), .ZN(n129) );
  INV_X1 U231 ( .A(n35), .ZN(n388) );
  AND2_X1 U232 ( .A1(n129), .A2(n388), .ZN(n179) );
  NAND2_X1 U233 ( .A1(n130), .A2(n158), .ZN(n131) );
  NOR4_X1 U234 ( .A1(n132), .A2(n171), .A3(n179), .A4(n131), .ZN(n147) );
  NOR2_X1 U235 ( .A1(n392), .A2(CS[0]), .ZN(n399) );
  NAND2_X1 U236 ( .A1(fetch_valid), .A2(n399), .ZN(n513) );
  INV_X1 U237 ( .A(n513), .ZN(n139) );
  NAND2_X1 U238 ( .A1(n521), .A2(n176), .ZN(n384) );
  INV_X1 U240 ( .A(fetch_valid), .ZN(n400) );
  AOI21_X1 U241 ( .B1(n176), .B2(n400), .A(n43), .ZN(n134) );
  INV_X1 U242 ( .A(n399), .ZN(n133) );
  NOR3_X1 U243 ( .A1(n888), .A2(n134), .A3(n133), .ZN(n138) );
  AOI211_X1 U244 ( .C1(n339), .C2(n400), .A(n345), .B(n888), .ZN(n136) );
  NAND2_X1 U245 ( .A1(n521), .A2(n358), .ZN(n340) );
  NAND2_X1 U246 ( .A1(n340), .A2(CS[2]), .ZN(n135) );
  AOI21_X1 U247 ( .B1(n136), .B2(n135), .A(n788), .ZN(n137) );
  AOI211_X1 U248 ( .C1(n139), .C2(n384), .A(n138), .B(n137), .ZN(n140) );
  NOR2_X1 U249 ( .A1(n140), .A2(n787), .ZN(n145) );
  NAND2_X1 U250 ( .A1(n888), .A2(n390), .ZN(n153) );
  OAI21_X1 U251 ( .B1(fetch_valid), .B2(n393), .A(n153), .ZN(n394) );
  INV_X1 U252 ( .A(n394), .ZN(n143) );
  INV_X1 U253 ( .A(n141), .ZN(n159) );
  NAND2_X1 U254 ( .A1(n888), .A2(n159), .ZN(n402) );
  NAND3_X1 U255 ( .A1(n888), .A2(n142), .A3(n400), .ZN(n366) );
  OAI211_X1 U256 ( .C1(n143), .C2(n788), .A(n402), .B(n366), .ZN(n144) );
  NAND2_X1 U257 ( .A1(n521), .A2(n171), .ZN(n156) );
  OAI21_X1 U258 ( .B1(n145), .B2(n144), .A(n156), .ZN(n146) );
  OAI211_X1 U259 ( .C1(n357), .C2(n147), .A(n172), .B(n146), .ZN(NS[0]) );
  AND2_X1 U260 ( .A1(n172), .A2(is_hwlp_q), .ZN(is_hwlp_o) );
  OAI21_X1 U261 ( .B1(fetch_gnt), .B2(n158), .A(n393), .ZN(n372) );
  AOI21_X1 U262 ( .B1(n793), .B2(n788), .A(CS[3]), .ZN(n148) );
  OAI21_X1 U263 ( .B1(n521), .B2(n149), .A(n148), .ZN(n150) );
  NOR2_X1 U264 ( .A1(n372), .A2(n150), .ZN(n522) );
  NAND2_X1 U265 ( .A1(n522), .A2(n151), .ZN(n324) );
  NAND2_X1 U266 ( .A1(n521), .A2(n322), .ZN(n155) );
  INV_X1 U267 ( .A(n155), .ZN(n152) );
  NAND2_X1 U268 ( .A1(n156), .A2(n172), .ZN(n520) );
  INV_X1 U269 ( .A(n520), .ZN(n514) );
  NAND3_X1 U270 ( .A1(n324), .A2(n152), .A3(n514), .ZN(n314) );
  INV_X1 U271 ( .A(n382), .ZN(n154) );
  OAI21_X1 U272 ( .B1(n154), .B2(n380), .A(n153), .ZN(n318) );
  AOI21_X1 U273 ( .B1(n324), .B2(n155), .A(n318), .ZN(n157) );
  OR2_X1 U275 ( .A1(n156), .A2(n320), .ZN(n160) );
  OR2_X1 U276 ( .A1(fetch_gnt), .A2(n160), .ZN(n378) );
  OAI21_X1 U277 ( .B1(n157), .B2(n520), .A(n378), .ZN(n310) );
  NAND2_X1 U278 ( .A1(n310), .A2(addr_o[2]), .ZN(n165) );
  NAND3_X1 U279 ( .A1(n521), .A2(n390), .A3(n787), .ZN(n349) );
  OAI21_X1 U280 ( .B1(n357), .B2(n158), .A(n349), .ZN(n516) );
  AND2_X1 U281 ( .A1(n521), .A2(n159), .ZN(n397) );
  NOR2_X1 U282 ( .A1(n516), .A2(n397), .ZN(n162) );
  INV_X1 U283 ( .A(n160), .ZN(n161) );
  NAND2_X1 U284 ( .A1(fetch_gnt), .A2(n161), .ZN(n517) );
  OAI21_X1 U285 ( .B1(n162), .B2(n520), .A(n517), .ZN(n163) );
  INV_X1 U286 ( .A(n163), .ZN(n330) );
  INV_X1 U287 ( .A(n330), .ZN(n237) );
  AOI22_X1 U288 ( .A1(n237), .A2(hwloop_target_i[2]), .B1(addr_i[2]), .B2(n320), .ZN(n164) );
  OAI211_X1 U289 ( .C1(addr_o[2]), .C2(n314), .A(n165), .B(n164), .ZN(
        addr_n[2]) );
  INV_X1 U290 ( .A(n185), .ZN(n170) );
  AOI22_X1 U291 ( .A1(rdata_L0[32]), .A2(n762), .B1(n890), .B2(n42), .ZN(n169)
         );
  AOI22_X1 U292 ( .A1(rdata_L0[0]), .A2(n31), .B1(rdata_L0[64]), .B2(n34), 
        .ZN(n168) );
  OAI211_X1 U293 ( .C1(n170), .C2(n765), .A(n169), .B(n168), .ZN(rdata_o[16])
         );
  NAND2_X1 U294 ( .A1(fetch_gnt), .A2(n171), .ZN(n353) );
  OR2_X1 U296 ( .A1(n521), .A2(n320), .ZN(n173) );
  AOI21_X1 U299 ( .B1(n343), .B2(n174), .A(hwloop_i), .ZN(n364) );
  NAND2_X1 U300 ( .A1(n382), .A2(n364), .ZN(n178) );
  OAI21_X1 U301 ( .B1(n175), .B2(n43), .A(n383), .ZN(n348) );
  INV_X1 U302 ( .A(n176), .ZN(n389) );
  NAND2_X1 U303 ( .A1(n389), .A2(n383), .ZN(n177) );
  NAND4_X1 U304 ( .A1(n178), .A2(n387), .A3(n348), .A4(n177), .ZN(n180) );
  OR2_X1 U306 ( .A1(n182), .A2(n521), .ZN(n181) );
  MUX2_X1 U313 ( .A(n185), .B(n186), .S(n537), .Z(rdata_o[0]) );
  AOI22_X1 U314 ( .A1(n768), .A2(n186), .B1(rdata_last_q[0]), .B2(n1042), .ZN(
        n188) );
  AOI22_X1 U315 ( .A1(n770), .A2(n890), .B1(n12), .B2(rdata_o[0]), .ZN(n187)
         );
  NAND2_X1 U316 ( .A1(n188), .A2(n187), .ZN(n823) );
  MUX2_X1 U317 ( .A(n189), .B(n334), .S(n765), .Z(rdata_o[1]) );
  AOI22_X1 U318 ( .A1(n768), .A2(n189), .B1(rdata_last_q[1]), .B2(n1042), .ZN(
        n191) );
  AOI22_X1 U319 ( .A1(n770), .A2(n863), .B1(n12), .B2(rdata_o[1]), .ZN(n190)
         );
  NAND2_X1 U320 ( .A1(n191), .A2(n190), .ZN(n824) );
  AOI22_X1 U321 ( .A1(n237), .A2(hwloop_target_i[31]), .B1(n192), .B2(n320), 
        .ZN(n201) );
  NAND2_X1 U322 ( .A1(addr_o[18]), .A2(addr_o[19]), .ZN(n460) );
  NAND2_X1 U323 ( .A1(addr_o[20]), .A2(addr_o[21]), .ZN(n471) );
  NOR2_X1 U324 ( .A1(n460), .A2(n471), .ZN(n232) );
  NAND2_X1 U325 ( .A1(n232), .A2(addr_o[22]), .ZN(n227) );
  NOR2_X1 U326 ( .A1(n227), .A2(n38), .ZN(n198) );
  NAND2_X1 U327 ( .A1(addr_o[10]), .A2(addr_o[11]), .ZN(n428) );
  NAND2_X1 U328 ( .A1(addr_o[13]), .A2(addr_o[12]), .ZN(n443) );
  NOR2_X1 U329 ( .A1(n428), .A2(n443), .ZN(n255) );
  NAND2_X1 U330 ( .A1(addr_o[14]), .A2(addr_o[15]), .ZN(n444) );
  NAND2_X1 U331 ( .A1(addr_o[16]), .A2(addr_o[17]), .ZN(n461) );
  NOR2_X1 U332 ( .A1(n444), .A2(n461), .ZN(n193) );
  NAND2_X1 U333 ( .A1(n255), .A2(n193), .ZN(n197) );
  NAND2_X1 U334 ( .A1(addr_o[8]), .A2(addr_o[9]), .ZN(n429) );
  NOR2_X1 U335 ( .A1(n194), .A2(n429), .ZN(n196) );
  NAND2_X1 U336 ( .A1(n196), .A2(n195), .ZN(n254) );
  NOR2_X1 U337 ( .A1(n197), .A2(n254), .ZN(n226) );
  AND2_X1 U338 ( .A1(n198), .A2(n226), .ZN(n223) );
  XOR2_X1 U339 ( .A(n199), .B(addr_o[31]), .Z(n503) );
  NAND2_X1 U340 ( .A1(n265), .A2(n503), .ZN(n200) );
  OAI211_X1 U341 ( .C1(n264), .C2(n853), .A(n201), .B(n200), .ZN(addr_n[31])
         );
  AOI22_X1 U342 ( .A1(n237), .A2(hwloop_target_i[30]), .B1(addr_i[30]), .B2(
        n320), .ZN(n205) );
  HA_X1 U343 ( .A(n203), .B(addr_o[30]), .CO(n199), .S(n502) );
  NAND2_X1 U344 ( .A1(n265), .A2(n502), .ZN(n204) );
  OAI211_X1 U345 ( .C1(n264), .C2(n846), .A(n205), .B(n204), .ZN(addr_n[30])
         );
  AOI22_X1 U346 ( .A1(n237), .A2(hwloop_target_i[29]), .B1(addr_i[29]), .B2(
        n320), .ZN(n208) );
  HA_X1 U347 ( .A(n206), .B(addr_o[29]), .CO(n203), .S(n499) );
  NAND2_X1 U348 ( .A1(n265), .A2(n499), .ZN(n207) );
  OAI211_X1 U349 ( .C1(n264), .C2(n843), .A(n208), .B(n207), .ZN(addr_n[29])
         );
  AOI22_X1 U350 ( .A1(n237), .A2(hwloop_target_i[28]), .B1(n209), .B2(n320), 
        .ZN(n212) );
  HA_X1 U351 ( .A(n210), .B(addr_o[28]), .CO(n206), .S(n496) );
  NAND2_X1 U352 ( .A1(n265), .A2(n496), .ZN(n211) );
  OAI211_X1 U353 ( .C1(n264), .C2(n845), .A(n212), .B(n211), .ZN(addr_n[28])
         );
  AOI22_X1 U354 ( .A1(n237), .A2(hwloop_target_i[27]), .B1(addr_i[27]), .B2(
        n320), .ZN(n215) );
  HA_X1 U355 ( .A(n213), .B(addr_o[27]), .CO(n210), .S(n493) );
  NAND2_X1 U356 ( .A1(n265), .A2(n493), .ZN(n214) );
  OAI211_X1 U357 ( .C1(n264), .C2(n850), .A(n215), .B(n214), .ZN(addr_n[27])
         );
  AOI22_X1 U358 ( .A1(n237), .A2(hwloop_target_i[26]), .B1(n216), .B2(n320), 
        .ZN(n219) );
  HA_X1 U359 ( .A(n217), .B(addr_o[26]), .CO(n213), .S(n490) );
  NAND2_X1 U360 ( .A1(n265), .A2(n490), .ZN(n218) );
  OAI211_X1 U361 ( .C1(n264), .C2(n851), .A(n219), .B(n218), .ZN(addr_n[26])
         );
  AOI22_X1 U362 ( .A1(n237), .A2(hwloop_target_i[25]), .B1(n40), .B2(n320), 
        .ZN(n222) );
  HA_X1 U363 ( .A(n220), .B(addr_o[25]), .CO(n217), .S(n487) );
  NAND2_X1 U364 ( .A1(n265), .A2(n487), .ZN(n221) );
  OAI211_X1 U365 ( .C1(n264), .C2(n791), .A(n222), .B(n221), .ZN(addr_n[25])
         );
  AOI22_X1 U366 ( .A1(n237), .A2(hwloop_target_i[24]), .B1(n889), .B2(n320), 
        .ZN(n225) );
  HA_X1 U367 ( .A(n223), .B(addr_o[24]), .CO(n220), .S(n484) );
  NAND2_X1 U368 ( .A1(n265), .A2(n484), .ZN(n224) );
  OAI211_X1 U369 ( .C1(n264), .C2(n790), .A(n225), .B(n224), .ZN(addr_n[24])
         );
  AOI22_X1 U370 ( .A1(n237), .A2(hwloop_target_i[23]), .B1(n891), .B2(n320), 
        .ZN(n230) );
  INV_X1 U371 ( .A(n226), .ZN(n250) );
  NOR2_X1 U372 ( .A1(n250), .A2(n227), .ZN(n228) );
  XNOR2_X1 U373 ( .A(n228), .B(n38), .ZN(n479) );
  NAND2_X1 U374 ( .A1(n265), .A2(n479), .ZN(n229) );
  OAI211_X1 U375 ( .C1(n264), .C2(n38), .A(n230), .B(n229), .ZN(addr_n[23]) );
  AOI22_X1 U376 ( .A1(n237), .A2(hwloop_target_i[22]), .B1(n231), .B2(n320), 
        .ZN(n236) );
  INV_X1 U377 ( .A(n232), .ZN(n233) );
  NOR2_X1 U378 ( .A1(n250), .A2(n233), .ZN(n234) );
  XNOR2_X1 U379 ( .A(n234), .B(n838), .ZN(n474) );
  NAND2_X1 U380 ( .A1(n265), .A2(n474), .ZN(n235) );
  OAI211_X1 U381 ( .C1(n264), .C2(n838), .A(n236), .B(n235), .ZN(addr_n[22])
         );
  AOI22_X1 U382 ( .A1(n237), .A2(hwloop_target_i[21]), .B1(addr_i[21]), .B2(
        n320), .ZN(n240) );
  NOR2_X1 U383 ( .A1(n250), .A2(n460), .ZN(n242) );
  NAND2_X1 U384 ( .A1(n242), .A2(addr_o[20]), .ZN(n238) );
  XOR2_X1 U385 ( .A(n238), .B(n852), .Z(n470) );
  NAND2_X1 U386 ( .A1(n265), .A2(n470), .ZN(n239) );
  OAI211_X1 U387 ( .C1(n264), .C2(n852), .A(n240), .B(n239), .ZN(addr_n[21])
         );
  INV_X1 U388 ( .A(n330), .ZN(n290) );
  AOI22_X1 U389 ( .A1(n290), .A2(hwloop_target_i[20]), .B1(n241), .B2(n320), 
        .ZN(n244) );
  XNOR2_X1 U390 ( .A(n242), .B(n789), .ZN(n467) );
  NAND2_X1 U391 ( .A1(n265), .A2(n467), .ZN(n243) );
  OAI211_X1 U392 ( .C1(n264), .C2(n789), .A(n244), .B(n243), .ZN(addr_n[20])
         );
  AOI22_X1 U393 ( .A1(n290), .A2(hwloop_target_i[19]), .B1(n245), .B2(n320), 
        .ZN(n248) );
  NOR2_X1 U394 ( .A1(n250), .A2(n841), .ZN(n246) );
  XNOR2_X1 U395 ( .A(n246), .B(n837), .ZN(n459) );
  NAND2_X1 U396 ( .A1(n265), .A2(n459), .ZN(n247) );
  OAI211_X1 U397 ( .C1(n264), .C2(n837), .A(n248), .B(n247), .ZN(addr_n[19])
         );
  AOI22_X1 U398 ( .A1(n290), .A2(hwloop_target_i[18]), .B1(addr_i[18]), .B2(
        n320), .ZN(n252) );
  XOR2_X1 U399 ( .A(n250), .B(n841), .Z(n455) );
  NAND2_X1 U400 ( .A1(n265), .A2(n455), .ZN(n251) );
  OAI211_X1 U401 ( .C1(n264), .C2(n841), .A(n252), .B(n251), .ZN(addr_n[18])
         );
  AOI22_X1 U402 ( .A1(n290), .A2(hwloop_target_i[17]), .B1(n253), .B2(n320), 
        .ZN(n259) );
  INV_X1 U403 ( .A(n254), .ZN(n286) );
  NAND2_X1 U404 ( .A1(n286), .A2(n255), .ZN(n266) );
  INV_X1 U405 ( .A(n266), .ZN(n271) );
  INV_X1 U406 ( .A(n444), .ZN(n256) );
  NAND2_X1 U407 ( .A1(n271), .A2(n256), .ZN(n261) );
  NOR2_X1 U408 ( .A1(n261), .A2(n842), .ZN(n257) );
  XNOR2_X1 U409 ( .A(n257), .B(n840), .ZN(n451) );
  NAND2_X1 U410 ( .A1(n265), .A2(n451), .ZN(n258) );
  OAI211_X1 U411 ( .C1(n264), .C2(n840), .A(n259), .B(n258), .ZN(addr_n[17])
         );
  AOI22_X1 U412 ( .A1(n290), .A2(hwloop_target_i[16]), .B1(n260), .B2(n320), 
        .ZN(n263) );
  XOR2_X1 U413 ( .A(n261), .B(n842), .Z(n447) );
  NAND2_X1 U414 ( .A1(n265), .A2(n447), .ZN(n262) );
  OAI211_X1 U415 ( .C1(n264), .C2(n842), .A(n263), .B(n262), .ZN(addr_n[16])
         );
  AOI22_X1 U416 ( .A1(n290), .A2(hwloop_target_i[15]), .B1(addr_i[15]), .B2(
        n320), .ZN(n269) );
  NOR2_X1 U417 ( .A1(n266), .A2(n849), .ZN(n267) );
  XNOR2_X1 U418 ( .A(n267), .B(n835), .ZN(n442) );
  NAND2_X1 U419 ( .A1(n265), .A2(n442), .ZN(n268) );
  OAI211_X1 U420 ( .C1(n264), .C2(n835), .A(n269), .B(n268), .ZN(addr_n[15])
         );
  AOI22_X1 U421 ( .A1(n290), .A2(hwloop_target_i[14]), .B1(n270), .B2(n320), 
        .ZN(n273) );
  XNOR2_X1 U422 ( .A(n271), .B(n849), .ZN(n438) );
  NAND2_X1 U423 ( .A1(n265), .A2(n438), .ZN(n272) );
  OAI211_X1 U424 ( .C1(n264), .C2(n849), .A(n273), .B(n272), .ZN(addr_n[14])
         );
  AOI22_X1 U425 ( .A1(n290), .A2(hwloop_target_i[13]), .B1(addr_i[13]), .B2(
        n320), .ZN(n277) );
  INV_X1 U426 ( .A(n428), .ZN(n274) );
  NAND2_X1 U427 ( .A1(n286), .A2(n274), .ZN(n278) );
  NOR2_X1 U428 ( .A1(n278), .A2(n834), .ZN(n275) );
  XNOR2_X1 U429 ( .A(n275), .B(n836), .ZN(n435) );
  NAND2_X1 U430 ( .A1(n265), .A2(n435), .ZN(n276) );
  OAI211_X1 U431 ( .C1(n264), .C2(n836), .A(n277), .B(n276), .ZN(addr_n[13])
         );
  AOI22_X1 U432 ( .A1(n290), .A2(hwloop_target_i[12]), .B1(addr_i[12]), .B2(
        n320), .ZN(n280) );
  XOR2_X1 U433 ( .A(n278), .B(n834), .Z(n432) );
  NAND2_X1 U434 ( .A1(n265), .A2(n432), .ZN(n279) );
  OAI211_X1 U435 ( .C1(n264), .C2(n834), .A(n280), .B(n279), .ZN(addr_n[12])
         );
  AOI22_X1 U436 ( .A1(n290), .A2(hwloop_target_i[11]), .B1(addr_i[11]), .B2(
        n320), .ZN(n283) );
  NAND2_X1 U437 ( .A1(n286), .A2(addr_o[10]), .ZN(n281) );
  XOR2_X1 U438 ( .A(n281), .B(n839), .Z(n427) );
  NAND2_X1 U439 ( .A1(n265), .A2(n427), .ZN(n282) );
  OAI211_X1 U440 ( .C1(n264), .C2(n839), .A(n283), .B(n282), .ZN(addr_n[11])
         );
  AOI22_X1 U441 ( .A1(n290), .A2(hwloop_target_i[10]), .B1(n285), .B2(n320), 
        .ZN(n288) );
  XNOR2_X1 U442 ( .A(n286), .B(n831), .ZN(n423) );
  NAND2_X1 U443 ( .A1(n265), .A2(n423), .ZN(n287) );
  OAI211_X1 U444 ( .C1(n264), .C2(n831), .A(n288), .B(n287), .ZN(addr_n[10])
         );
  AOI22_X1 U445 ( .A1(n290), .A2(hwloop_target_i[9]), .B1(n289), .B2(n320), 
        .ZN(n294) );
  NAND2_X1 U446 ( .A1(n291), .A2(addr_o[8]), .ZN(n292) );
  XOR2_X1 U447 ( .A(n292), .B(n844), .Z(n421) );
  NAND2_X1 U448 ( .A1(n265), .A2(n421), .ZN(n293) );
  OAI211_X1 U449 ( .C1(n264), .C2(n844), .A(n294), .B(n293), .ZN(addr_n[9]) );
  INV_X1 U450 ( .A(n330), .ZN(n519) );
  AOI22_X1 U451 ( .A1(n519), .A2(hwloop_target_i[8]), .B1(n295), .B2(n320), 
        .ZN(n298) );
  NAND2_X1 U452 ( .A1(n265), .A2(n296), .ZN(n297) );
  OAI211_X1 U453 ( .C1(n264), .C2(n832), .A(n298), .B(n297), .ZN(addr_n[8]) );
  AOI22_X1 U454 ( .A1(n519), .A2(hwloop_target_i[7]), .B1(addr_i[7]), .B2(n320), .ZN(n301) );
  NOR2_X1 U455 ( .A1(n302), .A2(n833), .ZN(n299) );
  XNOR2_X1 U456 ( .A(n299), .B(n847), .ZN(n419) );
  NAND2_X1 U457 ( .A1(n265), .A2(n419), .ZN(n300) );
  OAI211_X1 U458 ( .C1(n264), .C2(n847), .A(n301), .B(n300), .ZN(addr_n[7]) );
  AOI22_X1 U459 ( .A1(n519), .A2(hwloop_target_i[6]), .B1(addr_i[6]), .B2(n320), .ZN(n304) );
  XOR2_X1 U460 ( .A(n302), .B(n833), .Z(n415) );
  NAND2_X1 U461 ( .A1(n265), .A2(n415), .ZN(n303) );
  OAI211_X1 U462 ( .C1(n264), .C2(n833), .A(n304), .B(n303), .ZN(addr_n[6]) );
  AOI22_X1 U463 ( .A1(n519), .A2(hwloop_target_i[5]), .B1(addr_i[5]), .B2(n320), .ZN(n309) );
  NAND2_X1 U464 ( .A1(n123), .A2(addr_o[4]), .ZN(n307) );
  XOR2_X1 U465 ( .A(n307), .B(n848), .Z(n412) );
  NAND2_X1 U466 ( .A1(n265), .A2(n412), .ZN(n308) );
  OAI211_X1 U467 ( .C1(n264), .C2(n848), .A(n309), .B(n308), .ZN(addr_n[5]) );
  XNOR2_X1 U468 ( .A(n123), .B(n828), .ZN(n410) );
  INV_X1 U469 ( .A(n410), .ZN(n313) );
  NAND2_X1 U470 ( .A1(n310), .A2(addr_o[4]), .ZN(n312) );
  AOI22_X1 U471 ( .A1(n519), .A2(hwloop_target_i[4]), .B1(addr_i[4]), .B2(n320), .ZN(n311) );
  OAI211_X1 U472 ( .C1(n314), .C2(n313), .A(n312), .B(n311), .ZN(addr_n[4]) );
  AOI22_X1 U473 ( .A1(n519), .A2(hwloop_target_i[3]), .B1(addr_i[3]), .B2(n320), .ZN(n317) );
  NAND2_X1 U474 ( .A1(n265), .A2(n315), .ZN(n316) );
  OAI211_X1 U475 ( .C1(n264), .C2(n60), .A(n317), .B(n316), .ZN(addr_n[3]) );
  INV_X1 U476 ( .A(hwloop_target_i[1]), .ZN(n329) );
  INV_X1 U477 ( .A(n318), .ZN(n319) );
  OAI21_X1 U478 ( .B1(n319), .B2(n520), .A(n378), .ZN(n523) );
  AOI22_X1 U479 ( .A1(n523), .A2(addr_o[1]), .B1(n320), .B2(addr_i[1]), .ZN(
        n328) );
  INV_X1 U480 ( .A(n321), .ZN(n326) );
  INV_X1 U481 ( .A(n322), .ZN(n323) );
  MUX2_X1 U482 ( .A(addr_o[1]), .B(n323), .S(n521), .Z(n325) );
  OAI211_X1 U483 ( .C1(n326), .C2(n325), .A(n324), .B(n514), .ZN(n327) );
  OAI211_X1 U484 ( .C1(n330), .C2(n329), .A(n328), .B(n327), .ZN(addr_n[1]) );
  INV_X1 U485 ( .A(n334), .ZN(n333) );
  AOI22_X1 U486 ( .A1(rdata_L0[33]), .A2(n762), .B1(n863), .B2(n42), .ZN(n332)
         );
  AOI22_X1 U487 ( .A1(rdata_L0[1]), .A2(n31), .B1(rdata_L0[65]), .B2(n34), 
        .ZN(n331) );
  OAI211_X1 U488 ( .C1(n333), .C2(n765), .A(n332), .B(n331), .ZN(rdata_o[17])
         );
  INV_X1 U492 ( .A(n337), .ZN(n338) );
  NOR4_X1 U493 ( .A1(n340), .A2(n345), .A3(n339), .A4(n338), .ZN(n341) );
  OAI21_X1 U494 ( .B1(n343), .B2(n342), .A(n341), .ZN(n351) );
  INV_X1 U495 ( .A(n344), .ZN(n367) );
  NAND2_X1 U496 ( .A1(n346), .A2(n345), .ZN(n347) );
  NAND4_X1 U497 ( .A1(n348), .A2(n367), .A3(n513), .A4(n347), .ZN(n350) );
  NAND2_X1 U498 ( .A1(n397), .A2(fetch_valid), .ZN(n512) );
  NAND2_X1 U499 ( .A1(n512), .A2(n349), .ZN(n373) );
  AOI211_X1 U500 ( .C1(CS[3]), .C2(n351), .A(n350), .B(n373), .ZN(n355) );
  INV_X1 U501 ( .A(n352), .ZN(n371) );
  NAND2_X1 U502 ( .A1(n371), .A2(n364), .ZN(n354) );
  NAND2_X1 U503 ( .A1(n353), .A2(n514), .ZN(n409) );
  AOI21_X1 U504 ( .B1(n355), .B2(n354), .A(n409), .ZN(NS[3]) );
  AOI21_X1 U505 ( .B1(fetch_gnt), .B2(n384), .A(n43), .ZN(n356) );
  AOI211_X1 U506 ( .C1(n357), .C2(n888), .A(CS[0]), .B(n356), .ZN(n363) );
  OAI21_X1 U507 ( .B1(n389), .B2(n788), .A(n359), .ZN(n360) );
  NAND3_X1 U508 ( .A1(n521), .A2(CS[2]), .A3(n360), .ZN(n361) );
  OAI211_X1 U509 ( .C1(n363), .C2(n793), .A(n362), .B(n361), .ZN(n377) );
  OAI21_X1 U510 ( .B1(fetch_gnt), .B2(n43), .A(n364), .ZN(n370) );
  OAI22_X1 U511 ( .A1(n366), .A2(n793), .B1(n365), .B2(n513), .ZN(n369) );
  NOR3_X1 U512 ( .A1(fetch_gnt), .A2(n388), .A3(n367), .ZN(n368) );
  AOI211_X1 U513 ( .C1(n371), .C2(n370), .A(n369), .B(n368), .ZN(n375) );
  AOI21_X1 U514 ( .B1(n373), .B2(n36), .A(n372), .ZN(n374) );
  OAI21_X1 U515 ( .B1(n375), .B2(CS[3]), .A(n374), .ZN(n376) );
  AOI21_X1 U516 ( .B1(CS[3]), .B2(n377), .A(n376), .ZN(n379) );
  OAI211_X1 U517 ( .C1(n379), .C2(n520), .A(n378), .B(n594), .ZN(NS[1]) );
  NAND3_X1 U518 ( .A1(n382), .A2(n174), .A3(n380), .ZN(n386) );
  NAND3_X1 U519 ( .A1(n384), .A2(CS[1]), .A3(n383), .ZN(n385) );
  OAI211_X1 U520 ( .C1(n388), .C2(n387), .A(n386), .B(n385), .ZN(n407) );
  OAI21_X1 U521 ( .B1(n390), .B2(n399), .A(n389), .ZN(n391) );
  OAI211_X1 U522 ( .C1(n521), .C2(n392), .A(n391), .B(n393), .ZN(n396) );
  NOR2_X1 U523 ( .A1(n393), .A2(CS[0]), .ZN(n395) );
  AOI211_X1 U524 ( .C1(CS[3]), .C2(n396), .A(n395), .B(n394), .ZN(n404) );
  NAND2_X1 U525 ( .A1(n43), .A2(CS[3]), .ZN(n398) );
  AOI21_X1 U526 ( .B1(n399), .B2(n398), .A(n397), .ZN(n401) );
  MUX2_X1 U527 ( .A(n402), .B(n401), .S(n400), .Z(n403) );
  OAI211_X1 U528 ( .C1(n405), .C2(n43), .A(n404), .B(n403), .ZN(n406) );
  AOI21_X1 U529 ( .B1(fetch_gnt), .B2(n407), .A(n406), .ZN(n408) );
  NOR2_X1 U530 ( .A1(n409), .A2(n408), .ZN(NS[2]) );
  XNOR2_X1 U531 ( .A(n848), .B(addr_o[4]), .ZN(n411) );
  INV_X1 U532 ( .A(n413), .ZN(n416) );
  XNOR2_X1 U533 ( .A(n833), .B(n416), .ZN(n414) );
  MUX2_X1 U534 ( .A(n415), .B(n414), .S(n30), .Z(addr_real_next[6]) );
  NAND2_X1 U535 ( .A1(n416), .A2(addr_o[6]), .ZN(n417) );
  XOR2_X1 U536 ( .A(n417), .B(n847), .Z(n418) );
  NOR2_X1 U537 ( .A1(n422), .A2(n832), .ZN(n420) );
  NOR2_X1 U538 ( .A1(n422), .A2(n429), .ZN(n424) );
  NAND2_X1 U539 ( .A1(n424), .A2(addr_o[10]), .ZN(n425) );
  XOR2_X1 U540 ( .A(n425), .B(n839), .Z(n426) );
  MUX2_X1 U541 ( .A(n427), .B(n426), .S(n509), .Z(addr_real_next[11]) );
  NOR2_X1 U542 ( .A1(n429), .A2(n428), .ZN(n431) );
  NAND2_X1 U543 ( .A1(n431), .A2(n430), .ZN(n464) );
  INV_X1 U544 ( .A(n464), .ZN(n445) );
  NAND2_X1 U545 ( .A1(n445), .A2(addr_o[12]), .ZN(n433) );
  XOR2_X1 U546 ( .A(n433), .B(n836), .Z(n434) );
  MUX2_X1 U547 ( .A(n435), .B(n434), .S(n854), .Z(addr_real_next[13]) );
  INV_X1 U548 ( .A(n443), .ZN(n436) );
  NAND2_X1 U549 ( .A1(n445), .A2(n436), .ZN(n439) );
  XOR2_X1 U550 ( .A(n439), .B(n849), .Z(n437) );
  NOR2_X1 U551 ( .A1(n439), .A2(n849), .ZN(n440) );
  XNOR2_X1 U552 ( .A(n440), .B(n835), .ZN(n441) );
  MUX2_X1 U553 ( .A(n442), .B(n441), .S(n854), .Z(addr_real_next[15]) );
  NOR2_X1 U554 ( .A1(n444), .A2(n443), .ZN(n463) );
  NAND2_X1 U555 ( .A1(n445), .A2(n463), .ZN(n448) );
  INV_X1 U556 ( .A(n448), .ZN(n453) );
  XNOR2_X1 U557 ( .A(n453), .B(n842), .ZN(n446) );
  MUX2_X1 U558 ( .A(n447), .B(n446), .S(n7), .Z(addr_real_next[16]) );
  NOR2_X1 U559 ( .A1(n448), .A2(n842), .ZN(n449) );
  XNOR2_X1 U560 ( .A(n449), .B(n840), .ZN(n450) );
  MUX2_X1 U561 ( .A(n451), .B(n450), .S(n7), .Z(addr_real_next[17]) );
  INV_X1 U562 ( .A(n461), .ZN(n452) );
  NAND2_X1 U563 ( .A1(n453), .A2(n452), .ZN(n456) );
  XOR2_X1 U564 ( .A(n456), .B(n841), .Z(n454) );
  NOR2_X1 U565 ( .A1(n456), .A2(n841), .ZN(n457) );
  XNOR2_X1 U566 ( .A(n457), .B(n837), .ZN(n458) );
  MUX2_X1 U567 ( .A(n459), .B(n458), .S(n509), .Z(addr_real_next[19]) );
  NOR2_X1 U568 ( .A1(n461), .A2(n460), .ZN(n462) );
  NAND2_X1 U569 ( .A1(n463), .A2(n462), .ZN(n465) );
  NOR2_X1 U570 ( .A1(n465), .A2(n464), .ZN(n482) );
  INV_X1 U571 ( .A(n482), .ZN(n476) );
  XOR2_X1 U572 ( .A(n476), .B(n789), .Z(n466) );
  MUX2_X1 U573 ( .A(n467), .B(n466), .S(n854), .Z(addr_real_next[20]) );
  NOR2_X1 U574 ( .A1(n476), .A2(n789), .ZN(n468) );
  XNOR2_X1 U575 ( .A(n468), .B(n852), .ZN(n469) );
  MUX2_X1 U576 ( .A(n470), .B(n469), .S(n509), .Z(addr_real_next[21]) );
  INV_X1 U577 ( .A(n471), .ZN(n475) );
  NOR2_X1 U578 ( .A1(n476), .A2(n471), .ZN(n472) );
  XNOR2_X1 U579 ( .A(n472), .B(n838), .ZN(n473) );
  MUX2_X1 U580 ( .A(n474), .B(n473), .S(n854), .Z(addr_real_next[22]) );
  NAND2_X1 U581 ( .A1(n475), .A2(addr_o[22]), .ZN(n480) );
  NOR2_X1 U582 ( .A1(n476), .A2(n480), .ZN(n477) );
  XNOR2_X1 U583 ( .A(n477), .B(n38), .ZN(n478) );
  NOR2_X1 U585 ( .A1(n480), .A2(n38), .ZN(n481) );
  AND2_X1 U586 ( .A1(n482), .A2(n481), .ZN(n485) );
  HA_X1 U587 ( .A(n485), .B(addr_o[24]), .CO(n488), .S(n483) );
  MUX2_X1 U588 ( .A(n487), .B(n486), .S(n509), .Z(addr_real_next[25]) );
  HA_X1 U589 ( .A(n488), .B(addr_o[25]), .CO(n491), .S(n486) );
  MUX2_X1 U590 ( .A(n490), .B(n489), .S(n30), .Z(addr_real_next[26]) );
  HA_X1 U591 ( .A(n491), .B(addr_o[26]), .CO(n494), .S(n489) );
  MUX2_X1 U592 ( .A(n493), .B(n492), .S(n509), .Z(addr_real_next[27]) );
  HA_X1 U593 ( .A(n494), .B(addr_o[27]), .CO(n497), .S(n492) );
  MUX2_X1 U594 ( .A(n496), .B(n495), .S(n7), .Z(addr_real_next[28]) );
  HA_X1 U595 ( .A(n497), .B(addr_o[28]), .CO(n500), .S(n495) );
  MUX2_X1 U596 ( .A(n499), .B(n498), .S(n509), .Z(addr_real_next[29]) );
  HA_X1 U597 ( .A(n500), .B(addr_o[29]), .CO(n504), .S(n498) );
  MUX2_X1 U598 ( .A(n502), .B(n501), .S(n30), .Z(addr_real_next[30]) );
  INV_X1 U599 ( .A(n503), .ZN(n508) );
  HA_X1 U600 ( .A(n504), .B(addr_o[30]), .CO(n505), .S(n501) );
  XOR2_X1 U601 ( .A(n505), .B(addr_o[31]), .Z(n506) );
  NAND2_X1 U602 ( .A1(n509), .A2(n506), .ZN(n507) );
  OAI21_X1 U603 ( .B1(n854), .B2(n508), .A(n507), .ZN(addr_real_next[31]) );
  NAND2_X1 U604 ( .A1(n888), .A2(is_hwlp_q), .ZN(n511) );
  OAI211_X1 U605 ( .C1(CS[3]), .C2(n513), .A(n512), .B(n511), .ZN(n515) );
  OAI21_X1 U606 ( .B1(n516), .B2(n515), .A(n514), .ZN(n518) );
  NAND2_X1 U607 ( .A1(n518), .A2(n517), .ZN(is_hwlp_n) );
  NAND2_X1 U608 ( .A1(n519), .A2(hwloop_target_i[0]), .ZN(n526) );
  NOR3_X1 U609 ( .A1(n522), .A2(n521), .A3(n520), .ZN(n524) );
  OAI21_X1 U610 ( .B1(n524), .B2(n523), .A(addr_o[0]), .ZN(n525) );
  NAND2_X1 U611 ( .A1(n526), .A2(n525), .ZN(addr_n[0]) );
  AOI22_X1 U612 ( .A1(rdata_L0[113]), .A2(n755), .B1(rdata_last_q[18]), .B2(
        n871), .ZN(n531) );
  NAND2_X1 U613 ( .A1(rdata_L0[18]), .A2(n774), .ZN(n530) );
  NAND2_X1 U614 ( .A1(rdata_L0[81]), .A2(n756), .ZN(n529) );
  NAND2_X1 U615 ( .A1(rdata_L0[50]), .A2(n744), .ZN(n528) );
  AOI22_X1 U618 ( .A1(rdata_L0[34]), .A2(n762), .B1(rdata_L0[97]), .B2(n42), 
        .ZN(n533) );
  AOI22_X1 U619 ( .A1(rdata_L0[2]), .A2(n31), .B1(rdata_L0[66]), .B2(n34), 
        .ZN(n532) );
  OAI211_X1 U620 ( .C1(n883), .C2(n765), .A(n533), .B(n532), .ZN(rdata_o[18])
         );
  INV_X1 U625 ( .A(rdata_L0[66]), .ZN(n541) );
  NAND2_X1 U626 ( .A1(rdata_L0[34]), .A2(n744), .ZN(n540) );
  AOI22_X1 U627 ( .A1(rdata_L0[2]), .A2(n892), .B1(rdata_last_q[2]), .B2(n871), 
        .ZN(n539) );
  OAI211_X1 U628 ( .C1(n541), .C2(n777), .A(n540), .B(n539), .ZN(n544) );
  AOI22_X1 U629 ( .A1(n544), .A2(n537), .B1(rdata_L0[97]), .B2(n32), .ZN(n542)
         );
  OAI21_X1 U630 ( .B1(n883), .B2(n537), .A(n542), .ZN(rdata_o[2]) );
  INV_X1 U631 ( .A(n544), .ZN(n550) );
  AOI21_X1 U633 ( .B1(n755), .B2(n545), .A(n770), .ZN(n546) );
  NAND2_X1 U634 ( .A1(n782), .A2(rdata_L0[97]), .ZN(n549) );
  AOI22_X1 U635 ( .A1(n1042), .A2(rdata_last_q[2]), .B1(n12), .B2(rdata_o[2]), 
        .ZN(n548) );
  OAI211_X1 U636 ( .C1(n550), .C2(n785), .A(n549), .B(n548), .ZN(n822) );
  AOI22_X1 U637 ( .A1(rdata_L0[114]), .A2(n755), .B1(rdata_last_q[19]), .B2(
        n871), .ZN(n554) );
  NAND2_X1 U638 ( .A1(rdata_L0[19]), .A2(n892), .ZN(n553) );
  NAND2_X1 U639 ( .A1(rdata_L0[82]), .A2(n756), .ZN(n552) );
  NAND2_X1 U640 ( .A1(rdata_L0[51]), .A2(n744), .ZN(n551) );
  AOI22_X1 U643 ( .A1(rdata_L0[35]), .A2(n762), .B1(rdata_L0[98]), .B2(n42), 
        .ZN(n556) );
  AOI22_X1 U644 ( .A1(rdata_L0[3]), .A2(n31), .B1(rdata_L0[67]), .B2(n34), 
        .ZN(n555) );
  OAI211_X1 U645 ( .C1(n882), .C2(n765), .A(n556), .B(n555), .ZN(rdata_o[19])
         );
  INV_X1 U649 ( .A(rdata_L0[67]), .ZN(n562) );
  NAND2_X1 U650 ( .A1(rdata_L0[35]), .A2(n744), .ZN(n561) );
  AOI22_X1 U651 ( .A1(rdata_L0[3]), .A2(n892), .B1(rdata_last_q[3]), .B2(n871), 
        .ZN(n560) );
  OAI211_X1 U652 ( .C1(n562), .C2(n777), .A(n561), .B(n560), .ZN(n565) );
  AOI22_X1 U653 ( .A1(n565), .A2(n537), .B1(rdata_L0[98]), .B2(n32), .ZN(n563)
         );
  OAI21_X1 U654 ( .B1(n882), .B2(n537), .A(n563), .ZN(rdata_o[3]) );
  INV_X1 U655 ( .A(n565), .ZN(n568) );
  NAND2_X1 U656 ( .A1(n782), .A2(rdata_L0[98]), .ZN(n567) );
  AOI22_X1 U657 ( .A1(n1042), .A2(rdata_last_q[3]), .B1(n12), .B2(rdata_o[3]), 
        .ZN(n566) );
  OAI211_X1 U658 ( .C1(n568), .C2(n785), .A(n567), .B(n566), .ZN(n821) );
  AOI22_X1 U659 ( .A1(rdata_L0[115]), .A2(n755), .B1(rdata_last_q[20]), .B2(
        n871), .ZN(n572) );
  NAND2_X1 U660 ( .A1(rdata_L0[20]), .A2(n774), .ZN(n571) );
  NAND2_X1 U661 ( .A1(rdata_L0[83]), .A2(n756), .ZN(n570) );
  NAND2_X1 U662 ( .A1(rdata_L0[52]), .A2(n744), .ZN(n569) );
  AOI22_X1 U665 ( .A1(rdata_L0[36]), .A2(n762), .B1(rdata_L0[99]), .B2(n42), 
        .ZN(n574) );
  AOI22_X1 U666 ( .A1(rdata_L0[4]), .A2(n31), .B1(rdata_L0[68]), .B2(n34), 
        .ZN(n573) );
  OAI211_X1 U667 ( .C1(n881), .C2(n765), .A(n574), .B(n573), .ZN(rdata_o[20])
         );
  INV_X1 U671 ( .A(rdata_L0[68]), .ZN(n580) );
  NAND2_X1 U672 ( .A1(rdata_L0[36]), .A2(n744), .ZN(n579) );
  AOI22_X1 U673 ( .A1(rdata_L0[4]), .A2(n892), .B1(rdata_last_q[4]), .B2(n871), 
        .ZN(n578) );
  OAI211_X1 U674 ( .C1(n580), .C2(n777), .A(n579), .B(n578), .ZN(n583) );
  AOI22_X1 U675 ( .A1(n583), .A2(n537), .B1(rdata_L0[99]), .B2(n32), .ZN(n581)
         );
  OAI21_X1 U676 ( .B1(n881), .B2(n537), .A(n581), .ZN(rdata_o[4]) );
  INV_X1 U677 ( .A(n583), .ZN(n586) );
  NAND2_X1 U678 ( .A1(n782), .A2(rdata_L0[99]), .ZN(n585) );
  AOI22_X1 U679 ( .A1(n1042), .A2(rdata_last_q[4]), .B1(n12), .B2(rdata_o[4]), 
        .ZN(n584) );
  OAI211_X1 U680 ( .C1(n586), .C2(n785), .A(n585), .B(n584), .ZN(n820) );
  AOI22_X1 U681 ( .A1(rdata_L0[116]), .A2(n755), .B1(rdata_last_q[21]), .B2(
        n871), .ZN(n590) );
  NAND2_X1 U682 ( .A1(rdata_L0[21]), .A2(n892), .ZN(n589) );
  NAND2_X1 U683 ( .A1(rdata_L0[84]), .A2(n756), .ZN(n588) );
  NAND2_X1 U684 ( .A1(rdata_L0[53]), .A2(n744), .ZN(n587) );
  AOI22_X1 U687 ( .A1(rdata_L0[37]), .A2(n762), .B1(rdata_L0[100]), .B2(n42), 
        .ZN(n592) );
  AOI22_X1 U688 ( .A1(rdata_L0[5]), .A2(n31), .B1(rdata_L0[69]), .B2(n34), 
        .ZN(n591) );
  OAI211_X1 U689 ( .C1(n880), .C2(n765), .A(n592), .B(n591), .ZN(rdata_o[21])
         );
  INV_X1 U693 ( .A(rdata_L0[69]), .ZN(n599) );
  NAND2_X1 U694 ( .A1(rdata_L0[37]), .A2(n744), .ZN(n598) );
  AOI22_X1 U695 ( .A1(rdata_L0[5]), .A2(n892), .B1(rdata_last_q[5]), .B2(n871), 
        .ZN(n597) );
  OAI211_X1 U696 ( .C1(n599), .C2(n777), .A(n598), .B(n597), .ZN(n602) );
  AOI22_X1 U697 ( .A1(n602), .A2(n537), .B1(rdata_L0[100]), .B2(n32), .ZN(n600) );
  OAI21_X1 U698 ( .B1(n880), .B2(n537), .A(n600), .ZN(rdata_o[5]) );
  INV_X1 U699 ( .A(n602), .ZN(n605) );
  NAND2_X1 U700 ( .A1(n782), .A2(rdata_L0[100]), .ZN(n604) );
  AOI22_X1 U701 ( .A1(n547), .A2(rdata_last_q[5]), .B1(n12), .B2(rdata_o[5]), 
        .ZN(n603) );
  OAI211_X1 U702 ( .C1(n605), .C2(n785), .A(n604), .B(n603), .ZN(n819) );
  AOI22_X1 U703 ( .A1(rdata_L0[117]), .A2(n755), .B1(rdata_last_q[22]), .B2(
        n871), .ZN(n609) );
  NAND2_X1 U704 ( .A1(rdata_L0[22]), .A2(n892), .ZN(n608) );
  NAND2_X1 U705 ( .A1(rdata_L0[85]), .A2(n756), .ZN(n607) );
  NAND2_X1 U706 ( .A1(rdata_L0[54]), .A2(n773), .ZN(n606) );
  AOI22_X1 U709 ( .A1(rdata_L0[38]), .A2(n762), .B1(rdata_L0[101]), .B2(n42), 
        .ZN(n611) );
  AOI22_X1 U710 ( .A1(rdata_L0[6]), .A2(n31), .B1(rdata_L0[70]), .B2(n34), 
        .ZN(n610) );
  OAI211_X1 U711 ( .C1(n879), .C2(n765), .A(n611), .B(n610), .ZN(rdata_o[22])
         );
  INV_X1 U715 ( .A(rdata_L0[70]), .ZN(n617) );
  NAND2_X1 U716 ( .A1(rdata_L0[38]), .A2(n773), .ZN(n616) );
  AOI22_X1 U717 ( .A1(rdata_L0[6]), .A2(n892), .B1(rdata_last_q[6]), .B2(n871), 
        .ZN(n615) );
  OAI211_X1 U718 ( .C1(n617), .C2(n777), .A(n616), .B(n615), .ZN(n620) );
  AOI22_X1 U719 ( .A1(n620), .A2(n537), .B1(rdata_L0[101]), .B2(n32), .ZN(n618) );
  OAI21_X1 U720 ( .B1(n879), .B2(n537), .A(n618), .ZN(rdata_o[6]) );
  INV_X1 U721 ( .A(n620), .ZN(n623) );
  NAND2_X1 U722 ( .A1(n782), .A2(rdata_L0[101]), .ZN(n622) );
  AOI22_X1 U723 ( .A1(n547), .A2(rdata_last_q[6]), .B1(n12), .B2(rdata_o[6]), 
        .ZN(n621) );
  OAI211_X1 U724 ( .C1(n623), .C2(n785), .A(n622), .B(n621), .ZN(n818) );
  AOI22_X1 U725 ( .A1(rdata_L0[118]), .A2(n755), .B1(rdata_last_q[23]), .B2(
        n871), .ZN(n627) );
  NAND2_X1 U726 ( .A1(rdata_L0[23]), .A2(n892), .ZN(n626) );
  NAND2_X1 U727 ( .A1(rdata_L0[86]), .A2(n756), .ZN(n625) );
  NAND2_X1 U728 ( .A1(rdata_L0[55]), .A2(n744), .ZN(n624) );
  AOI22_X1 U731 ( .A1(rdata_L0[39]), .A2(n762), .B1(rdata_L0[102]), .B2(n42), 
        .ZN(n629) );
  AOI22_X1 U732 ( .A1(rdata_L0[7]), .A2(n31), .B1(rdata_L0[71]), .B2(n34), 
        .ZN(n628) );
  OAI211_X1 U733 ( .C1(n878), .C2(n765), .A(n629), .B(n628), .ZN(rdata_o[23])
         );
  INV_X1 U737 ( .A(rdata_L0[71]), .ZN(n635) );
  NAND2_X1 U738 ( .A1(rdata_L0[39]), .A2(n744), .ZN(n634) );
  AOI22_X1 U739 ( .A1(rdata_L0[7]), .A2(n892), .B1(rdata_last_q[7]), .B2(n871), 
        .ZN(n633) );
  OAI211_X1 U740 ( .C1(n635), .C2(n777), .A(n634), .B(n633), .ZN(n638) );
  AOI22_X1 U741 ( .A1(n638), .A2(n537), .B1(rdata_L0[102]), .B2(n32), .ZN(n636) );
  OAI21_X1 U742 ( .B1(n878), .B2(n537), .A(n636), .ZN(rdata_o[7]) );
  INV_X1 U743 ( .A(n638), .ZN(n641) );
  NAND2_X1 U744 ( .A1(n782), .A2(rdata_L0[102]), .ZN(n640) );
  AOI22_X1 U745 ( .A1(n547), .A2(rdata_last_q[7]), .B1(n12), .B2(rdata_o[7]), 
        .ZN(n639) );
  OAI211_X1 U746 ( .C1(n641), .C2(n785), .A(n640), .B(n639), .ZN(n817) );
  AOI22_X1 U747 ( .A1(rdata_L0[119]), .A2(n755), .B1(rdata_last_q[24]), .B2(
        n538), .ZN(n645) );
  NAND2_X1 U748 ( .A1(rdata_L0[24]), .A2(n892), .ZN(n644) );
  NAND2_X1 U749 ( .A1(rdata_L0[87]), .A2(n756), .ZN(n643) );
  NAND2_X1 U750 ( .A1(rdata_L0[56]), .A2(n773), .ZN(n642) );
  AOI22_X1 U753 ( .A1(rdata_L0[40]), .A2(n762), .B1(rdata_L0[103]), .B2(n42), 
        .ZN(n647) );
  AOI22_X1 U754 ( .A1(rdata_L0[8]), .A2(n31), .B1(rdata_L0[72]), .B2(n34), 
        .ZN(n646) );
  OAI211_X1 U755 ( .C1(n886), .C2(n765), .A(n647), .B(n646), .ZN(rdata_o[24])
         );
  INV_X1 U759 ( .A(rdata_L0[72]), .ZN(n653) );
  NAND2_X1 U760 ( .A1(rdata_L0[40]), .A2(n744), .ZN(n652) );
  AOI22_X1 U761 ( .A1(rdata_L0[8]), .A2(n892), .B1(rdata_last_q[8]), .B2(n871), 
        .ZN(n651) );
  OAI211_X1 U762 ( .C1(n653), .C2(n777), .A(n652), .B(n651), .ZN(n656) );
  AOI22_X1 U763 ( .A1(n656), .A2(n537), .B1(rdata_L0[103]), .B2(n32), .ZN(n654) );
  OAI21_X1 U764 ( .B1(n886), .B2(n537), .A(n654), .ZN(rdata_o[8]) );
  INV_X1 U765 ( .A(n656), .ZN(n659) );
  NAND2_X1 U766 ( .A1(n782), .A2(rdata_L0[103]), .ZN(n658) );
  AOI22_X1 U767 ( .A1(n547), .A2(rdata_last_q[8]), .B1(n12), .B2(rdata_o[8]), 
        .ZN(n657) );
  OAI211_X1 U768 ( .C1(n659), .C2(n785), .A(n658), .B(n657), .ZN(n816) );
  AOI22_X1 U769 ( .A1(rdata_L0[120]), .A2(n755), .B1(rdata_last_q[25]), .B2(
        n871), .ZN(n663) );
  NAND2_X1 U770 ( .A1(rdata_L0[25]), .A2(n892), .ZN(n662) );
  NAND2_X1 U771 ( .A1(rdata_L0[88]), .A2(n756), .ZN(n661) );
  NAND2_X1 U772 ( .A1(rdata_L0[57]), .A2(n744), .ZN(n660) );
  AOI22_X1 U775 ( .A1(rdata_L0[41]), .A2(n762), .B1(rdata_L0[104]), .B2(n42), 
        .ZN(n665) );
  AOI22_X1 U776 ( .A1(rdata_L0[9]), .A2(n31), .B1(rdata_L0[73]), .B2(n34), 
        .ZN(n664) );
  OAI211_X1 U777 ( .C1(n877), .C2(n765), .A(n665), .B(n664), .ZN(rdata_o[25])
         );
  INV_X1 U781 ( .A(rdata_L0[73]), .ZN(n671) );
  NAND2_X1 U782 ( .A1(rdata_L0[41]), .A2(n744), .ZN(n670) );
  AOI22_X1 U783 ( .A1(rdata_L0[9]), .A2(n774), .B1(rdata_last_q[9]), .B2(n871), 
        .ZN(n669) );
  OAI211_X1 U784 ( .C1(n671), .C2(n777), .A(n670), .B(n669), .ZN(n674) );
  AOI22_X1 U785 ( .A1(n674), .A2(n537), .B1(rdata_L0[104]), .B2(n32), .ZN(n672) );
  OAI21_X1 U786 ( .B1(n877), .B2(n537), .A(n672), .ZN(rdata_o[9]) );
  INV_X1 U787 ( .A(n674), .ZN(n677) );
  NAND2_X1 U788 ( .A1(n782), .A2(rdata_L0[104]), .ZN(n676) );
  AOI22_X1 U789 ( .A1(n547), .A2(rdata_last_q[9]), .B1(n12), .B2(rdata_o[9]), 
        .ZN(n675) );
  OAI211_X1 U790 ( .C1(n677), .C2(n785), .A(n676), .B(n675), .ZN(n815) );
  AOI22_X1 U791 ( .A1(rdata_L0[121]), .A2(n755), .B1(rdata_last_q[26]), .B2(
        n871), .ZN(n681) );
  NAND2_X1 U792 ( .A1(rdata_L0[26]), .A2(n774), .ZN(n680) );
  NAND2_X1 U793 ( .A1(rdata_L0[89]), .A2(n756), .ZN(n679) );
  NAND2_X1 U794 ( .A1(rdata_L0[58]), .A2(n773), .ZN(n678) );
  AOI22_X1 U797 ( .A1(rdata_L0[42]), .A2(n762), .B1(rdata_L0[105]), .B2(n42), 
        .ZN(n683) );
  AOI22_X1 U798 ( .A1(rdata_L0[10]), .A2(n31), .B1(rdata_L0[74]), .B2(n34), 
        .ZN(n682) );
  OAI211_X1 U799 ( .C1(n876), .C2(n765), .A(n683), .B(n682), .ZN(rdata_o[26])
         );
  INV_X1 U803 ( .A(rdata_L0[74]), .ZN(n689) );
  NAND2_X1 U804 ( .A1(rdata_L0[42]), .A2(n773), .ZN(n688) );
  AOI22_X1 U805 ( .A1(rdata_L0[10]), .A2(n892), .B1(rdata_last_q[10]), .B2(
        n871), .ZN(n687) );
  OAI211_X1 U806 ( .C1(n689), .C2(n777), .A(n688), .B(n687), .ZN(n692) );
  AOI22_X1 U807 ( .A1(n692), .A2(n537), .B1(rdata_L0[105]), .B2(n32), .ZN(n690) );
  OAI21_X1 U808 ( .B1(n876), .B2(n537), .A(n690), .ZN(rdata_o[10]) );
  INV_X1 U809 ( .A(n692), .ZN(n695) );
  NAND2_X1 U810 ( .A1(n782), .A2(rdata_L0[105]), .ZN(n694) );
  AOI22_X1 U811 ( .A1(n547), .A2(rdata_last_q[10]), .B1(n12), .B2(rdata_o[10]), 
        .ZN(n693) );
  OAI211_X1 U812 ( .C1(n695), .C2(n785), .A(n694), .B(n693), .ZN(n814) );
  AOI22_X1 U813 ( .A1(rdata_L0[122]), .A2(n755), .B1(rdata_last_q[27]), .B2(
        n871), .ZN(n699) );
  NAND2_X1 U814 ( .A1(rdata_L0[27]), .A2(n892), .ZN(n698) );
  NAND2_X1 U815 ( .A1(rdata_L0[90]), .A2(n756), .ZN(n697) );
  NAND2_X1 U816 ( .A1(rdata_L0[59]), .A2(n744), .ZN(n696) );
  AOI22_X1 U819 ( .A1(rdata_L0[43]), .A2(n762), .B1(rdata_L0[106]), .B2(n42), 
        .ZN(n701) );
  AOI22_X1 U820 ( .A1(rdata_L0[11]), .A2(n31), .B1(rdata_L0[75]), .B2(n34), 
        .ZN(n700) );
  OAI211_X1 U821 ( .C1(n875), .C2(n765), .A(n701), .B(n700), .ZN(rdata_o[27])
         );
  INV_X1 U825 ( .A(rdata_L0[75]), .ZN(n707) );
  NAND2_X1 U826 ( .A1(rdata_L0[43]), .A2(n744), .ZN(n706) );
  AOI22_X1 U827 ( .A1(rdata_L0[11]), .A2(n892), .B1(rdata_last_q[11]), .B2(
        n871), .ZN(n705) );
  OAI211_X1 U828 ( .C1(n707), .C2(n777), .A(n706), .B(n705), .ZN(n710) );
  AOI22_X1 U829 ( .A1(n710), .A2(n537), .B1(rdata_L0[106]), .B2(n32), .ZN(n708) );
  OAI21_X1 U830 ( .B1(n875), .B2(n537), .A(n708), .ZN(rdata_o[11]) );
  INV_X1 U831 ( .A(n710), .ZN(n713) );
  NAND2_X1 U832 ( .A1(n782), .A2(rdata_L0[106]), .ZN(n712) );
  AOI22_X1 U833 ( .A1(n547), .A2(rdata_last_q[11]), .B1(n769), .B2(rdata_o[11]), .ZN(n711) );
  OAI211_X1 U834 ( .C1(n713), .C2(n785), .A(n712), .B(n711), .ZN(n813) );
  AOI22_X1 U835 ( .A1(rdata_L0[44]), .A2(n762), .B1(rdata_L0[107]), .B2(n42), 
        .ZN(n715) );
  AOI22_X1 U836 ( .A1(rdata_L0[12]), .A2(n31), .B1(rdata_L0[76]), .B2(n34), 
        .ZN(n714) );
  OAI211_X1 U837 ( .C1(n885), .C2(n765), .A(n715), .B(n714), .ZN(rdata_o[28])
         );
  INV_X1 U841 ( .A(n720), .ZN(n723) );
  NAND2_X1 U842 ( .A1(n782), .A2(rdata_L0[107]), .ZN(n722) );
  AOI22_X1 U843 ( .A1(n547), .A2(rdata_last_q[12]), .B1(n769), .B2(rdata_o[12]), .ZN(n721) );
  OAI211_X1 U844 ( .C1(n723), .C2(n785), .A(n722), .B(n721), .ZN(n812) );
  AOI22_X1 U845 ( .A1(rdata_L0[45]), .A2(n762), .B1(rdata_L0[108]), .B2(n42), 
        .ZN(n725) );
  AOI22_X1 U846 ( .A1(rdata_L0[13]), .A2(n31), .B1(rdata_L0[77]), .B2(n34), 
        .ZN(n724) );
  OAI211_X1 U847 ( .C1(n884), .C2(n765), .A(n725), .B(n724), .ZN(rdata_o[29])
         );
  INV_X1 U851 ( .A(n730), .ZN(n733) );
  NAND2_X1 U852 ( .A1(n782), .A2(rdata_L0[108]), .ZN(n732) );
  AOI22_X1 U853 ( .A1(n547), .A2(rdata_last_q[13]), .B1(n769), .B2(rdata_o[13]), .ZN(n731) );
  OAI211_X1 U854 ( .C1(n733), .C2(n785), .A(n732), .B(n731), .ZN(n811) );
  AOI22_X1 U855 ( .A1(rdata_L0[125]), .A2(n755), .B1(rdata_last_q[30]), .B2(
        n871), .ZN(n738) );
  NAND2_X1 U856 ( .A1(rdata_L0[30]), .A2(n892), .ZN(n737) );
  NAND2_X1 U857 ( .A1(rdata_L0[93]), .A2(n756), .ZN(n736) );
  NAND2_X1 U858 ( .A1(rdata_L0[62]), .A2(n773), .ZN(n735) );
  AOI22_X1 U861 ( .A1(rdata_L0[46]), .A2(n762), .B1(rdata_L0[109]), .B2(n42), 
        .ZN(n740) );
  AOI22_X1 U862 ( .A1(rdata_L0[14]), .A2(n31), .B1(rdata_L0[78]), .B2(n34), 
        .ZN(n739) );
  OAI211_X1 U863 ( .C1(n874), .C2(n765), .A(n740), .B(n739), .ZN(rdata_o[30])
         );
  INV_X1 U867 ( .A(rdata_L0[78]), .ZN(n747) );
  NAND2_X1 U868 ( .A1(rdata_L0[46]), .A2(n744), .ZN(n746) );
  AOI22_X1 U869 ( .A1(rdata_L0[14]), .A2(n892), .B1(rdata_last_q[14]), .B2(
        n871), .ZN(n745) );
  OAI211_X1 U870 ( .C1(n747), .C2(n777), .A(n746), .B(n745), .ZN(n750) );
  AOI22_X1 U871 ( .A1(n750), .A2(n537), .B1(rdata_L0[109]), .B2(n32), .ZN(n748) );
  OAI21_X1 U872 ( .B1(n874), .B2(n537), .A(n748), .ZN(rdata_o[14]) );
  INV_X1 U873 ( .A(n750), .ZN(n753) );
  NAND2_X1 U874 ( .A1(n782), .A2(rdata_L0[109]), .ZN(n752) );
  AOI22_X1 U875 ( .A1(n547), .A2(rdata_last_q[14]), .B1(n769), .B2(rdata_o[14]), .ZN(n751) );
  OAI211_X1 U876 ( .C1(n753), .C2(n785), .A(n752), .B(n751), .ZN(n810) );
  AOI22_X1 U877 ( .A1(rdata_L0[126]), .A2(n755), .B1(rdata_last_q[31]), .B2(
        n871), .ZN(n760) );
  NAND2_X1 U878 ( .A1(rdata_L0[31]), .A2(n892), .ZN(n759) );
  NAND2_X1 U879 ( .A1(rdata_L0[94]), .A2(n756), .ZN(n758) );
  NAND2_X1 U880 ( .A1(rdata_L0[63]), .A2(n773), .ZN(n757) );
  NAND4_X1 U881 ( .A1(n760), .A2(n759), .A3(n758), .A4(n757), .ZN(n767) );
  INV_X1 U882 ( .A(n767), .ZN(n780) );
  AOI22_X1 U883 ( .A1(rdata_L0[47]), .A2(n762), .B1(rdata_L0[110]), .B2(n42), 
        .ZN(n764) );
  AOI22_X1 U884 ( .A1(rdata_L0[15]), .A2(n31), .B1(rdata_L0[79]), .B2(n34), 
        .ZN(n763) );
  OAI211_X1 U885 ( .C1(n780), .C2(n765), .A(n764), .B(n763), .ZN(rdata_o[31])
         );
  AOI22_X1 U886 ( .A1(n768), .A2(n767), .B1(n1042), .B2(rdata_last_q[31]), 
        .ZN(n772) );
  AOI22_X1 U887 ( .A1(n770), .A2(rdata_L0[126]), .B1(n769), .B2(rdata_o[31]), 
        .ZN(n771) );
  NAND2_X1 U888 ( .A1(n772), .A2(n771), .ZN(n792) );
  INV_X1 U889 ( .A(rdata_L0[79]), .ZN(n778) );
  NAND2_X1 U890 ( .A1(rdata_L0[47]), .A2(n773), .ZN(n776) );
  AOI22_X1 U891 ( .A1(rdata_L0[15]), .A2(n892), .B1(rdata_last_q[15]), .B2(
        n871), .ZN(n775) );
  OAI211_X1 U892 ( .C1(n778), .C2(n777), .A(n776), .B(n775), .ZN(n781) );
  AOI22_X1 U893 ( .A1(n781), .A2(n537), .B1(rdata_L0[110]), .B2(n32), .ZN(n779) );
  OAI21_X1 U894 ( .B1(n780), .B2(n537), .A(n779), .ZN(rdata_o[15]) );
  INV_X1 U895 ( .A(n781), .ZN(n786) );
  NAND2_X1 U896 ( .A1(n782), .A2(rdata_L0[110]), .ZN(n784) );
  AOI22_X1 U897 ( .A1(n547), .A2(rdata_last_q[15]), .B1(n12), .B2(rdata_o[15]), 
        .ZN(n783) );
  OAI211_X1 U898 ( .C1(n786), .C2(n785), .A(n784), .B(n783), .ZN(n809) );
  SDFFR_X1 rdata_last_q_reg_17_ ( .D(n1207), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[17]) );
  SDFFR_X1 rdata_last_q_reg_0_ ( .D(n823), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[0]) );
  SDFFR_X1 CS_reg_2_ ( .D(NS[2]), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(rst_n), 
        .Q(CS[2]), .QN(n829) );
  SDFFR_X1 addr_q_reg_0_ ( .D(addr_n[0]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[0]) );
  SDFFR_X1 addr_q_reg_3_ ( .D(addr_n[3]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[3]), .QN(n60) );
  SDFFR_X1 addr_q_reg_5_ ( .D(addr_n[5]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[5]), .QN(n848) );
  SDFFR_X1 addr_q_reg_6_ ( .D(addr_n[6]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[6]), .QN(n833) );
  SDFFR_X1 addr_q_reg_7_ ( .D(addr_n[7]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[7]), .QN(n847) );
  SDFFR_X1 addr_q_reg_8_ ( .D(addr_n[8]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[8]), .QN(n832) );
  SDFFR_X1 addr_q_reg_9_ ( .D(addr_n[9]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[9]), .QN(n844) );
  SDFFR_X1 addr_q_reg_10_ ( .D(addr_n[10]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[10]), .QN(n831) );
  SDFFR_X1 addr_q_reg_11_ ( .D(addr_n[11]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[11]), .QN(n839) );
  SDFFR_X1 addr_q_reg_12_ ( .D(addr_n[12]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[12]), .QN(n834) );
  SDFFR_X1 addr_q_reg_13_ ( .D(addr_n[13]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[13]), .QN(n836) );
  SDFFR_X1 addr_q_reg_14_ ( .D(addr_n[14]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[14]), .QN(n849) );
  SDFFR_X1 addr_q_reg_15_ ( .D(addr_n[15]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[15]), .QN(n835) );
  SDFFR_X1 addr_q_reg_16_ ( .D(addr_n[16]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[16]), .QN(n842) );
  SDFFR_X1 addr_q_reg_17_ ( .D(addr_n[17]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[17]), .QN(n840) );
  SDFFR_X1 addr_q_reg_18_ ( .D(addr_n[18]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[18]), .QN(n841) );
  SDFFR_X1 addr_q_reg_19_ ( .D(addr_n[19]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[19]), .QN(n837) );
  SDFFR_X1 addr_q_reg_20_ ( .D(addr_n[20]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[20]), .QN(n789) );
  SDFFR_X1 addr_q_reg_21_ ( .D(addr_n[21]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[21]), .QN(n852) );
  SDFFR_X1 addr_q_reg_22_ ( .D(addr_n[22]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[22]), .QN(n838) );
  SDFFR_X1 addr_q_reg_23_ ( .D(addr_n[23]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[23]), .QN(n38) );
  SDFFR_X1 addr_q_reg_24_ ( .D(addr_n[24]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[24]), .QN(n790) );
  SDFFR_X1 addr_q_reg_25_ ( .D(addr_n[25]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[25]), .QN(n791) );
  SDFFR_X1 addr_q_reg_26_ ( .D(addr_n[26]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[26]), .QN(n851) );
  SDFFR_X1 addr_q_reg_27_ ( .D(addr_n[27]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[27]), .QN(n850) );
  SDFFR_X1 rdata_last_q_reg_1_ ( .D(n824), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[1]) );
  SDFFR_X1 is_hwlp_q_reg ( .D(is_hwlp_n), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(is_hwlp_q) );
  SDFFR_X1 rdata_last_q_reg_16_ ( .D(n1208), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[16]), .QN(n830) );
  SDFFR_X1 rdata_last_q_reg_18_ ( .D(n1209), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[18]) );
  SDFFR_X1 rdata_last_q_reg_19_ ( .D(n1210), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[19]) );
  SDFFR_X1 rdata_last_q_reg_20_ ( .D(n1211), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[20]) );
  SDFFR_X1 rdata_last_q_reg_21_ ( .D(n1212), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[21]) );
  SDFFR_X1 rdata_last_q_reg_22_ ( .D(n1213), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[22]) );
  SDFFR_X1 rdata_last_q_reg_6_ ( .D(n818), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[6]) );
  SDFFR_X1 rdata_last_q_reg_23_ ( .D(n1214), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[23]) );
  SDFFR_X1 rdata_last_q_reg_7_ ( .D(n817), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[7]) );
  SDFFR_X1 rdata_last_q_reg_24_ ( .D(n1215), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[24]) );
  SDFFR_X1 rdata_last_q_reg_8_ ( .D(n816), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[8]) );
  SDFFR_X1 rdata_last_q_reg_25_ ( .D(n1216), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[25]) );
  SDFFR_X1 rdata_last_q_reg_9_ ( .D(n815), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[9]) );
  SDFFR_X1 rdata_last_q_reg_26_ ( .D(n1217), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[26]) );
  SDFFR_X1 rdata_last_q_reg_10_ ( .D(n814), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[10]) );
  SDFFR_X1 rdata_last_q_reg_27_ ( .D(n1218), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[27]) );
  SDFFR_X1 rdata_last_q_reg_11_ ( .D(n813), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[11]) );
  SDFFR_X1 rdata_last_q_reg_28_ ( .D(n1219), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[28]) );
  SDFFR_X1 rdata_last_q_reg_12_ ( .D(n812), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[12]) );
  SDFFR_X1 rdata_last_q_reg_29_ ( .D(n1220), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[29]) );
  SDFFR_X1 rdata_last_q_reg_13_ ( .D(n811), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[13]) );
  SDFFR_X1 rdata_last_q_reg_30_ ( .D(n1221), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[30]) );
  SDFFR_X1 rdata_last_q_reg_14_ ( .D(n810), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[14]) );
  SDFFR_X1 rdata_last_q_reg_31_ ( .D(n792), .SI(1'b0), .SE(1'b0), .CK(n1222), 
        .RN(rst_n), .Q(rdata_last_q[31]) );
  SDFFR_X1 rdata_last_q_reg_15_ ( .D(n809), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[15]) );
  SDFFR_X1 CS_reg_1_ ( .D(NS[1]), .SI(1'b0), .SE(1'b0), .CK(n1201), .RN(rst_n), 
        .Q(CS[1]), .QN(n793) );
  SDFFR_X1 addr_q_reg_4_ ( .D(addr_n[4]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[4]), .QN(n828) );
  SDFFR_X1 addr_q_reg_2_ ( .D(addr_n[2]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[2]), .QN(n826) );
  SDFFR_X1 CS_reg_3_ ( .D(NS[3]), .SI(1'b0), .SE(1'b0), .CK(n1201), .RN(rst_n), 
        .Q(CS[3]), .QN(n787) );
  SDFFR_X1 addr_q_reg_31_ ( .D(addr_n[31]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[31]), .QN(n853) );
  SDFFR_X1 addr_q_reg_30_ ( .D(addr_n[30]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[30]), .QN(n846) );
  SDFFR_X1 addr_q_reg_28_ ( .D(addr_n[28]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[28]), .QN(n845) );
  SDFFR_X1 addr_q_reg_29_ ( .D(addr_n[29]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[29]), .QN(n843) );
  SDFFR_X1 addr_q_reg_1_ ( .D(addr_n[1]), .SI(1'b0), .SE(1'b0), .CK(n1201), 
        .RN(rst_n), .Q(addr_o[1]), .QN(n827) );
  SDFFR_X1 CS_reg_0_ ( .D(NS[0]), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(rst_n), 
        .Q(CS[0]), .QN(n788) );
  AND2_X2 U112 ( .A1(n66), .A2(n826), .ZN(n756) );
  SDFFR_X2 rdata_last_q_reg_2_ ( .D(n822), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[2]) );
  SDFFR_X2 rdata_last_q_reg_3_ ( .D(n821), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[3]) );
  SDFFR_X2 rdata_last_q_reg_4_ ( .D(n820), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[4]) );
  SDFFR_X2 rdata_last_q_reg_5_ ( .D(n819), .SI(1'b0), .SE(1'b0), .CK(n1204), 
        .RN(rst_n), .Q(rdata_last_q[5]) );
  riscv_L0_buffer_RDATA_IN_WIDTH128 L0_buffer_i ( .clk(clk), .rst_n(rst_n), 
        .prefetch_i(n825), .prefetch_addr_i({addr_real_next, n43, 1'b0}), 
        .branch_i(branch_i), .branch_addr_i({addr_i[31:1], 1'b0}), .hwlp_i(
        n_0_net_), .hwlp_addr_i({hwloop_target_i[31:1], 1'b0}), .fetch_gnt_o(
        fetch_gnt), .fetch_valid_o(fetch_valid), .rdata_o({rdata_L0[126:97], 
        n872, rdata_L0[95:81], n855, rdata_L0[80:0]}), .addr_o({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, addr_L0, 
        SYNOPSYS_UNCONNECTED__28}), .instr_req_o(instr_req_o), .instr_addr_o({
        instr_addr_o[31:4], SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32}), .instr_gnt_i(
        instr_gnt_i), .instr_rvalid_i(instr_rvalid_i), .instr_rdata_i(
        instr_rdata_i), .busy_o(busy_o) );
  SNPS_CLOCK_GATE_HIGH_riscv_prefetch_L0_buffer_0 clk_gate_rdata_last_q_reg_31_ ( 
        .CLK(clk), .EN(n1224), .ENCLK(n1222), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_prefetch_L0_buffer_1 clk_gate_rdata_last_q_reg_15_ ( 
        .CLK(clk), .EN(n1206), .ENCLK(n1204), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_prefetch_L0_buffer_2 clk_gate_is_hwlp_q_reg ( 
        .CLK(clk), .EN(n1203), .ENCLK(n1201), .TE(1'b0) );
  OR2_X1 U7 ( .A1(n47), .A2(n71), .ZN(n124) );
  AND2_X1 U8 ( .A1(n39), .A2(n124), .ZN(n28) );
  CLKBUF_X1 U20 ( .A(n509), .Z(n43) );
  INV_X1 U3 ( .A(n594), .ZN(n12) );
  NOR2_X2 U309 ( .A1(n769), .A2(n545), .ZN(n547) );
  BUF_X1 U4 ( .A(n872), .Z(n863) );
  OAI211_X1 U5 ( .C1(n105), .C2(n64), .A(n894), .B(rdata_L0[111]), .ZN(n39) );
  NOR2_X1 U6 ( .A1(n769), .A2(n545), .ZN(n1042) );
  INV_X1 U9 ( .A(n182), .ZN(n545) );
  AND2_X2 U10 ( .A1(n39), .A2(n124), .ZN(n381) );
  INV_X4 U16 ( .A(n594), .ZN(n769) );
  NOR2_X1 U18 ( .A1(n182), .A2(n888), .ZN(n770) );
  INV_X1 U19 ( .A(n768), .ZN(n785) );
  INV_X1 U26 ( .A(n182), .ZN(n1197) );
  OR2_X1 U51 ( .A1(n353), .A2(n173), .ZN(n594) );
  AOI21_X2 U58 ( .B1(fetch_gnt), .B2(n180), .A(n179), .ZN(n182) );
  NOR2_X2 U65 ( .A1(n521), .A2(n306), .ZN(n873) );
  BUF_X2 U74 ( .A(ready_i), .Z(n521) );
  CLKBUF_X1 U82 ( .A(addr_i[24]), .Z(n889) );
  BUF_X1 U84 ( .A(n774), .Z(n892) );
  BUF_X4 U128 ( .A(n538), .Z(n871) );
  CLKBUF_X1 U132 ( .A(rdata_L0[111]), .Z(n893) );
  INV_X1 U138 ( .A(n381), .ZN(n7) );
  CLKBUF_X1 U139 ( .A(n773), .Z(n744) );
  INV_X2 U144 ( .A(n521), .ZN(n888) );
  INV_X2 U183 ( .A(n310), .ZN(n264) );
  AND4_X1 U184 ( .A1(n738), .A2(n737), .A3(n736), .A4(n735), .ZN(n874) );
  AND4_X1 U239 ( .A1(n699), .A2(n698), .A3(n697), .A4(n696), .ZN(n875) );
  AND4_X1 U274 ( .A1(n681), .A2(n680), .A3(n679), .A4(n678), .ZN(n876) );
  AND4_X1 U295 ( .A1(n663), .A2(n662), .A3(n661), .A4(n660), .ZN(n877) );
  AND4_X1 U297 ( .A1(n627), .A2(n626), .A3(n625), .A4(n624), .ZN(n878) );
  AND4_X1 U298 ( .A1(n609), .A2(n608), .A3(n607), .A4(n606), .ZN(n879) );
  AND4_X1 U305 ( .A1(n590), .A2(n589), .A3(n588), .A4(n587), .ZN(n880) );
  AND4_X1 U307 ( .A1(n572), .A2(n571), .A3(n570), .A4(n569), .ZN(n881) );
  AND4_X1 U308 ( .A1(n554), .A2(n553), .A3(n552), .A4(n551), .ZN(n882) );
  AND4_X1 U310 ( .A1(n531), .A2(n530), .A3(n529), .A4(n528), .ZN(n883) );
  AND4_X1 U311 ( .A1(n98), .A2(n97), .A3(n96), .A4(n95), .ZN(n884) );
  AND4_X1 U312 ( .A1(n76), .A2(n75), .A3(n74), .A4(n73), .ZN(n885) );
  AND4_X1 U489 ( .A1(n645), .A2(n644), .A3(n643), .A4(n642), .ZN(n886) );
  INV_X1 U490 ( .A(n521), .ZN(n887) );
  INV_X1 U491 ( .A(n521), .ZN(n510) );
  NOR2_X1 U584 ( .A1(n769), .A2(n181), .ZN(n768) );
  MUX2_X1 U616 ( .A(n478), .B(n479), .S(n381), .Z(addr_real_next[23]) );
  CLKBUF_X1 U617 ( .A(rdata_L0[95]), .Z(n890) );
  CLKBUF_X1 U621 ( .A(addr_i[23]), .Z(n891) );
  AND2_X1 U622 ( .A1(rdata_L0[112]), .A2(n63), .ZN(n894) );
  NAND3_X1 U623 ( .A1(n70), .A2(rdata_L0[111]), .A3(rdata_L0[112]), .ZN(n47)
         );
  OAI21_X1 U624 ( .B1(n1060), .B2(n1061), .A(n887), .ZN(n1059) );
  INV_X1 U632 ( .A(n1184), .ZN(n895) );
  NOR2_X1 U641 ( .A1(n182), .A2(n1186), .ZN(n896) );
  MUX2_X1 U642 ( .A(n895), .B(n896), .S(n1185), .Z(n1221) );
  INV_X2 U646 ( .A(n172), .ZN(n320) );
  OAI211_X1 U985 ( .C1(n829), .C2(CS[0]), .A(n1035), .B(n1036), .ZN(n1203) );
  NOR2_X1 U986 ( .A1(fetch_gnt), .A2(n1037), .ZN(n1036) );
  NAND3_X1 U987 ( .A1(CS[3]), .A2(n788), .A3(n172), .ZN(n1037) );
  NOR2_X1 U988 ( .A1(n521), .A2(CS[1]), .ZN(n1035) );
  OAI221_X1 U989 ( .B1(n769), .B2(n1038), .C1(n1185), .C2(n537), .A(n1039), 
        .ZN(n1206) );
  NOR2_X1 U990 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
  OAI21_X1 U991 ( .B1(n1042), .B2(n871), .A(n1043), .ZN(n1041) );
  OAI221_X1 U992 ( .B1(n1044), .B2(n892), .C1(n1044), .C2(rdata_L0[14]), .A(
        n1045), .ZN(n1043) );
  NAND2_X1 U993 ( .A1(n181), .A2(n1042), .ZN(n1045) );
  OAI21_X1 U994 ( .B1(n777), .B2(n747), .A(n746), .ZN(n1044) );
  AOI21_X1 U995 ( .B1(n1185), .B2(n546), .A(n1046), .ZN(n1040) );
  OAI21_X1 U996 ( .B1(n32), .B2(n1185), .A(rdata_L0[109]), .ZN(n1046) );
  NAND2_X1 U997 ( .A1(n181), .A2(n545), .ZN(n1038) );
  OAI21_X1 U998 ( .B1(n887), .B2(n1047), .A(n1048), .ZN(n1207) );
  AOI22_X1 U999 ( .A1(n888), .A2(n1049), .B1(n12), .B2(rdata_o[17]), .ZN(n1048) );
  NOR3_X1 U1000 ( .A1(n1050), .A2(n182), .A3(n769), .ZN(n1049) );
  OAI22_X1 U1001 ( .A1(n1051), .A2(n1052), .B1(n510), .B2(n1053), .ZN(n1050)
         );
  NAND3_X1 U1002 ( .A1(n120), .A2(n118), .A3(n117), .ZN(n1052) );
  NOR2_X1 U1003 ( .A1(n306), .A2(n1053), .ZN(n1051) );
  INV_X1 U1004 ( .A(n41), .ZN(n1053) );
  NAND2_X1 U1005 ( .A1(n41), .A2(n1197), .ZN(n1047) );
  OAI21_X1 U1006 ( .B1(n1054), .B2(n769), .A(n1055), .ZN(n1208) );
  OAI221_X1 U1007 ( .B1(rdata_o[16]), .B2(n893), .C1(rdata_o[16]), .C2(n770), 
        .A(n769), .ZN(n1055) );
  AOI21_X1 U1008 ( .B1(n1056), .B2(n1197), .A(n1057), .ZN(n1054) );
  AOI21_X1 U1009 ( .B1(n1058), .B2(n1059), .A(n182), .ZN(n1057) );
  OAI21_X1 U1010 ( .B1(n306), .B2(n1062), .A(n112), .ZN(n1061) );
  NAND2_X1 U1011 ( .A1(n115), .A2(n114), .ZN(n1060) );
  OAI211_X1 U1012 ( .C1(n1063), .C2(n1064), .A(n887), .B(n1062), .ZN(n1058) );
  INV_X1 U1013 ( .A(n112), .ZN(n1064) );
  AOI21_X1 U1014 ( .B1(n115), .B2(n114), .A(n1165), .ZN(n1063) );
  NOR2_X1 U1015 ( .A1(n888), .A2(n1062), .ZN(n1056) );
  INV_X1 U1016 ( .A(n893), .ZN(n1062) );
  OAI21_X1 U1017 ( .B1(n510), .B2(n1065), .A(n1066), .ZN(n1209) );
  AOI22_X1 U1018 ( .A1(n1134), .A2(n1067), .B1(n12), .B2(rdata_o[18]), .ZN(
        n1066) );
  OAI21_X1 U1019 ( .B1(n1068), .B2(n1069), .A(n1070), .ZN(n1067) );
  OAI211_X1 U1020 ( .C1(n887), .C2(n1071), .A(n510), .B(n1068), .ZN(n1070) );
  INV_X1 U1021 ( .A(rdata_L0[113]), .ZN(n1071) );
  NAND3_X1 U1022 ( .A1(rdata_L0[113]), .A2(n873), .A3(n510), .ZN(n1069) );
  NAND3_X1 U1023 ( .A1(n528), .A2(n530), .A3(n529), .ZN(n1068) );
  NAND2_X1 U1024 ( .A1(rdata_L0[113]), .A2(n1197), .ZN(n1065) );
  OAI21_X1 U1025 ( .B1(n888), .B2(n1072), .A(n1073), .ZN(n1210) );
  AOI22_X1 U1026 ( .A1(n1134), .A2(n1074), .B1(n12), .B2(rdata_o[19]), .ZN(
        n1073) );
  OAI21_X1 U1027 ( .B1(n1075), .B2(n1076), .A(n1077), .ZN(n1074) );
  OAI211_X1 U1028 ( .C1(n887), .C2(n1078), .A(n888), .B(n1075), .ZN(n1077) );
  INV_X1 U1029 ( .A(rdata_L0[114]), .ZN(n1078) );
  NAND3_X1 U1030 ( .A1(rdata_L0[114]), .A2(n873), .A3(n887), .ZN(n1076) );
  NAND3_X1 U1031 ( .A1(n551), .A2(n553), .A3(n552), .ZN(n1075) );
  NAND2_X1 U1032 ( .A1(rdata_L0[114]), .A2(n1197), .ZN(n1072) );
  OAI21_X1 U1033 ( .B1(n888), .B2(n1079), .A(n1080), .ZN(n1211) );
  AOI22_X1 U1034 ( .A1(n1134), .A2(n1081), .B1(n12), .B2(rdata_o[20]), .ZN(
        n1080) );
  OAI21_X1 U1035 ( .B1(n1082), .B2(n1083), .A(n1084), .ZN(n1081) );
  OAI211_X1 U1036 ( .C1(n888), .C2(n1085), .A(n887), .B(n1082), .ZN(n1084) );
  INV_X1 U1037 ( .A(rdata_L0[115]), .ZN(n1085) );
  NAND3_X1 U1038 ( .A1(rdata_L0[115]), .A2(n873), .A3(n510), .ZN(n1083) );
  NAND3_X1 U1039 ( .A1(n569), .A2(n571), .A3(n570), .ZN(n1082) );
  NAND2_X1 U1040 ( .A1(rdata_L0[115]), .A2(n1197), .ZN(n1079) );
  OAI21_X1 U1041 ( .B1(n887), .B2(n1086), .A(n1087), .ZN(n1212) );
  AOI22_X1 U1042 ( .A1(n1134), .A2(n1088), .B1(n12), .B2(rdata_o[21]), .ZN(
        n1087) );
  OAI21_X1 U1043 ( .B1(n1089), .B2(n1090), .A(n1091), .ZN(n1088) );
  OAI211_X1 U1044 ( .C1(n510), .C2(n1092), .A(n888), .B(n1089), .ZN(n1091) );
  INV_X1 U1045 ( .A(rdata_L0[116]), .ZN(n1092) );
  NAND3_X1 U1046 ( .A1(rdata_L0[116]), .A2(n873), .A3(n888), .ZN(n1090) );
  NAND3_X1 U1047 ( .A1(n587), .A2(n589), .A3(n588), .ZN(n1089) );
  NAND2_X1 U1048 ( .A1(rdata_L0[116]), .A2(n1197), .ZN(n1086) );
  OAI21_X1 U1049 ( .B1(n510), .B2(n1093), .A(n1094), .ZN(n1213) );
  AOI22_X1 U1050 ( .A1(rdata_o[22]), .A2(n12), .B1(n1134), .B2(n1095), .ZN(
        n1094) );
  OAI33_X1 U1051 ( .A1(n1096), .A2(n1181), .A3(n1097), .B1(n1098), .B2(n1099), 
        .B3(n1100), .ZN(n1095) );
  AOI22_X1 U1052 ( .A1(n1101), .A2(rdata_L0[117]), .B1(n888), .B2(n1102), .ZN(
        n1100) );
  AND3_X1 U1053 ( .A1(n607), .A2(n873), .A3(n608), .ZN(n1101) );
  AOI21_X1 U1054 ( .B1(n888), .B2(n1103), .A(n1104), .ZN(n1099) );
  OAI22_X1 U1055 ( .A1(n871), .A2(n1098), .B1(n1103), .B2(n1102), .ZN(n1097)
         );
  NAND2_X1 U1056 ( .A1(n608), .A2(n607), .ZN(n1102) );
  INV_X1 U1057 ( .A(n871), .ZN(n1103) );
  NOR2_X1 U1058 ( .A1(n167), .A2(n1105), .ZN(n1098) );
  INV_X1 U1059 ( .A(rdata_L0[54]), .ZN(n1105) );
  NOR2_X1 U1060 ( .A1(n510), .A2(n1104), .ZN(n1096) );
  INV_X1 U1061 ( .A(rdata_L0[117]), .ZN(n1104) );
  NAND2_X1 U1062 ( .A1(rdata_L0[117]), .A2(n1197), .ZN(n1093) );
  OAI21_X1 U1063 ( .B1(n888), .B2(n1106), .A(n1107), .ZN(n1214) );
  AOI22_X1 U1064 ( .A1(n1134), .A2(n1108), .B1(n12), .B2(rdata_o[23]), .ZN(
        n1107) );
  OAI21_X1 U1065 ( .B1(n1109), .B2(n1110), .A(n1111), .ZN(n1108) );
  OAI211_X1 U1066 ( .C1(n888), .C2(n1112), .A(n887), .B(n1109), .ZN(n1111) );
  INV_X1 U1067 ( .A(rdata_L0[118]), .ZN(n1112) );
  NAND3_X1 U1068 ( .A1(rdata_L0[118]), .A2(n873), .A3(n510), .ZN(n1110) );
  NAND3_X1 U1069 ( .A1(n624), .A2(n626), .A3(n625), .ZN(n1109) );
  NAND2_X1 U1070 ( .A1(rdata_L0[118]), .A2(n1197), .ZN(n1106) );
  OAI21_X1 U1071 ( .B1(n887), .B2(n1113), .A(n1114), .ZN(n1215) );
  AOI22_X1 U1072 ( .A1(rdata_o[24]), .A2(n12), .B1(n1134), .B2(n1115), .ZN(
        n1114) );
  OAI33_X1 U1073 ( .A1(n1116), .A2(n1181), .A3(n1117), .B1(n1118), .B2(n1119), 
        .B3(n1120), .ZN(n1115) );
  AOI22_X1 U1074 ( .A1(n1121), .A2(rdata_L0[119]), .B1(n888), .B2(n1122), .ZN(
        n1120) );
  AND3_X1 U1075 ( .A1(n643), .A2(n873), .A3(n644), .ZN(n1121) );
  AOI21_X1 U1076 ( .B1(n887), .B2(n1103), .A(n1123), .ZN(n1119) );
  OAI22_X1 U1077 ( .A1(n871), .A2(n1118), .B1(n1103), .B2(n1122), .ZN(n1117)
         );
  NAND2_X1 U1078 ( .A1(n644), .A2(n643), .ZN(n1122) );
  NOR2_X1 U1079 ( .A1(n167), .A2(n1124), .ZN(n1118) );
  INV_X1 U1080 ( .A(rdata_L0[56]), .ZN(n1124) );
  NOR2_X1 U1081 ( .A1(n888), .A2(n1123), .ZN(n1116) );
  INV_X1 U1082 ( .A(rdata_L0[119]), .ZN(n1123) );
  NAND2_X1 U1083 ( .A1(rdata_L0[119]), .A2(n1197), .ZN(n1113) );
  OAI21_X1 U1084 ( .B1(n510), .B2(n1125), .A(n1126), .ZN(n1216) );
  AOI22_X1 U1085 ( .A1(n1134), .A2(n1127), .B1(n12), .B2(rdata_o[25]), .ZN(
        n1126) );
  OAI21_X1 U1086 ( .B1(n1128), .B2(n1129), .A(n1130), .ZN(n1127) );
  OAI211_X1 U1087 ( .C1(n510), .C2(n1131), .A(n888), .B(n1128), .ZN(n1130) );
  INV_X1 U1088 ( .A(rdata_L0[120]), .ZN(n1131) );
  NAND3_X1 U1089 ( .A1(rdata_L0[120]), .A2(n873), .A3(n510), .ZN(n1129) );
  NAND3_X1 U1090 ( .A1(n660), .A2(n662), .A3(n661), .ZN(n1128) );
  NAND2_X1 U1091 ( .A1(rdata_L0[120]), .A2(n1197), .ZN(n1125) );
  OAI21_X1 U1092 ( .B1(n888), .B2(n1132), .A(n1133), .ZN(n1217) );
  AOI22_X1 U1093 ( .A1(rdata_o[26]), .A2(n12), .B1(n1134), .B2(n1135), .ZN(
        n1133) );
  OAI33_X1 U1094 ( .A1(n1136), .A2(n1165), .A3(n1137), .B1(n1138), .B2(n1139), 
        .B3(n1140), .ZN(n1135) );
  AOI22_X1 U1095 ( .A1(n1141), .A2(rdata_L0[121]), .B1(n888), .B2(n1142), .ZN(
        n1140) );
  AND3_X1 U1096 ( .A1(n679), .A2(n873), .A3(n680), .ZN(n1141) );
  AOI21_X1 U1097 ( .B1(n888), .B2(n1103), .A(n1143), .ZN(n1139) );
  OAI22_X1 U1098 ( .A1(n871), .A2(n1138), .B1(n1103), .B2(n1142), .ZN(n1137)
         );
  NAND2_X1 U1099 ( .A1(n680), .A2(n679), .ZN(n1142) );
  NOR2_X1 U1100 ( .A1(n167), .A2(n1144), .ZN(n1138) );
  INV_X1 U1101 ( .A(rdata_L0[58]), .ZN(n1144) );
  NOR2_X1 U1102 ( .A1(n887), .A2(n1143), .ZN(n1136) );
  INV_X1 U1103 ( .A(rdata_L0[121]), .ZN(n1143) );
  NOR2_X1 U1104 ( .A1(n182), .A2(n769), .ZN(n1134) );
  NAND2_X1 U1105 ( .A1(rdata_L0[121]), .A2(n1197), .ZN(n1132) );
  OAI21_X1 U1106 ( .B1(n769), .B2(n1145), .A(n1146), .ZN(n1218) );
  OAI221_X1 U1107 ( .B1(rdata_o[27]), .B2(rdata_L0[122]), .C1(rdata_o[27]), 
        .C2(n770), .A(n769), .ZN(n1146) );
  AOI22_X1 U1108 ( .A1(rdata_L0[122]), .A2(n1147), .B1(n1225), .B2(n1148), 
        .ZN(n1145) );
  NOR2_X1 U1109 ( .A1(rdata_L0[122]), .A2(n182), .ZN(n1148) );
  OAI22_X1 U1110 ( .A1(n182), .A2(n1149), .B1(n888), .B2(n1150), .ZN(n1147) );
  INV_X1 U1111 ( .A(n1197), .ZN(n1150) );
  OAI221_X1 U1112 ( .B1(n1151), .B2(n888), .C1(n1152), .C2(n873), .A(n888), 
        .ZN(n1149) );
  INV_X1 U1113 ( .A(n1152), .ZN(n1151) );
  NAND3_X1 U1114 ( .A1(n696), .A2(n698), .A3(n697), .ZN(n1152) );
  OAI21_X1 U1115 ( .B1(n1153), .B2(n769), .A(n1154), .ZN(n1219) );
  OAI221_X1 U1116 ( .B1(rdata_o[28]), .B2(n770), .C1(rdata_o[28]), .C2(
        rdata_L0[123]), .A(n769), .ZN(n1154) );
  AOI21_X1 U1117 ( .B1(n1155), .B2(n1197), .A(n1156), .ZN(n1153) );
  AOI221_X1 U1118 ( .B1(n1158), .B2(n1157), .C1(n1155), .C2(n1158), .A(n182), 
        .ZN(n1156) );
  OAI221_X1 U1119 ( .B1(rdata_L0[123]), .B2(n1159), .C1(n1160), .C2(n1161), 
        .A(n1162), .ZN(n1158) );
  AOI211_X1 U1120 ( .C1(n1163), .C2(n1164), .A(n871), .B(n1165), .ZN(n1161) );
  INV_X1 U1121 ( .A(n510), .ZN(n1165) );
  NAND3_X1 U1122 ( .A1(n75), .A2(n74), .A3(n873), .ZN(n1164) );
  INV_X1 U1123 ( .A(n1159), .ZN(n1163) );
  AOI21_X1 U1124 ( .B1(n75), .B2(n74), .A(n1165), .ZN(n1159) );
  OAI211_X1 U1125 ( .C1(n871), .C2(n1166), .A(n1167), .B(n888), .ZN(n1157) );
  NAND3_X1 U1126 ( .A1(n75), .A2(n74), .A3(n871), .ZN(n1167) );
  INV_X1 U1127 ( .A(n1162), .ZN(n1166) );
  NAND2_X1 U1128 ( .A1(rdata_L0[60]), .A2(n1168), .ZN(n1162) );
  INV_X1 U1129 ( .A(n167), .ZN(n1168) );
  NOR2_X1 U1130 ( .A1(n887), .A2(n1160), .ZN(n1155) );
  INV_X1 U1131 ( .A(rdata_L0[123]), .ZN(n1160) );
  OAI21_X1 U1132 ( .B1(n1169), .B2(n769), .A(n1170), .ZN(n1220) );
  OAI221_X1 U1133 ( .B1(rdata_o[29]), .B2(n770), .C1(rdata_o[29]), .C2(
        rdata_L0[124]), .A(n769), .ZN(n1170) );
  AOI21_X1 U1134 ( .B1(n1171), .B2(n1197), .A(n1172), .ZN(n1169) );
  AOI221_X1 U1135 ( .B1(n1173), .B2(n1174), .C1(n1171), .C2(n1174), .A(n182), 
        .ZN(n1172) );
  OAI221_X1 U1136 ( .B1(rdata_L0[124]), .B2(n1175), .C1(n1176), .C2(n1177), 
        .A(n1178), .ZN(n1174) );
  AOI211_X1 U1137 ( .C1(n1179), .C2(n1180), .A(n871), .B(n1181), .ZN(n1177) );
  INV_X1 U1138 ( .A(n887), .ZN(n1181) );
  NAND3_X1 U1139 ( .A1(n97), .A2(n96), .A3(n873), .ZN(n1180) );
  INV_X1 U1140 ( .A(n1175), .ZN(n1179) );
  AOI21_X1 U1141 ( .B1(n97), .B2(n96), .A(n1181), .ZN(n1175) );
  OAI211_X1 U1142 ( .C1(n871), .C2(n1182), .A(n1183), .B(n888), .ZN(n1173) );
  NAND3_X1 U1143 ( .A1(n97), .A2(n96), .A3(n871), .ZN(n1183) );
  INV_X1 U1144 ( .A(n1178), .ZN(n1182) );
  NAND2_X1 U1145 ( .A1(rdata_L0[61]), .A2(n1168), .ZN(n1178) );
  NOR2_X1 U1146 ( .A1(n888), .A2(n1176), .ZN(n1171) );
  INV_X1 U1147 ( .A(rdata_L0[124]), .ZN(n1176) );
  AOI221_X1 U1148 ( .B1(n1187), .B2(n510), .C1(n1188), .C2(n887), .A(n1189), 
        .ZN(n1186) );
  AOI221_X1 U1149 ( .B1(n1190), .B2(n888), .C1(n1191), .C2(n888), .A(n1192), 
        .ZN(n1189) );
  INV_X1 U1150 ( .A(rdata_L0[125]), .ZN(n1192) );
  NAND4_X1 U1151 ( .A1(n873), .A2(n737), .A3(n1103), .A4(n1193), .ZN(n1191) );
  INV_X1 U1152 ( .A(n736), .ZN(n1190) );
  NAND2_X1 U1153 ( .A1(n736), .A2(n737), .ZN(n1188) );
  NOR2_X1 U1154 ( .A1(n871), .A2(n1193), .ZN(n1187) );
  NAND2_X1 U1155 ( .A1(rdata_L0[62]), .A2(n1168), .ZN(n1193) );
  INV_X1 U1156 ( .A(n769), .ZN(n1185) );
  AOI21_X1 U1157 ( .B1(n770), .B2(rdata_L0[125]), .A(rdata_o[30]), .ZN(n1184)
         );
  NAND2_X1 U1158 ( .A1(n1194), .A2(n1195), .ZN(n1224) );
  AOI21_X1 U1159 ( .B1(n1196), .B2(n545), .A(n769), .ZN(n1195) );
  NAND3_X1 U1160 ( .A1(n871), .A2(n1197), .A3(n510), .ZN(n1196) );
  OAI221_X1 U1161 ( .B1(n1225), .B2(rdata_L0[122]), .C1(n1225), .C2(n1198), 
        .A(n1197), .ZN(n1194) );
  OAI21_X1 U1162 ( .B1(n871), .B2(n1199), .A(n887), .ZN(n1198) );
  INV_X1 U1163 ( .A(n873), .ZN(n1199) );
  AND2_X1 U1164 ( .A1(n1200), .A2(n510), .ZN(n1225) );
  NAND3_X1 U1165 ( .A1(n698), .A2(n697), .A3(n696), .ZN(n1200) );
endmodule


module riscv_pmp_N_PMP_ENTRIES16 ( clk, rst_n, pmp_privil_mode_i, pmp_addr_i, 
        pmp_cfg_i, data_req_i, data_addr_i, data_we_i, data_gnt_o, data_req_o, 
        data_gnt_i, instr_req_i, instr_addr_i, instr_gnt_o, instr_req_o, 
        instr_gnt_i, instr_err_o, data_err_ack_i_BAR, data_err_o_BAR, 
        instr_addr_o_31_, instr_addr_o_30_, instr_addr_o_29_, instr_addr_o_28_, 
        instr_addr_o_27_, instr_addr_o_26_, instr_addr_o_25_, instr_addr_o_24_, 
        instr_addr_o_23_, instr_addr_o_22_, instr_addr_o_21_, instr_addr_o_20_, 
        instr_addr_o_19_, instr_addr_o_17_, instr_addr_o_16_, instr_addr_o_15_, 
        instr_addr_o_13_, instr_addr_o_12_, instr_addr_o_11_, instr_addr_o_10_, 
        instr_addr_o_9_, instr_addr_o_8_, instr_addr_o_7_, instr_addr_o_6_, 
        instr_addr_o_5_, instr_addr_o_3_, instr_addr_o_2_, instr_addr_o_1_, 
        instr_addr_o_0_, data_addr_o_30_, data_addr_o_29_, data_addr_o_28_, 
        data_addr_o_27_, data_addr_o_26_, data_addr_o_25_, data_addr_o_24_, 
        data_addr_o_23_, data_addr_o_22_, data_addr_o_21_, data_addr_o_20_, 
        data_addr_o_19_, data_addr_o_18_, data_addr_o_17_, data_addr_o_16_, 
        data_addr_o_15_, data_addr_o_14_, data_addr_o_13_, data_addr_o_12_, 
        data_addr_o_11_, data_addr_o_10_, data_addr_o_9_, data_addr_o_8_, 
        data_addr_o_7_, data_addr_o_6_, data_addr_o_5_, data_addr_o_4_, 
        data_addr_o_3_, data_addr_o_2_, data_addr_o_1_, data_addr_o_0_, 
        instr_addr_o_18_, instr_addr_o_14_, instr_addr_o_4_, data_addr_o_31_
 );
  input [1:0] pmp_privil_mode_i;
  input [511:0] pmp_addr_i;
  input [127:0] pmp_cfg_i;
  input [31:0] data_addr_i;
  input [31:0] instr_addr_i;
  input clk, rst_n, data_req_i, data_we_i, data_gnt_i, instr_req_i,
         instr_gnt_i, data_err_ack_i_BAR;
  output data_gnt_o, data_req_o, instr_gnt_o, instr_req_o, instr_err_o,
         data_err_o_BAR, instr_addr_o_31_, instr_addr_o_30_, instr_addr_o_29_,
         instr_addr_o_28_, instr_addr_o_27_, instr_addr_o_26_,
         instr_addr_o_25_, instr_addr_o_24_, instr_addr_o_23_,
         instr_addr_o_22_, instr_addr_o_21_, instr_addr_o_20_,
         instr_addr_o_19_, instr_addr_o_17_, instr_addr_o_16_,
         instr_addr_o_15_, instr_addr_o_13_, instr_addr_o_12_,
         instr_addr_o_11_, instr_addr_o_10_, instr_addr_o_9_, instr_addr_o_8_,
         instr_addr_o_7_, instr_addr_o_6_, instr_addr_o_5_, instr_addr_o_3_,
         instr_addr_o_2_, instr_addr_o_1_, instr_addr_o_0_, data_addr_o_30_,
         data_addr_o_29_, data_addr_o_28_, data_addr_o_27_, data_addr_o_26_,
         data_addr_o_25_, data_addr_o_24_, data_addr_o_23_, data_addr_o_22_,
         data_addr_o_21_, data_addr_o_20_, data_addr_o_19_, data_addr_o_18_,
         data_addr_o_17_, data_addr_o_16_, data_addr_o_15_, data_addr_o_14_,
         data_addr_o_13_, data_addr_o_12_, data_addr_o_11_, data_addr_o_10_,
         data_addr_o_9_, data_addr_o_8_, data_addr_o_7_, data_addr_o_6_,
         data_addr_o_5_, data_addr_o_4_, data_addr_o_3_, data_addr_o_2_,
         data_addr_o_1_, data_addr_o_0_, instr_addr_o_18_, instr_addr_o_14_,
         instr_addr_o_4_, data_addr_o_31_;
  wire   data_err_state_q, n4177, gte_x_382_A_16_, n12260, n1, n2, n3, n4, n7,
         n8, n9, n10, n11, n12, n13, n15, n16, n17, n18, n19, n20,
         data_addr_o_31__BAR, n22, n23, n24, n29, n31, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n142, n143,
         n146, n147, n149, n150, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n191, n192, n193,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n12265, n210, n212, n213, n214, n215, n217, n218,
         n219, n220, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n233, n234, n235, n236, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         instr_addr_o_4__BAR, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n12266, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4541, n4542, n4543, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n12263, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, instr_addr_o_18__BAR, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5432,
         n5433, n5434, n5436, n5437, n5439, n5440, n5441, n5442, n5443, n5444,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, instr_addr_o_14__BAR, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5999, n6000,
         n6001, n6002, n6003, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12150, n12152, n12267,
         n12156, n12157, n12158, n12264, n12161, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12192, n12193, n12194, n12195, n12197, n12198, n12199,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257;
  assign data_addr_o_8_ = data_addr_i[8];
  assign data_addr_o_1_ = data_addr_i[1];
  assign data_addr_o_0_ = data_addr_i[0];
  assign data_addr_o_22_ = data_addr_i[22];
  assign data_addr_o_24_ = data_addr_i[24];
  assign data_addr_o_19_ = data_addr_i[19];
  assign data_addr_o_28_ = data_addr_i[28];
  assign data_addr_o_21_ = data_addr_i[21];
  assign data_addr_o_27_ = data_addr_i[27];
  assign data_addr_o_31_ = n24;
  assign instr_addr_o_17_ = n4069;
  assign instr_addr_o_7_ = n4605;
  assign instr_addr_o_18_ = n4908;
  assign instr_addr_o_4_ = n5291;
  assign instr_addr_o_30_ = n5980;
  assign data_addr_o_18_ = n10967;
  assign data_addr_o_25_ = n11320;

  AOI21_X1 U5 ( .B1(n1291), .B2(n1290), .A(n1289), .ZN(n1301) );
  AND2_X1 U6 ( .A1(n4234), .A2(n8254), .ZN(n4966) );
  OAI21_X1 U7 ( .B1(n5663), .B2(n4266), .A(n1976), .ZN(n6314) );
  NOR2_X1 U14 ( .A1(n267), .A2(n1), .ZN(n127) );
  NAND4_X1 U15 ( .A1(n129), .A2(n4683), .A3(n4679), .A4(n4682), .ZN(n1) );
  NAND4_X1 U17 ( .A1(n5828), .A2(n2), .A3(n198), .A4(n5827), .ZN(n6041) );
  OAI211_X1 U19 ( .C1(n5055), .C2(n3), .A(n5079), .B(n5054), .ZN(n5082) );
  NAND2_X1 U20 ( .A1(n5045), .A2(n5044), .ZN(n3) );
  INV_X2 U21 ( .A(n511), .ZN(n4866) );
  OR2_X1 U22 ( .A1(n4234), .A2(n7322), .ZN(n4254) );
  NAND4_X1 U23 ( .A1(n67), .A2(n234), .A3(n5013), .A4(n4), .ZN(n5015) );
  NOR3_X1 U24 ( .A1(n4945), .A2(n4947), .A3(n4946), .ZN(n4) );
  NAND2_X1 U31 ( .A1(n2035), .A2(n8), .ZN(n233) );
  AND2_X1 U32 ( .A1(n3846), .A2(pmp_addr_i[487]), .ZN(n4088) );
  NOR2_X1 U35 ( .A1(n2033), .A2(n2032), .ZN(n8) );
  NAND2_X1 U36 ( .A1(n2013), .A2(n9), .ZN(n2030) );
  NAND3_X1 U40 ( .A1(n10), .A2(n2118), .A3(n2110), .ZN(n2133) );
  OAI21_X1 U41 ( .B1(n2108), .B2(n2107), .A(n2106), .ZN(n10) );
  OAI211_X1 U43 ( .C1(n1568), .C2(n1567), .A(n12), .B(n11), .ZN(n1569) );
  NAND2_X1 U44 ( .A1(instr_addr_o_18__BAR), .A2(pmp_addr_i[400]), .ZN(n11) );
  NAND2_X1 U45 ( .A1(n1564), .A2(n1565), .ZN(n12) );
  NAND3_X1 U46 ( .A1(n238), .A2(n321), .A3(n2747), .ZN(n308) );
  NAND3_X1 U47 ( .A1(n13), .A2(n1146), .A3(n315), .ZN(n1405) );
  NAND2_X1 U48 ( .A1(n96), .A2(n1040), .ZN(n13) );
  AND2_X1 U49 ( .A1(n4234), .A2(n10290), .ZN(n3002) );
  NAND2_X1 U50 ( .A1(n15), .A2(n9019), .ZN(n9023) );
  NAND2_X2 U55 ( .A1(n11595), .A2(n9009), .ZN(n5783) );
  INV_X2 U56 ( .A(n3531), .ZN(n208) );
  INV_X1 U58 ( .A(n12152), .ZN(n16) );
  INV_X2 U59 ( .A(n466), .ZN(n12152) );
  INV_X4 U61 ( .A(n142), .ZN(instr_addr_o_6_) );
  OR2_X1 U63 ( .A1(n5041), .A2(n7346), .ZN(n4785) );
  INV_X1 U64 ( .A(instr_addr_i[18]), .ZN(n17) );
  AND2_X1 U67 ( .A1(n4234), .A2(n9842), .ZN(n4500) );
  NOR2_X1 U68 ( .A1(n5187), .A2(n4328), .ZN(n4331) );
  AND2_X1 U69 ( .A1(n4234), .A2(n11793), .ZN(n3952) );
  NAND2_X1 U70 ( .A1(instr_addr_o_11_), .A2(n1284), .ZN(n5607) );
  OR2_X1 U71 ( .A1(n3100), .A2(n7301), .ZN(n5387) );
  AND2_X1 U72 ( .A1(n4153), .A2(n6484), .ZN(n18) );
  INV_X2 U73 ( .A(n2739), .ZN(n206) );
  AND4_X1 U74 ( .A1(n3370), .A2(n3369), .A3(n3368), .A4(n3367), .ZN(n19) );
  INV_X2 U76 ( .A(n1431), .ZN(n5069) );
  AND3_X1 U77 ( .A1(n5333), .A2(n5331), .A3(n5332), .ZN(n5334) );
  AND4_X1 U78 ( .A1(n4678), .A2(n4677), .A3(n4676), .A4(n4675), .ZN(n4679) );
  INV_X1 U79 ( .A(n3531), .ZN(n5057) );
  NAND2_X1 U80 ( .A1(n5192), .A2(pmp_addr_i[372]), .ZN(n69) );
  INV_X2 U86 ( .A(n467), .ZN(n5293) );
  INV_X1 U88 ( .A(n5031), .ZN(n4596) );
  INV_X1 U89 ( .A(n5031), .ZN(n5280) );
  CLKBUF_X1 U90 ( .A(n12130), .Z(n12140) );
  INV_X2 U91 ( .A(n3876), .ZN(n5899) );
  INV_X1 U92 ( .A(n5031), .ZN(n20) );
  INV_X1 U93 ( .A(n9918), .ZN(n9860) );
  INV_X1 U95 ( .A(n9947), .ZN(n31) );
  INV_X2 U96 ( .A(data_addr_i[31]), .ZN(data_addr_o_31__BAR) );
  CLKBUF_X1 U97 ( .A(data_addr_i[25]), .Z(n11320) );
  BUF_X1 U99 ( .A(data_addr_i[18]), .Z(n10967) );
  CLKBUF_X1 U101 ( .A(data_addr_i[27]), .Z(n10746) );
  BUF_X2 U102 ( .A(data_addr_i[12]), .Z(data_addr_o_12_) );
  CLKBUF_X2 U104 ( .A(data_addr_i[14]), .Z(data_addr_o_14_) );
  INV_X2 U108 ( .A(n7923), .ZN(n23) );
  OR2_X2 U109 ( .A1(n471), .A2(pmp_cfg_i[60]), .ZN(n432) );
  AOI22_X1 U111 ( .A1(n49), .A2(n48), .B1(n4650), .B2(n47), .ZN(n46) );
  AOI21_X1 U112 ( .B1(n2382), .B2(n2381), .A(n2380), .ZN(n2383) );
  AOI21_X1 U113 ( .B1(n5139), .B2(n5138), .A(n5137), .ZN(n5140) );
  NAND4_X1 U114 ( .A1(n131), .A2(n2841), .A3(n133), .A4(n2860), .ZN(n2924) );
  AOI21_X1 U115 ( .B1(n4665), .B2(n4666), .A(n4664), .ZN(n50) );
  NOR2_X1 U116 ( .A1(n1768), .A2(n1767), .ZN(n85) );
  NOR2_X1 U117 ( .A1(n2864), .A2(n132), .ZN(n131) );
  INV_X1 U118 ( .A(n2107), .ZN(n2102) );
  INV_X1 U119 ( .A(n1861), .ZN(n1856) );
  NOR2_X1 U120 ( .A1(n588), .A2(n512), .ZN(n606) );
  INV_X1 U121 ( .A(n2748), .ZN(n94) );
  AND3_X1 U122 ( .A1(n4729), .A2(n124), .A3(n4728), .ZN(n123) );
  OAI211_X1 U123 ( .C1(n5048), .C2(n9842), .A(n3574), .B(n4514), .ZN(n3566) );
  OR2_X1 U125 ( .A1(n1537), .A2(n1486), .ZN(n1509) );
  OR2_X1 U126 ( .A1(n5633), .A2(n5634), .ZN(n57) );
  AOI22_X1 U127 ( .A1(n4388), .A2(n4398), .B1(n4602), .B2(pmp_addr_i[104]), 
        .ZN(n4400) );
  BUF_X1 U129 ( .A(n362), .Z(instr_addr_o_19_) );
  NAND2_X1 U130 ( .A1(n4498), .A2(n4497), .ZN(n4514) );
  AND2_X1 U131 ( .A1(n4726), .A2(n4727), .ZN(n125) );
  AOI22_X1 U132 ( .A1(n4088), .A2(n4098), .B1(n4602), .B2(pmp_addr_i[488]), 
        .ZN(n4100) );
  NOR2_X1 U133 ( .A1(n12179), .A2(n7651), .ZN(n3268) );
  INV_X1 U134 ( .A(n2441), .ZN(n3284) );
  OR2_X1 U135 ( .A1(n2467), .A2(n2441), .ZN(n2465) );
  NOR2_X1 U136 ( .A1(n1662), .A2(n1700), .ZN(n1693) );
  AND2_X1 U137 ( .A1(n2070), .A2(n66), .ZN(n65) );
  OAI21_X1 U138 ( .B1(n5048), .B2(pmp_addr_i[367]), .A(n3111), .ZN(n3113) );
  OR2_X1 U139 ( .A1(n1544), .A2(n1482), .ZN(n1537) );
  AND4_X1 U140 ( .A1(n5545), .A2(n5544), .A3(n5543), .A4(n5555), .ZN(n43) );
  INV_X1 U141 ( .A(n4475), .ZN(n82) );
  AND2_X1 U142 ( .A1(n616), .A2(n9940), .ZN(n4508) );
  INV_X2 U143 ( .A(n499), .ZN(n12265) );
  AND2_X1 U144 ( .A1(n3000), .A2(n10298), .ZN(n3014) );
  NOR2_X1 U145 ( .A1(n5187), .A2(n4529), .ZN(n4532) );
  OR2_X1 U146 ( .A1(n4147), .A2(pmp_addr_i[345]), .ZN(n61) );
  OR2_X1 U148 ( .A1(n5052), .A2(pmp_addr_i[73]), .ZN(n66) );
  OR2_X1 U149 ( .A1(n5094), .A2(pmp_addr_i[185]), .ZN(n64) );
  CLKBUF_X2 U150 ( .A(n5163), .Z(n4438) );
  NOR2_X1 U151 ( .A1(n5974), .A2(n7666), .ZN(n2441) );
  INV_X1 U152 ( .A(n2423), .ZN(n3298) );
  OR2_X1 U153 ( .A1(n616), .A2(pmp_addr_i[268]), .ZN(n1825) );
  OR2_X1 U157 ( .A1(n4658), .A2(pmp_addr_i[508]), .ZN(n4151) );
  BUF_X2 U158 ( .A(n5240), .Z(n149) );
  OR2_X1 U159 ( .A1(n3839), .A2(pmp_addr_i[227]), .ZN(n91) );
  OR2_X1 U161 ( .A1(n5250), .A2(n1285), .ZN(n5527) );
  AND2_X1 U162 ( .A1(n3819), .A2(n7296), .ZN(n360) );
  CLKBUF_X2 U163 ( .A(n937), .Z(instr_addr_o_13_) );
  INV_X1 U165 ( .A(n1131), .ZN(instr_addr_o_26_) );
  NOR2_X1 U167 ( .A1(n12152), .A2(n7656), .ZN(n2423) );
  INV_X1 U169 ( .A(instr_addr_i[23]), .ZN(n5086) );
  INV_X1 U171 ( .A(n467), .ZN(n6015) );
  INV_X1 U172 ( .A(instr_addr_i[5]), .ZN(n5031) );
  AND2_X1 U173 ( .A1(n11026), .A2(n106), .ZN(n11027) );
  CLKBUF_X1 U174 ( .A(data_addr_i[31]), .Z(n10662) );
  CLKBUF_X1 U176 ( .A(data_addr_i[23]), .Z(n10737) );
  INV_X1 U177 ( .A(n9941), .ZN(n11309) );
  CLKBUF_X1 U179 ( .A(data_addr_i[13]), .Z(data_addr_o_13_) );
  CLKBUF_X1 U180 ( .A(data_addr_i[18]), .Z(n11298) );
  INV_X1 U182 ( .A(n10494), .ZN(n29) );
  BUF_X4 U183 ( .A(data_addr_i[9]), .Z(data_addr_o_9_) );
  CLKBUF_X1 U184 ( .A(data_addr_i[13]), .Z(n6649) );
  OAI21_X2 U185 ( .B1(n11564), .B2(n625), .A(pmp_cfg_i[52]), .ZN(n4893) );
  CLKBUF_X1 U186 ( .A(data_addr_i[6]), .Z(n10953) );
  CLKBUF_X1 U187 ( .A(data_addr_i[6]), .Z(n10655) );
  INV_X1 U188 ( .A(data_addr_i[5]), .ZN(n11291) );
  CLKBUF_X1 U189 ( .A(data_addr_i[6]), .Z(n10358) );
  CLKBUF_X1 U190 ( .A(data_addr_i[6]), .Z(data_addr_o_6_) );
  NOR2_X1 U191 ( .A1(n2727), .A2(n2726), .ZN(n325) );
  NOR2_X1 U192 ( .A1(n11963), .A2(n3507), .ZN(n11947) );
  INV_X1 U193 ( .A(n10260), .ZN(n34) );
  CLKBUF_X1 U194 ( .A(data_addr_i[6]), .Z(n11331) );
  OAI21_X2 U196 ( .B1(n11510), .B2(n2716), .A(pmp_cfg_i[12]), .ZN(n4996) );
  INV_X1 U197 ( .A(data_addr_i[4]), .ZN(n12058) );
  NAND2_X1 U198 ( .A1(n5951), .A2(n5963), .ZN(n6011) );
  OR2_X1 U199 ( .A1(n1959), .A2(n6257), .ZN(n101) );
  INV_X1 U200 ( .A(data_addr_i[2]), .ZN(n10651) );
  NOR2_X1 U201 ( .A1(n11989), .A2(n3499), .ZN(n11992) );
  OAI21_X1 U202 ( .B1(n12041), .B2(n112), .A(n5948), .ZN(n5951) );
  OR4_X1 U203 ( .A1(n12041), .A2(n2996), .A3(n2992), .A4(n116), .ZN(n111) );
  OR3_X1 U204 ( .A1(n12041), .A2(n116), .A3(n2992), .ZN(n115) );
  NAND2_X1 U205 ( .A1(n217), .A2(n218), .ZN(n3476) );
  OR2_X1 U206 ( .A1(n5384), .A2(n1727), .ZN(n11050) );
  AOI21_X2 U208 ( .B1(n1911), .B2(n11155), .A(n6096), .ZN(n5663) );
  AND2_X1 U209 ( .A1(n7246), .A2(pmp_cfg_i[58]), .ZN(n143) );
  INV_X1 U211 ( .A(n2219), .ZN(n6935) );
  AND2_X1 U212 ( .A1(n119), .A2(n117), .ZN(n12018) );
  NOR2_X1 U213 ( .A1(n4891), .A2(n611), .ZN(n4842) );
  INV_X1 U214 ( .A(n4892), .ZN(n878) );
  NOR2_X1 U215 ( .A1(n11062), .A2(n1741), .ZN(n11068) );
  NOR2_X1 U216 ( .A1(n11975), .A2(n3497), .ZN(n3511) );
  NOR3_X1 U217 ( .A1(n5933), .A2(n2959), .A3(n3127), .ZN(n119) );
  NOR2_X2 U218 ( .A1(n5283), .A2(pmp_cfg_i[44]), .ZN(n161) );
  OR2_X2 U219 ( .A1(n2227), .A2(pmp_cfg_i[76]), .ZN(n2219) );
  INV_X2 U220 ( .A(n156), .ZN(n35) );
  NOR2_X2 U221 ( .A1(n11659), .A2(pmp_cfg_i[84]), .ZN(n9329) );
  NOR2_X1 U222 ( .A1(n2394), .A2(pmp_cfg_i[116]), .ZN(n7923) );
  OR2_X1 U223 ( .A1(n663), .A2(pmp_cfg_i[52]), .ZN(n4892) );
  INV_X2 U224 ( .A(n160), .ZN(n36) );
  NOR2_X1 U225 ( .A1(n4194), .A2(pmp_cfg_i[28]), .ZN(n7551) );
  NOR2_X1 U226 ( .A1(n1948), .A2(pmp_cfg_i[19]), .ZN(n6096) );
  AND3_X1 U227 ( .A1(pmp_addr_i[427]), .A2(pmp_addr_i[426]), .A3(
        pmp_addr_i[428]), .ZN(n60) );
  INV_X1 U228 ( .A(pmp_addr_i[365]), .ZN(n116) );
  INV_X1 U229 ( .A(pmp_addr_i[291]), .ZN(n89) );
  NAND4_X1 U230 ( .A1(n37), .A2(n53), .A3(n4619), .A4(n4620), .ZN(n52) );
  OAI211_X1 U231 ( .C1(n4610), .C2(n4611), .A(n4618), .B(n4609), .ZN(n37) );
  NAND4_X1 U232 ( .A1(n3186), .A2(n38), .A3(n3174), .A4(n3175), .ZN(n3202) );
  OAI211_X1 U233 ( .C1(n3172), .C2(n3173), .A(n69), .B(n68), .ZN(n38) );
  NAND3_X1 U234 ( .A1(n39), .A2(n1347), .A3(n1348), .ZN(n1362) );
  NAND2_X1 U235 ( .A1(n1338), .A2(n1337), .ZN(n39) );
  NAND3_X1 U236 ( .A1(n40), .A2(n83), .A3(n82), .ZN(n277) );
  OAI21_X1 U237 ( .B1(n4472), .B2(n4471), .A(n4470), .ZN(n40) );
  NOR2_X1 U238 ( .A1(n41), .A2(n2067), .ZN(n2064) );
  NAND2_X1 U239 ( .A1(n65), .A2(n2071), .ZN(n41) );
  NAND2_X1 U240 ( .A1(n2073), .A2(n2057), .ZN(n2075) );
  NAND4_X1 U241 ( .A1(n42), .A2(n4436), .A3(n4426), .A4(n4427), .ZN(n4450) );
  OAI21_X1 U242 ( .B1(n4425), .B2(n4424), .A(n4423), .ZN(n42) );
  NAND4_X1 U243 ( .A1(n5556), .A2(n43), .A3(n5554), .A4(n5542), .ZN(n5565) );
  OAI21_X1 U244 ( .B1(n4638), .B2(n4637), .A(n4636), .ZN(n48) );
  AND2_X1 U245 ( .A1(n5313), .A2(pmp_addr_i[433]), .ZN(n4633) );
  OAI21_X1 U246 ( .B1(n3961), .B2(n4698), .A(n45), .ZN(n3962) );
  NAND3_X1 U247 ( .A1(n3956), .A2(n44), .A3(n3966), .ZN(n4704) );
  AND2_X1 U248 ( .A1(n4703), .A2(n45), .ZN(n44) );
  NAND2_X1 U249 ( .A1(n206), .A2(n4733), .ZN(n45) );
  OAI211_X1 U250 ( .C1(n51), .C2(n4630), .A(n50), .B(n46), .ZN(n4667) );
  NOR2_X1 U251 ( .A1(n291), .A2(n4640), .ZN(n47) );
  NOR3_X1 U252 ( .A1(n291), .A2(n293), .A3(n290), .ZN(n49) );
  AND2_X1 U253 ( .A1(n52), .A2(n54), .ZN(n51) );
  NAND2_X1 U254 ( .A1(n4618), .A2(n4617), .ZN(n53) );
  AOI21_X1 U255 ( .B1(n4619), .B2(n56), .A(n55), .ZN(n54) );
  OAI21_X1 U256 ( .B1(n4592), .B2(n4593), .A(n4591), .ZN(n55) );
  OAI21_X1 U257 ( .B1(n4586), .B2(n4614), .A(n4585), .ZN(n56) );
  NAND2_X1 U258 ( .A1(n4615), .A2(n4616), .ZN(n4617) );
  NOR2_X1 U260 ( .A1(n5635), .A2(n57), .ZN(n5655) );
  OAI21_X1 U261 ( .B1(n5972), .B2(n58), .A(n5971), .ZN(n6038) );
  NAND3_X1 U263 ( .A1(n242), .A2(n4453), .A3(n241), .ZN(n5021) );
  AND2_X1 U264 ( .A1(n3846), .A2(pmp_addr_i[103]), .ZN(n4388) );
  INV_X2 U265 ( .A(n1431), .ZN(n3934) );
  NAND2_X1 U267 ( .A1(n9866), .A2(n9781), .ZN(n9868) );
  NAND4_X1 U268 ( .A1(n59), .A2(n941), .A3(n908), .A4(n940), .ZN(n936) );
  OR2_X1 U269 ( .A1(n915), .A2(n895), .ZN(n59) );
  NAND2_X1 U270 ( .A1(n11992), .A2(n60), .ZN(n3535) );
  NAND2_X1 U271 ( .A1(n1843), .A2(n1858), .ZN(n1861) );
  NAND3_X1 U272 ( .A1(n9912), .A2(n9911), .A3(n9913), .ZN(n9997) );
  NAND3_X1 U273 ( .A1(n1124), .A2(n1116), .A3(n61), .ZN(n1056) );
  NAND2_X1 U274 ( .A1(instr_addr_o_28_), .A2(n3047), .ZN(n1116) );
  INV_X2 U275 ( .A(n499), .ZN(n12156) );
  NAND2_X1 U276 ( .A1(n62), .A2(n3801), .ZN(n179) );
  OAI21_X1 U277 ( .B1(n181), .B2(n180), .A(n3800), .ZN(n62) );
  AND2_X1 U278 ( .A1(n5052), .A2(n8517), .ZN(n3442) );
  BUF_X2 U281 ( .A(n1632), .Z(n4658) );
  AND2_X1 U283 ( .A1(n1935), .A2(n1937), .ZN(n63) );
  NAND2_X1 U284 ( .A1(n270), .A2(n3567), .ZN(n99) );
  NAND3_X1 U286 ( .A1(n5113), .A2(n5122), .A3(n64), .ZN(n5095) );
  NAND2_X1 U287 ( .A1(n4901), .A2(n5093), .ZN(n5113) );
  NAND4_X1 U288 ( .A1(n5450), .A2(n5453), .A3(n5451), .A4(n5452), .ZN(n5454)
         );
  NAND2_X1 U289 ( .A1(n12203), .A2(n6875), .ZN(n5450) );
  INV_X2 U290 ( .A(n3876), .ZN(n3836) );
  INV_X2 U292 ( .A(n212), .ZN(n5262) );
  INV_X2 U293 ( .A(n511), .ZN(n6018) );
  NAND2_X1 U294 ( .A1(n5031), .A2(n9980), .ZN(n83) );
  INV_X1 U295 ( .A(n2901), .ZN(n2913) );
  NAND2_X1 U296 ( .A1(n2797), .A2(n2807), .ZN(n307) );
  NOR3_X1 U297 ( .A1(n4986), .A2(n4987), .A3(n4985), .ZN(n67) );
  NAND3_X1 U298 ( .A1(n4161), .A2(n4160), .A3(n4159), .ZN(n4162) );
  NAND2_X1 U299 ( .A1(n3170), .A2(n3171), .ZN(n68) );
  BUF_X2 U301 ( .A(n5041), .Z(n4602) );
  NAND3_X1 U302 ( .A1(n7552), .A2(n7553), .A3(n7551), .ZN(n7618) );
  NAND2_X1 U303 ( .A1(n3406), .A2(n97), .ZN(n76) );
  OAI211_X1 U304 ( .C1(n7493), .C2(n7492), .A(n71), .B(n70), .ZN(n7494) );
  NAND2_X1 U305 ( .A1(n7490), .A2(n7491), .ZN(n70) );
  INV_X1 U306 ( .A(n7489), .ZN(n71) );
  OAI211_X1 U307 ( .C1(n1307), .C2(n1306), .A(n1304), .B(n1305), .ZN(n72) );
  NOR2_X1 U309 ( .A1(n3757), .A2(n73), .ZN(n3869) );
  NAND2_X1 U311 ( .A1(n4435), .A2(n4436), .ZN(n4449) );
  NAND2_X1 U313 ( .A1(n74), .A2(n177), .ZN(n1280) );
  AND3_X1 U314 ( .A1(n1252), .A2(n1261), .A3(n1159), .ZN(n74) );
  NAND4_X1 U315 ( .A1(n5334), .A2(n5345), .A3(n75), .A4(n175), .ZN(n5363) );
  INV_X1 U316 ( .A(n5335), .ZN(n75) );
  INV_X1 U317 ( .A(n5667), .ZN(n103) );
  OAI21_X1 U318 ( .B1(n3408), .B2(n3407), .A(n76), .ZN(n3757) );
  NAND3_X1 U319 ( .A1(n19), .A2(n3379), .A3(n77), .ZN(n3404) );
  NOR2_X1 U320 ( .A1(n3371), .A2(n78), .ZN(n77) );
  NAND2_X1 U321 ( .A1(n3378), .A2(n3380), .ZN(n78) );
  NAND3_X1 U322 ( .A1(n195), .A2(n4443), .A3(n196), .ZN(n4445) );
  NAND3_X1 U323 ( .A1(n4165), .A2(n4166), .A3(n4164), .ZN(n5022) );
  NAND3_X1 U324 ( .A1(n610), .A2(n79), .A3(n143), .ZN(n1407) );
  BUF_X2 U326 ( .A(n537), .Z(n1431) );
  OR2_X1 U327 ( .A1(n1431), .A2(n7325), .ZN(n4765) );
  NOR2_X1 U328 ( .A1(n80), .A2(n5012), .ZN(n234) );
  NAND4_X1 U329 ( .A1(n5006), .A2(n5007), .A3(n5004), .A4(n5005), .ZN(n80) );
  INV_X2 U331 ( .A(n3290), .ZN(instr_addr_o_20_) );
  NAND2_X1 U333 ( .A1(n86), .A2(n85), .ZN(n84) );
  NAND2_X1 U334 ( .A1(n1769), .A2(n1770), .ZN(n86) );
  NAND4_X1 U335 ( .A1(n564), .A2(n566), .A3(n567), .A4(n565), .ZN(n87) );
  NAND3_X1 U336 ( .A1(n2316), .A2(n2317), .A3(n88), .ZN(n2320) );
  NAND2_X1 U337 ( .A1(n4596), .A2(n89), .ZN(n88) );
  NAND3_X1 U338 ( .A1(n90), .A2(n555), .A3(n556), .ZN(n558) );
  NAND3_X1 U339 ( .A1(n553), .A2(n554), .A3(n91), .ZN(n90) );
  AND4_X2 U340 ( .A1(n1406), .A2(n1407), .A3(n1405), .A4(n1404), .ZN(n12135)
         );
  OAI22_X1 U341 ( .A1(n332), .A2(n2930), .B1(n92), .B2(n2929), .ZN(n12131) );
  AOI21_X1 U342 ( .B1(n305), .B2(n306), .A(n170), .ZN(n92) );
  NAND2_X1 U343 ( .A1(n93), .A2(n2747), .ZN(n2757) );
  OAI21_X1 U344 ( .B1(n2746), .B2(n2745), .A(n94), .ZN(n93) );
  AND2_X1 U345 ( .A1(n2733), .A2(n8208), .ZN(n2743) );
  OR2_X1 U347 ( .A1(n3846), .A2(n9801), .ZN(n4484) );
  NAND3_X1 U348 ( .A1(n4155), .A2(n4154), .A3(n18), .ZN(n4156) );
  NAND2_X1 U349 ( .A1(n2895), .A2(n2898), .ZN(n2901) );
  NAND2_X1 U350 ( .A1(n95), .A2(n4832), .ZN(n5017) );
  OAI21_X1 U353 ( .B1(n990), .B2(n989), .A(n988), .ZN(n96) );
  AND2_X1 U354 ( .A1(n3000), .A2(n9199), .ZN(n943) );
  OAI22_X1 U355 ( .A1(n3404), .A2(n3405), .B1(n3403), .B2(n3402), .ZN(n97) );
  NAND2_X1 U356 ( .A1(n2092), .A2(n2104), .ZN(n2107) );
  NAND3_X1 U357 ( .A1(n1337), .A2(n309), .A3(n311), .ZN(n258) );
  NAND4_X1 U359 ( .A1(n4504), .A2(n4484), .A3(n4506), .A4(n4473), .ZN(n98) );
  OAI21_X1 U361 ( .B1(n3569), .B2(n3568), .A(n99), .ZN(n3638) );
  NAND2_X1 U362 ( .A1(n409), .A2(n410), .ZN(n412) );
  NAND3_X1 U363 ( .A1(n2479), .A2(n2477), .A3(n2478), .ZN(n247) );
  BUF_X4 U364 ( .A(instr_addr_i[23]), .Z(n5208) );
  NAND3_X1 U365 ( .A1(n100), .A2(n1960), .A3(n5648), .ZN(n1961) );
  NAND2_X1 U366 ( .A1(n1958), .A2(n101), .ZN(n100) );
  OAI21_X1 U367 ( .B1(n2116), .B2(n102), .A(n2115), .ZN(n2117) );
  AOI22_X1 U368 ( .A1(n2111), .A2(n2112), .B1(pmp_addr_i[86]), .B2(n2580), 
        .ZN(n102) );
  AND2_X1 U369 ( .A1(n5313), .A2(pmp_addr_i[113]), .ZN(n4420) );
  BUF_X2 U370 ( .A(n372), .Z(n3045) );
  NAND2_X1 U371 ( .A1(n103), .A2(n5646), .ZN(n1920) );
  NAND2_X1 U372 ( .A1(n104), .A2(n5646), .ZN(n204) );
  INV_X1 U374 ( .A(n5720), .ZN(n104) );
  NOR2_X1 U375 ( .A1(n105), .A2(n10227), .ZN(n10228) );
  OAI21_X1 U376 ( .B1(n10251), .B2(n105), .A(n10250), .ZN(n10252) );
  NAND2_X1 U377 ( .A1(n10226), .A2(n10249), .ZN(n105) );
  NAND2_X1 U378 ( .A1(n108), .A2(n107), .ZN(n106) );
  INV_X1 U379 ( .A(n12054), .ZN(n107) );
  NAND2_X1 U380 ( .A1(n110), .A2(n109), .ZN(n108) );
  NAND2_X1 U381 ( .A1(n12007), .A2(n10331), .ZN(n109) );
  NAND3_X1 U382 ( .A1(n10257), .A2(n10256), .A3(n10332), .ZN(n110) );
  NAND2_X1 U383 ( .A1(n114), .A2(n113), .ZN(n112) );
  NOR2_X1 U384 ( .A1(n2996), .A2(n2997), .ZN(n113) );
  NOR2_X1 U385 ( .A1(n116), .A2(n2992), .ZN(n114) );
  NOR2_X1 U386 ( .A1(n12041), .A2(n2992), .ZN(n12024) );
  NOR3_X1 U387 ( .A1(n12042), .A2(n2990), .A3(n2950), .ZN(n117) );
  NAND2_X1 U388 ( .A1(n119), .A2(n120), .ZN(n12014) );
  NOR2_X1 U389 ( .A1(n12042), .A2(n2950), .ZN(n120) );
  NOR2_X1 U390 ( .A1(n5933), .A2(n2950), .ZN(n12021) );
  NAND2_X1 U391 ( .A1(n120), .A2(n118), .ZN(n12009) );
  NOR2_X1 U392 ( .A1(n5933), .A2(n2959), .ZN(n118) );
  OAI211_X1 U393 ( .C1(n127), .C2(n4739), .A(n4738), .B(n121), .ZN(n5018) );
  NOR2_X1 U394 ( .A1(n122), .A2(n4737), .ZN(n121) );
  NAND4_X1 U395 ( .A1(n126), .A2(n125), .A3(n4736), .A4(n123), .ZN(n122) );
  INV_X1 U396 ( .A(n4735), .ZN(n124) );
  INV_X1 U397 ( .A(n4734), .ZN(n126) );
  INV_X1 U398 ( .A(n4680), .ZN(n129) );
  NOR2_X1 U399 ( .A1(n130), .A2(n2864), .ZN(n2858) );
  NAND3_X1 U400 ( .A1(n133), .A2(n2866), .A3(n2860), .ZN(n130) );
  NAND2_X1 U401 ( .A1(n4901), .A2(n2767), .ZN(n2860) );
  NAND3_X1 U402 ( .A1(n2850), .A2(n2866), .A3(n2840), .ZN(n132) );
  NAND2_X1 U403 ( .A1(n134), .A2(n2769), .ZN(n133) );
  INV_X1 U404 ( .A(n4147), .ZN(n134) );
  INV_X1 U405 ( .A(n3992), .ZN(n136) );
  INV_X1 U406 ( .A(n3992), .ZN(n137) );
  INV_X1 U407 ( .A(n5163), .ZN(n138) );
  AND3_X1 U408 ( .A1(n3165), .A2(n3164), .A3(n3194), .ZN(n139) );
  INV_X2 U409 ( .A(n1026), .ZN(n5985) );
  INV_X1 U412 ( .A(n4234), .ZN(n4069) );
  OR2_X1 U413 ( .A1(n12211), .A2(pmp_addr_i[509]), .ZN(n4152) );
  AND2_X1 U414 ( .A1(n376), .A2(n6637), .ZN(n4041) );
  INV_X1 U415 ( .A(instr_addr_i[6]), .ZN(n142) );
  INV_X2 U416 ( .A(instr_addr_i[20]), .ZN(n3290) );
  INV_X2 U417 ( .A(n3290), .ZN(n4802) );
  BUF_X2 U418 ( .A(n17), .Z(instr_addr_o_18__BAR) );
  BUF_X2 U420 ( .A(instr_addr_o_18__BAR), .Z(n1922) );
  BUF_X2 U422 ( .A(n5979), .Z(n146) );
  INV_X2 U423 ( .A(n2103), .ZN(n5181) );
  INV_X2 U425 ( .A(n2707), .ZN(instr_addr_o_8_) );
  INV_X2 U426 ( .A(n2707), .ZN(n5342) );
  INV_X1 U431 ( .A(n543), .ZN(n5996) );
  BUF_X2 U432 ( .A(instr_addr_i[13]), .Z(n5997) );
  OR2_X1 U433 ( .A1(n376), .A2(pmp_addr_i[124]), .ZN(n4441) );
  AND2_X1 U434 ( .A1(n10614), .A2(n597), .ZN(n7097) );
  NOR2_X1 U435 ( .A1(n6027), .A2(n2776), .ZN(n2800) );
  OR2_X1 U436 ( .A1(n4406), .A2(pmp_addr_i[123]), .ZN(n278) );
  INV_X1 U437 ( .A(n3209), .ZN(n3253) );
  OR2_X1 U438 ( .A1(n4623), .A2(pmp_addr_i[379]), .ZN(n263) );
  AND2_X1 U439 ( .A1(n4658), .A2(n8055), .ZN(n180) );
  AND2_X1 U440 ( .A1(n3799), .A2(n182), .ZN(n181) );
  INV_X1 U441 ( .A(n3800), .ZN(n184) );
  AND3_X1 U442 ( .A1(n5812), .A2(n5808), .A3(n5811), .ZN(n200) );
  INV_X1 U443 ( .A(n5893), .ZN(n280) );
  INV_X1 U444 ( .A(n5903), .ZN(n283) );
  INV_X1 U445 ( .A(n5833), .ZN(n285) );
  AND2_X1 U446 ( .A1(n2733), .A2(n9204), .ZN(n3321) );
  AND2_X1 U447 ( .A1(n5086), .A2(pmp_addr_i[437]), .ZN(n4642) );
  OR2_X1 U448 ( .A1(n312), .A2(n1395), .ZN(n1378) );
  AND3_X1 U449 ( .A1(n675), .A2(n4833), .A3(n676), .ZN(n253) );
  NOR2_X1 U450 ( .A1(n426), .A2(n418), .ZN(n448) );
  OR2_X1 U451 ( .A1(n1972), .A2(n2019), .ZN(n1993) );
  BUF_X2 U452 ( .A(n362), .Z(n3793) );
  OR2_X1 U453 ( .A1(n10614), .A2(n597), .ZN(n7095) );
  AND2_X1 U454 ( .A1(n5023), .A2(pmp_addr_i[164]), .ZN(n246) );
  INV_X1 U455 ( .A(pmp_cfg_i[99]), .ZN(n1454) );
  OR2_X1 U456 ( .A1(instr_addr_o_18__BAR), .A2(n9939), .ZN(n4517) );
  AND2_X1 U457 ( .A1(n3000), .A2(n7571), .ZN(n4255) );
  AND2_X1 U458 ( .A1(n5023), .A2(n7333), .ZN(n4183) );
  AND2_X1 U459 ( .A1(n5000), .A2(n11510), .ZN(n236) );
  OR2_X1 U460 ( .A1(n616), .A2(n9940), .ZN(n4506) );
  OR2_X1 U461 ( .A1(n4200), .A2(n10830), .ZN(n5889) );
  INV_X1 U462 ( .A(n5889), .ZN(n286) );
  NOR2_X1 U463 ( .A1(n213), .A2(n8229), .ZN(n4965) );
  NOR2_X1 U464 ( .A1(n12152), .A2(n327), .ZN(n4958) );
  INV_X1 U465 ( .A(n4641), .ZN(n293) );
  OR2_X1 U466 ( .A1(n4651), .A2(n4639), .ZN(n291) );
  AND3_X1 U467 ( .A1(n277), .A2(n4473), .A3(n276), .ZN(n4491) );
  OR2_X1 U468 ( .A1(n4474), .A2(n4475), .ZN(n276) );
  OR2_X1 U469 ( .A1(instr_addr_o_18__BAR), .A2(n6648), .ZN(n3968) );
  OAI21_X1 U470 ( .B1(n4658), .B2(n197), .A(n192), .ZN(n196) );
  INV_X1 U471 ( .A(n193), .ZN(n192) );
  OAI22_X1 U472 ( .A1(n4778), .A2(n11713), .B1(n4779), .B2(n11722), .ZN(n235)
         );
  NOR3_X1 U473 ( .A1(n3322), .A2(n3321), .A3(n3320), .ZN(n314) );
  AND2_X1 U474 ( .A1(n5163), .A2(n10266), .ZN(n3080) );
  AND2_X1 U475 ( .A1(n1269), .A2(n8034), .ZN(n225) );
  AND2_X1 U476 ( .A1(n5947), .A2(n111), .ZN(n239) );
  OAI21_X1 U477 ( .B1(n5895), .B2(n11362), .A(n287), .ZN(n5877) );
  NOR2_X1 U478 ( .A1(n5873), .A2(n10806), .ZN(n288) );
  NOR2_X1 U479 ( .A1(n5847), .A2(n294), .ZN(n5853) );
  AND2_X1 U480 ( .A1(n5096), .A2(n5139), .ZN(n264) );
  AND2_X1 U481 ( .A1(n2896), .A2(n11681), .ZN(n3320) );
  INV_X1 U482 ( .A(n2800), .ZN(n178) );
  NOR2_X1 U483 ( .A1(n4965), .A2(n4949), .ZN(n2711) );
  INV_X1 U485 ( .A(n4129), .ZN(n4124) );
  NOR2_X2 U486 ( .A1(n3895), .A2(pmp_cfg_i[124]), .ZN(n6624) );
  NOR3_X1 U487 ( .A1(n4418), .A2(n4417), .A3(n4437), .ZN(n4436) );
  INV_X1 U488 ( .A(n4424), .ZN(n4411) );
  OR2_X1 U489 ( .A1(n3237), .A2(n240), .ZN(n3245) );
  INV_X1 U490 ( .A(n2968), .ZN(n269) );
  NOR2_X1 U491 ( .A1(n3798), .A2(n184), .ZN(n183) );
  AND2_X1 U492 ( .A1(n5698), .A2(n5697), .ZN(n229) );
  NOR2_X1 U493 ( .A1(n281), .A2(n280), .ZN(n279) );
  AND2_X1 U494 ( .A1(n5070), .A2(pmp_addr_i[74]), .ZN(n231) );
  INV_X1 U495 ( .A(n1767), .ZN(n1745) );
  NOR2_X1 U496 ( .A1(n5799), .A2(n5815), .ZN(n1775) );
  INV_X1 U497 ( .A(n1715), .ZN(n1677) );
  INV_X1 U498 ( .A(n1509), .ZN(n1508) );
  AND2_X1 U499 ( .A1(n2463), .A2(n2471), .ZN(n2464) );
  AOI21_X1 U500 ( .B1(n2470), .B2(n2469), .A(n2468), .ZN(n2478) );
  NOR3_X1 U501 ( .A1(n2892), .A2(n2908), .A3(n164), .ZN(n296) );
  AND4_X1 U502 ( .A1(n2658), .A2(n2649), .A3(n2640), .A4(n2635), .ZN(n274) );
  NOR2_X1 U503 ( .A1(n2637), .A2(n2654), .ZN(n275) );
  AND2_X1 U504 ( .A1(n7551), .A2(pmp_cfg_i[26]), .ZN(n241) );
  AOI21_X1 U505 ( .B1(n3198), .B2(n3199), .A(n228), .ZN(n3200) );
  AND2_X1 U506 ( .A1(n10256), .A2(pmp_cfg_i[90]), .ZN(n254) );
  NOR3_X1 U507 ( .A1(n5364), .A2(n271), .A3(n5373), .ZN(n5412) );
  NOR2_X1 U508 ( .A1(n1056), .A2(n1121), .ZN(n1141) );
  AND2_X1 U509 ( .A1(n1377), .A2(n255), .ZN(n1361) );
  AND2_X1 U510 ( .A1(n1360), .A2(n1376), .ZN(n255) );
  INV_X1 U511 ( .A(n1378), .ZN(n1377) );
  AND3_X1 U512 ( .A1(n678), .A2(n319), .A3(n252), .ZN(n738) );
  OR2_X1 U513 ( .A1(n489), .A2(n488), .ZN(n490) );
  INV_X1 U514 ( .A(n1993), .ZN(n1992) );
  OR2_X1 U515 ( .A1(n2338), .A2(n2337), .ZN(n2347) );
  AND2_X1 U516 ( .A1(n9584), .A2(pmp_cfg_i[34]), .ZN(n226) );
  AND2_X1 U517 ( .A1(n878), .A2(pmp_cfg_i[50]), .ZN(n272) );
  CLKBUF_X1 U519 ( .A(n12133), .Z(n6047) );
  INV_X1 U520 ( .A(instr_addr_i[30]), .ZN(n1632) );
  BUF_X2 U522 ( .A(data_addr_i[23]), .Z(n10898) );
  INV_X1 U523 ( .A(n1150), .ZN(n9584) );
  OR2_X2 U524 ( .A1(n1215), .A2(pmp_cfg_i[36]), .ZN(n1150) );
  NOR2_X1 U525 ( .A1(n1742), .A2(pmp_cfg_i[68]), .ZN(n156) );
  INV_X2 U526 ( .A(n3819), .ZN(instr_addr_o_21_) );
  INV_X1 U527 ( .A(n3984), .ZN(n5183) );
  AND2_X1 U528 ( .A1(n4179), .A2(n4178), .ZN(n157) );
  NAND2_X1 U529 ( .A1(n3665), .A2(pmp_addr_i[7]), .ZN(n158) );
  NAND2_X1 U530 ( .A1(n3679), .A2(pmp_addr_i[6]), .ZN(n159) );
  OR2_X1 U531 ( .A1(n2695), .A2(pmp_cfg_i[12]), .ZN(n160) );
  AND2_X1 U533 ( .A1(n9911), .A2(pmp_cfg_i[106]), .ZN(n162) );
  AND3_X1 U534 ( .A1(n11420), .A2(n1419), .A3(n1415), .ZN(n163) );
  AND2_X1 U535 ( .A1(instr_addr_o_11_), .A2(n4981), .ZN(n164) );
  AND4_X1 U536 ( .A1(n5825), .A2(n5824), .A3(n5823), .A4(n5822), .ZN(n165) );
  AND4_X1 U537 ( .A1(n5716), .A2(n5715), .A3(n5714), .A4(n5713), .ZN(n166) );
  AND4_X1 U538 ( .A1(n1627), .A2(n1618), .A3(n1626), .A4(n1604), .ZN(n167) );
  AND2_X1 U539 ( .A1(n156), .A2(pmp_cfg_i[66]), .ZN(n168) );
  NOR2_X1 U541 ( .A1(n773), .A2(n702), .ZN(n169) );
  AND2_X1 U542 ( .A1(n2824), .A2(n2823), .ZN(n170) );
  AND2_X1 U543 ( .A1(n2151), .A2(n2175), .ZN(n171) );
  OR2_X1 U544 ( .A1(n5069), .A2(n7266), .ZN(n172) );
  OR2_X1 U545 ( .A1(n12202), .A2(n5261), .ZN(n173) );
  AND2_X1 U546 ( .A1(n3195), .A2(n10111), .ZN(n174) );
  AND2_X1 U547 ( .A1(n5343), .A2(n5344), .ZN(n175) );
  OR2_X1 U548 ( .A1(pmp_addr_i[125]), .A2(n197), .ZN(n176) );
  AOI21_X1 U549 ( .B1(n1260), .B2(n177), .A(n1259), .ZN(n1263) );
  NAND3_X1 U551 ( .A1(n2806), .A2(n2783), .A3(n178), .ZN(n2784) );
  AND2_X1 U553 ( .A1(n4406), .A2(n8054), .ZN(n182) );
  NAND2_X1 U554 ( .A1(n186), .A2(n3797), .ZN(n185) );
  NAND3_X1 U555 ( .A1(n3796), .A2(n4147), .A3(n8049), .ZN(n186) );
  INV_X1 U556 ( .A(n187), .ZN(n188) );
  OAI21_X1 U557 ( .B1(n1054), .B2(n1069), .A(n1053), .ZN(n187) );
  NAND2_X1 U559 ( .A1(n1070), .A2(n1071), .ZN(n189) );
  NAND2_X1 U561 ( .A1(n191), .A2(n4407), .ZN(n4442) );
  INV_X1 U562 ( .A(n3295), .ZN(n191) );
  OAI22_X1 U563 ( .A1(n12211), .A2(n176), .B1(n197), .B2(pmp_addr_i[124]), 
        .ZN(n193) );
  INV_X2 U564 ( .A(n376), .ZN(n12161) );
  NAND4_X1 U565 ( .A1(n4656), .A2(pmp_addr_i[123]), .A3(n4442), .A4(n4441), 
        .ZN(n195) );
  INV_X1 U566 ( .A(n4444), .ZN(n197) );
  NAND3_X1 U567 ( .A1(n448), .A2(n172), .A3(n447), .ZN(n5364) );
  NAND4_X1 U568 ( .A1(n5809), .A2(n5817), .A3(n5807), .A4(n5816), .ZN(n201) );
  NOR2_X1 U569 ( .A1(n201), .A2(n199), .ZN(n198) );
  NAND2_X1 U570 ( .A1(n200), .A2(n5813), .ZN(n199) );
  AND2_X1 U571 ( .A1(n2896), .A2(n7320), .ZN(n4250) );
  AND2_X1 U572 ( .A1(n1014), .A2(n333), .ZN(n202) );
  AND2_X1 U573 ( .A1(n5023), .A2(n10814), .ZN(n5837) );
  OR2_X1 U575 ( .A1(n4623), .A2(n6664), .ZN(n4040) );
  AND2_X1 U576 ( .A1(n3846), .A2(n7819), .ZN(n3260) );
  AND2_X1 U577 ( .A1(n4652), .A2(pmp_addr_i[121]), .ZN(n299) );
  AND2_X1 U578 ( .A1(n12203), .A2(n11194), .ZN(n203) );
  NAND2_X1 U579 ( .A1(n204), .A2(n5715), .ZN(n1925) );
  BUF_X1 U580 ( .A(n2339), .Z(n3025) );
  NOR2_X1 U582 ( .A1(n5047), .A2(n6557), .ZN(n3969) );
  INV_X2 U583 ( .A(n3894), .ZN(n205) );
  INV_X1 U585 ( .A(instr_addr_i[15]), .ZN(n207) );
  NAND3_X1 U587 ( .A1(n1894), .A2(n1893), .A3(n168), .ZN(n2389) );
  INV_X2 U588 ( .A(n1131), .ZN(n210) );
  AND2_X1 U589 ( .A1(n4234), .A2(n9045), .ZN(n3322) );
  NOR2_X2 U591 ( .A1(n3536), .A2(pmp_cfg_i[108]), .ZN(n9911) );
  OR2_X1 U592 ( .A1(n511), .A2(pmp_addr_i[445]), .ZN(n4659) );
  INV_X2 U594 ( .A(n3041), .ZN(n5149) );
  OR2_X1 U595 ( .A1(n5094), .A2(pmp_addr_i[441]), .ZN(n292) );
  OR2_X1 U596 ( .A1(n5094), .A2(pmp_addr_i[153]), .ZN(n313) );
  OR2_X1 U597 ( .A1(n5094), .A2(pmp_addr_i[121]), .ZN(n298) );
  OR2_X1 U598 ( .A1(n5094), .A2(pmp_addr_i[377]), .ZN(n266) );
  INV_X1 U599 ( .A(instr_addr_i[10]), .ZN(n212) );
  INV_X1 U600 ( .A(n5041), .ZN(n214) );
  INV_X2 U601 ( .A(n3275), .ZN(n6028) );
  AND3_X1 U602 ( .A1(n2912), .A2(n2895), .A3(n2904), .ZN(n297) );
  OAI21_X1 U603 ( .B1(pmp_cfg_i[43]), .B2(n5255), .A(n11381), .ZN(n215) );
  INV_X1 U605 ( .A(n1454), .ZN(n219) );
  INV_X1 U606 ( .A(pmp_cfg_i[100]), .ZN(n220) );
  NAND2_X1 U607 ( .A1(n219), .A2(n220), .ZN(n217) );
  NAND2_X1 U608 ( .A1(n219), .A2(n163), .ZN(n218) );
  INV_X1 U610 ( .A(n4234), .ZN(n5062) );
  NOR2_X1 U611 ( .A1(n1553), .A2(n1552), .ZN(n223) );
  OAI21_X1 U612 ( .B1(n224), .B2(n3810), .A(n3809), .ZN(n3811) );
  AOI21_X1 U613 ( .B1(n3803), .B2(n3804), .A(n225), .ZN(n224) );
  BUF_X2 U614 ( .A(n937), .Z(n4061) );
  INV_X1 U615 ( .A(n2214), .ZN(n227) );
  NAND3_X1 U616 ( .A1(n2183), .A2(n2184), .A3(n171), .ZN(n2214) );
  NAND3_X1 U617 ( .A1(n3197), .A2(n3196), .A3(n174), .ZN(n228) );
  AND2_X1 U618 ( .A1(n4234), .A2(pmp_addr_i[495]), .ZN(n4070) );
  AND2_X1 U619 ( .A1(n1438), .A2(n1468), .ZN(n259) );
  AOI21_X1 U620 ( .B1(n203), .B2(n11193), .A(n229), .ZN(n5708) );
  OAI21_X1 U622 ( .B1(n1362), .B2(n1363), .A(n1361), .ZN(n230) );
  AOI21_X1 U623 ( .B1(n2069), .B2(n2070), .A(n231), .ZN(n2076) );
  NAND4_X1 U624 ( .A1(n233), .A2(n2136), .A3(n6376), .A4(pmp_cfg_i[18]), .ZN(
        n2388) );
  OR2_X1 U625 ( .A1(instr_addr_o_18__BAR), .A2(n10298), .ZN(n3013) );
  NAND2_X1 U626 ( .A1(n4111), .A2(n4126), .ZN(n4129) );
  AND2_X1 U627 ( .A1(n3000), .A2(n9939), .ZN(n4519) );
  BUF_X2 U628 ( .A(n500), .Z(n3000) );
  NOR2_X1 U629 ( .A1(n4786), .A2(n235), .ZN(n4798) );
  OR2_X1 U630 ( .A1(instr_addr_o_18__BAR), .A2(n7571), .ZN(n4253) );
  INV_X2 U631 ( .A(n699), .ZN(n4644) );
  NAND2_X1 U632 ( .A1(n12156), .A2(n236), .ZN(n5001) );
  OR2_X1 U633 ( .A1(n4452), .A2(n4451), .ZN(n242) );
  NAND2_X1 U634 ( .A1(n2713), .A2(n2712), .ZN(n238) );
  AOI21_X1 U635 ( .B1(n5946), .B2(n12009), .A(n239), .ZN(n5954) );
  NAND2_X1 U636 ( .A1(n3239), .A2(n3238), .ZN(n240) );
  NAND2_X1 U637 ( .A1(n3225), .A2(n7927), .ZN(n3237) );
  NAND3_X1 U638 ( .A1(n2333), .A2(n244), .A3(n243), .ZN(n2348) );
  INV_X1 U639 ( .A(n2307), .ZN(n243) );
  NAND3_X1 U642 ( .A1(n2348), .A2(n2346), .A3(n2347), .ZN(n245) );
  NAND2_X1 U643 ( .A1(n1302), .A2(n1303), .ZN(n1304) );
  INV_X2 U645 ( .A(n2424), .ZN(n4605) );
  INV_X1 U646 ( .A(n5302), .ZN(n5847) );
  AOI21_X1 U647 ( .B1(n5024), .B2(n5030), .A(n246), .ZN(n5035) );
  NAND2_X1 U648 ( .A1(n12152), .A2(n648), .ZN(n5030) );
  NAND2_X1 U649 ( .A1(n247), .A2(n2515), .ZN(n2561) );
  BUF_X2 U650 ( .A(n2739), .Z(instr_addr_o_14__BAR) );
  NAND3_X1 U651 ( .A1(n5142), .A2(n5140), .A3(n5141), .ZN(n5324) );
  NAND2_X1 U652 ( .A1(n248), .A2(n167), .ZN(n1642) );
  OAI21_X1 U653 ( .B1(n3098), .B2(n3097), .A(n3096), .ZN(n249) );
  NAND2_X1 U654 ( .A1(n5723), .A2(n5722), .ZN(n257) );
  NAND3_X1 U655 ( .A1(n166), .A2(n256), .A3(n5724), .ZN(n5725) );
  NAND3_X1 U656 ( .A1(n3753), .A2(n250), .A3(n3752), .ZN(n3754) );
  NOR2_X1 U657 ( .A1(n3751), .A2(n3750), .ZN(n250) );
  AND2_X1 U658 ( .A1(n5031), .A2(n6833), .ZN(n2249) );
  NAND4_X1 U659 ( .A1(n5324), .A2(n251), .A3(n5322), .A4(n5323), .ZN(n6045) );
  NAND4_X1 U660 ( .A1(n5311), .A2(n5308), .A3(n5310), .A4(n5309), .ZN(n251) );
  NAND2_X1 U661 ( .A1(n5300), .A2(n5301), .ZN(n5307) );
  NOR2_X1 U663 ( .A1(n5717), .A2(n257), .ZN(n256) );
  AOI21_X1 U664 ( .B1(n1329), .B2(n322), .A(n258), .ZN(n1363) );
  NAND3_X1 U665 ( .A1(n1469), .A2(n1439), .A3(n259), .ZN(n1465) );
  NAND3_X1 U666 ( .A1(n1775), .A2(n5803), .A3(n5808), .ZN(n1736) );
  NAND2_X1 U667 ( .A1(n261), .A2(n260), .ZN(n310) );
  NAND2_X1 U668 ( .A1(n154), .A2(n1322), .ZN(n260) );
  NAND2_X1 U669 ( .A1(n213), .A2(n5261), .ZN(n261) );
  AOI22_X1 U670 ( .A1(n5730), .A2(n5729), .B1(n5728), .B2(n262), .ZN(n6043) );
  OAI21_X1 U671 ( .B1(n5726), .B2(n5727), .A(n5725), .ZN(n262) );
  NAND2_X1 U672 ( .A1(n12203), .A2(n11194), .ZN(n5715) );
  INV_X1 U673 ( .A(n3188), .ZN(n3165) );
  NAND2_X1 U674 ( .A1(n3193), .A2(n263), .ZN(n3188) );
  INV_X2 U675 ( .A(n2739), .ZN(n4788) );
  NAND2_X1 U676 ( .A1(n265), .A2(n264), .ZN(n5142) );
  NAND2_X1 U678 ( .A1(n3189), .A2(n266), .ZN(n3163) );
  NAND2_X1 U679 ( .A1(n5979), .A2(n3146), .ZN(n3189) );
  INV_X2 U680 ( .A(n537), .ZN(instr_addr_o_11_) );
  INV_X2 U681 ( .A(n3192), .ZN(n5550) );
  INV_X2 U682 ( .A(n3846), .ZN(n5040) );
  OR2_X1 U683 ( .A1(n4687), .A2(n4688), .ZN(n267) );
  OR2_X1 U685 ( .A1(n3000), .A2(pmp_addr_i[432]), .ZN(n4590) );
  INV_X2 U686 ( .A(n1658), .ZN(n4859) );
  INV_X2 U687 ( .A(n3192), .ZN(n4900) );
  OAI211_X1 U688 ( .C1(n2972), .C2(n2971), .A(n269), .B(n268), .ZN(n3023) );
  NAND2_X1 U689 ( .A1(n2969), .A2(n2970), .ZN(n268) );
  NAND2_X1 U690 ( .A1(n5366), .A2(n5367), .ZN(n271) );
  OR2_X1 U692 ( .A1(n4234), .A2(n9842), .ZN(n4518) );
  OAI211_X1 U694 ( .C1(n2639), .C2(n2638), .A(n275), .B(n274), .ZN(n2663) );
  NAND3_X1 U695 ( .A1(n6038), .A2(n6036), .A3(n6037), .ZN(n6039) );
  NAND2_X1 U697 ( .A1(n4441), .A2(n278), .ZN(n4437) );
  OAI21_X1 U698 ( .B1(n285), .B2(n282), .A(n279), .ZN(n5254) );
  NOR2_X1 U699 ( .A1(n5252), .A2(n5891), .ZN(n281) );
  AOI21_X1 U700 ( .B1(n284), .B2(n5302), .A(n283), .ZN(n282) );
  INV_X1 U701 ( .A(n289), .ZN(n284) );
  NAND2_X1 U703 ( .A1(n5295), .A2(n286), .ZN(n295) );
  NAND4_X1 U704 ( .A1(n5895), .A2(n5893), .A3(n5894), .A4(n289), .ZN(n5896) );
  NAND2_X1 U705 ( .A1(instr_addr_o_11_), .A2(n10946), .ZN(n289) );
  NAND2_X1 U706 ( .A1(instr_addr_o_11_), .A2(n288), .ZN(n287) );
  NAND2_X1 U707 ( .A1(n4621), .A2(n4646), .ZN(n4648) );
  NAND2_X1 U708 ( .A1(n4653), .A2(n292), .ZN(n4640) );
  NAND4_X1 U709 ( .A1(n4621), .A2(n4653), .A3(n4646), .A4(n292), .ZN(n290) );
  NAND2_X1 U710 ( .A1(instr_addr_o_28_), .A2(n2511), .ZN(n4653) );
  INV_X1 U711 ( .A(n5295), .ZN(n294) );
  NAND2_X1 U712 ( .A1(n295), .A2(n5895), .ZN(n5273) );
  OAI211_X1 U713 ( .C1(n2894), .C2(n2893), .A(n297), .B(n296), .ZN(n2917) );
  NAND2_X1 U714 ( .A1(n12266), .A2(n2891), .ZN(n2912) );
  INV_X2 U715 ( .A(instr_addr_i[14]), .ZN(n2739) );
  NAND2_X1 U716 ( .A1(n300), .A2(n298), .ZN(n4418) );
  NAND2_X1 U717 ( .A1(n300), .A2(n299), .ZN(n4440) );
  NAND2_X1 U718 ( .A1(n5979), .A2(n1155), .ZN(n300) );
  NAND2_X1 U719 ( .A1(n301), .A2(n336), .ZN(n7319) );
  NAND3_X1 U720 ( .A1(n302), .A2(n7245), .A3(n7246), .ZN(n301) );
  OAI211_X1 U721 ( .C1(n7125), .C2(n7124), .A(n304), .B(n303), .ZN(n302) );
  INV_X1 U722 ( .A(n7121), .ZN(n303) );
  NAND2_X1 U723 ( .A1(n7123), .A2(n7122), .ZN(n304) );
  NAND4_X1 U724 ( .A1(n308), .A2(n2756), .A3(n331), .A4(n2757), .ZN(n305) );
  NAND2_X1 U725 ( .A1(n307), .A2(n331), .ZN(n306) );
  NAND2_X1 U726 ( .A1(n310), .A2(n173), .ZN(n309) );
  NOR2_X1 U727 ( .A1(n1335), .A2(n1326), .ZN(n311) );
  NAND3_X1 U728 ( .A1(n1391), .A2(n1398), .A3(n313), .ZN(n312) );
  NAND2_X1 U729 ( .A1(n138), .A2(n1350), .ZN(n1391) );
  INV_X2 U730 ( .A(n2896), .ZN(n3100) );
  NAND2_X1 U731 ( .A1(n314), .A2(n3323), .ZN(n3324) );
  INV_X1 U732 ( .A(n4504), .ZN(n3503) );
  AND2_X1 U733 ( .A1(n9329), .A2(pmp_cfg_i[82]), .ZN(n315) );
  OR2_X1 U734 ( .A1(n5814), .A2(n1744), .ZN(n316) );
  OR2_X1 U735 ( .A1(n8063), .A2(n8066), .ZN(n317) );
  NOR2_X1 U736 ( .A1(n1186), .A2(n1275), .ZN(n1266) );
  AND2_X1 U737 ( .A1(n4660), .A2(n8062), .ZN(n318) );
  AND3_X1 U738 ( .A1(n685), .A2(n4861), .A3(n4869), .ZN(n319) );
  OR2_X1 U739 ( .A1(instr_addr_o_9_), .A2(n4848), .ZN(n320) );
  AND2_X1 U740 ( .A1(n2742), .A2(n2744), .ZN(n321) );
  AND4_X1 U741 ( .A1(n1321), .A2(n173), .A3(n1320), .A4(n1319), .ZN(n322) );
  AND2_X1 U742 ( .A1(n3883), .A2(n3882), .ZN(n323) );
  OR2_X1 U743 ( .A1(n3675), .A2(n3654), .ZN(n324) );
  NOR2_X1 U744 ( .A1(n2732), .A2(n2731), .ZN(n326) );
  NOR2_X1 U745 ( .A1(n2679), .A2(n2678), .ZN(n327) );
  OR2_X1 U746 ( .A1(n3683), .A2(n3687), .ZN(n328) );
  OR2_X1 U747 ( .A1(n3683), .A2(n3651), .ZN(n329) );
  OR2_X1 U748 ( .A1(n3661), .A2(n3652), .ZN(n330) );
  OR2_X1 U749 ( .A1(n2838), .A2(n2837), .ZN(n331) );
  AND3_X1 U750 ( .A1(n2561), .A2(n2560), .A3(n2559), .ZN(n332) );
  AND3_X1 U751 ( .A1(n1005), .A2(n986), .A3(n1015), .ZN(n333) );
  XOR2_X1 U752 ( .A(n6019), .B(n9199), .Z(n334) );
  OR2_X1 U753 ( .A1(n11082), .A2(n7316), .ZN(n336) );
  AND2_X1 U754 ( .A1(n4234), .A2(n7322), .ZN(n337) );
  AND2_X1 U755 ( .A1(n1641), .A2(n1640), .ZN(n338) );
  AND3_X1 U756 ( .A1(n1617), .A2(n1616), .A3(n1615), .ZN(n339) );
  NOR2_X1 U757 ( .A1(n10211), .A2(n10123), .ZN(n10214) );
  NOR2_X1 U758 ( .A1(n11769), .A2(n11761), .ZN(n4671) );
  AND2_X1 U759 ( .A1(n2398), .A2(n3278), .ZN(n2428) );
  INV_X1 U760 ( .A(n11068), .ZN(n5356) );
  NOR2_X1 U761 ( .A1(n318), .A2(n317), .ZN(n3801) );
  INV_X1 U762 ( .A(n4506), .ZN(n3502) );
  AND2_X1 U763 ( .A1(n2462), .A2(n3300), .ZN(n2471) );
  AND3_X1 U764 ( .A1(n3312), .A2(n3311), .A3(n3310), .ZN(n3328) );
  OR2_X1 U765 ( .A1(n5262), .A2(n7659), .ZN(n3278) );
  OR2_X1 U766 ( .A1(n1668), .A2(n1674), .ZN(n1715) );
  AND2_X1 U767 ( .A1(n2472), .A2(n2471), .ZN(n2476) );
  OR2_X1 U769 ( .A1(n1171), .A2(n1248), .ZN(n1243) );
  AND2_X1 U770 ( .A1(n676), .A2(n645), .ZN(n646) );
  NOR2_X1 U771 ( .A1(n11487), .A2(n2693), .ZN(n11476) );
  INV_X1 U772 ( .A(n4637), .ZN(n4627) );
  NOR3_X1 U773 ( .A1(n4146), .A2(n4120), .A3(n4119), .ZN(n4145) );
  INV_X1 U774 ( .A(n3172), .ZN(n3157) );
  OR2_X1 U775 ( .A1(n1346), .A2(n1345), .ZN(n1347) );
  AND2_X1 U776 ( .A1(n851), .A2(n837), .ZN(n838) );
  NOR2_X1 U777 ( .A1(n485), .A2(n489), .ZN(n486) );
  NOR2_X1 U778 ( .A1(n2273), .A2(n2272), .ZN(n2274) );
  AND3_X1 U779 ( .A1(n5305), .A2(n5304), .A3(n5833), .ZN(n5306) );
  AND2_X1 U780 ( .A1(n5098), .A2(n5139), .ZN(n5124) );
  AND3_X1 U781 ( .A1(n9338), .A2(n9337), .A3(n9336), .ZN(n9339) );
  OR2_X1 U782 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U783 ( .A1(n4890), .A2(n4889), .ZN(n4917) );
  INV_X1 U784 ( .A(n4326), .ZN(n4359) );
  NOR3_X1 U786 ( .A1(n2345), .A2(n2349), .A3(n2370), .ZN(n2346) );
  OR2_X1 U787 ( .A1(n2558), .A2(n2557), .ZN(n2559) );
  INV_X1 U788 ( .A(instr_addr_i[10]), .ZN(n545) );
  INV_X2 U789 ( .A(n212), .ZN(n5270) );
  INV_X1 U790 ( .A(instr_addr_i[8]), .ZN(n2707) );
  INV_X1 U791 ( .A(n2707), .ZN(n2623) );
  INV_X1 U792 ( .A(instr_addr_i[16]), .ZN(n433) );
  INV_X2 U794 ( .A(n3228), .ZN(n5229) );
  INV_X1 U796 ( .A(instr_addr_i[21]), .ZN(n3984) );
  INV_X1 U797 ( .A(n3984), .ZN(n5191) );
  INV_X2 U799 ( .A(instr_addr_o_4__BAR), .ZN(n12150) );
  INV_X1 U800 ( .A(instr_addr_i[22]), .ZN(n3288) );
  INV_X2 U801 ( .A(n3288), .ZN(n12157) );
  INV_X1 U802 ( .A(instr_addr_i[27]), .ZN(n580) );
  INV_X1 U804 ( .A(instr_addr_i[15]), .ZN(n3531) );
  INV_X2 U805 ( .A(n3531), .ZN(instr_addr_o_15_) );
  INV_X1 U806 ( .A(instr_addr_i[9]), .ZN(n543) );
  INV_X1 U807 ( .A(instr_addr_i[26]), .ZN(n1131) );
  INV_X2 U808 ( .A(n1131), .ZN(n12158) );
  INV_X1 U809 ( .A(instr_addr_i[30]), .ZN(n376) );
  INV_X1 U810 ( .A(instr_addr_i[28]), .ZN(n372) );
  INV_X2 U811 ( .A(n3045), .ZN(instr_addr_o_28_) );
  INV_X1 U812 ( .A(instr_addr_i[29]), .ZN(n3041) );
  INV_X1 U813 ( .A(instr_addr_i[11]), .ZN(n537) );
  INV_X1 U814 ( .A(instr_addr_i[17]), .ZN(n687) );
  INV_X1 U815 ( .A(instr_addr_i[6]), .ZN(n466) );
  INV_X1 U817 ( .A(instr_addr_i[24]), .ZN(n3275) );
  INV_X1 U818 ( .A(instr_addr_i[7]), .ZN(n811) );
  INV_X1 U819 ( .A(instr_addr_i[12]), .ZN(n679) );
  INV_X1 U820 ( .A(instr_addr_i[23]), .ZN(n1658) );
  BUF_X1 U821 ( .A(instr_addr_i[23]), .Z(instr_addr_o_23_) );
  INV_X1 U822 ( .A(instr_addr_i[19]), .ZN(n2339) );
  INV_X1 U823 ( .A(n2339), .ZN(n362) );
  INV_X1 U824 ( .A(instr_addr_i[5]), .ZN(n467) );
  INV_X1 U825 ( .A(n467), .ZN(instr_addr_o_5_) );
  BUF_X1 U826 ( .A(instr_addr_i[13]), .Z(n937) );
  INV_X1 U827 ( .A(instr_addr_i[18]), .ZN(n500) );
  INV_X1 U828 ( .A(n3000), .ZN(gte_x_382_A_16_) );
  INV_X1 U829 ( .A(pmp_cfg_i[59]), .ZN(n471) );
  INV_X1 U830 ( .A(pmp_addr_i[220]), .ZN(n723) );
  AND3_X1 U831 ( .A1(pmp_addr_i[228]), .A2(pmp_addr_i[227]), .A3(
        pmp_addr_i[226]), .ZN(n450) );
  AND2_X1 U832 ( .A1(pmp_addr_i[224]), .A2(pmp_addr_i[225]), .ZN(n11037) );
  NAND4_X1 U833 ( .A1(n450), .A2(n11037), .A3(pmp_addr_i[229]), .A4(
        pmp_addr_i[230]), .ZN(n11062) );
  INV_X1 U834 ( .A(pmp_addr_i[231]), .ZN(n1741) );
  NAND3_X1 U835 ( .A1(pmp_addr_i[233]), .A2(pmp_addr_i[236]), .A3(
        pmp_addr_i[232]), .ZN(n341) );
  NAND2_X1 U836 ( .A1(pmp_addr_i[235]), .A2(pmp_addr_i[234]), .ZN(n340) );
  NOR2_X1 U837 ( .A1(n341), .A2(n340), .ZN(n413) );
  NAND2_X1 U838 ( .A1(n11068), .A2(n413), .ZN(n5405) );
  OR2_X1 U839 ( .A1(n5405), .A2(n497), .ZN(n5384) );
  INV_X1 U840 ( .A(pmp_addr_i[238]), .ZN(n1727) );
  OAI21_X1 U841 ( .B1(n11050), .B2(n501), .A(pmp_cfg_i[60]), .ZN(n5326) );
  NAND2_X1 U842 ( .A1(n5326), .A2(pmp_cfg_i[59]), .ZN(n5337) );
  NAND2_X1 U843 ( .A1(n5337), .A2(pmp_addr_i[252]), .ZN(n342) );
  OAI21_X1 U844 ( .B1(n432), .B2(n723), .A(n342), .ZN(n7247) );
  INV_X1 U845 ( .A(n7247), .ZN(n343) );
  NOR2_X1 U846 ( .A1(n4753), .A2(n343), .ZN(n378) );
  INV_X2 U847 ( .A(n3041), .ZN(instr_addr_o_29_) );
  INV_X1 U848 ( .A(pmp_addr_i[219]), .ZN(n726) );
  NAND2_X1 U849 ( .A1(n5337), .A2(pmp_addr_i[251]), .ZN(n344) );
  OAI21_X1 U850 ( .B1(n432), .B2(n726), .A(n344), .ZN(n7290) );
  INV_X1 U851 ( .A(n7290), .ZN(n375) );
  NOR2_X1 U852 ( .A1(n5149), .A2(n375), .ZN(n345) );
  NOR2_X1 U853 ( .A1(n378), .A2(n345), .ZN(n381) );
  INV_X1 U854 ( .A(pmp_addr_i[221]), .ZN(n728) );
  NAND2_X1 U855 ( .A1(n5337), .A2(pmp_addr_i[253]), .ZN(n12089) );
  OAI21_X1 U856 ( .B1(n432), .B2(n728), .A(n12089), .ZN(n7309) );
  NOR2_X1 U857 ( .A1(pmp_addr_i[222]), .A2(pmp_addr_i[223]), .ZN(n10453) );
  INV_X1 U858 ( .A(n10453), .ZN(n397) );
  AOI21_X1 U859 ( .B1(n4005), .B2(n7309), .A(n397), .ZN(n382) );
  INV_X2 U860 ( .A(n372), .ZN(n5368) );
  INV_X1 U861 ( .A(pmp_addr_i[218]), .ZN(n730) );
  NAND2_X1 U862 ( .A1(n5337), .A2(pmp_addr_i[250]), .ZN(n346) );
  OAI21_X1 U863 ( .B1(n432), .B2(n730), .A(n346), .ZN(n7295) );
  INV_X1 U864 ( .A(n7295), .ZN(n347) );
  OR2_X1 U865 ( .A1(n5368), .A2(n347), .ZN(n370) );
  INV_X1 U866 ( .A(instr_addr_i[27]), .ZN(n4000) );
  BUF_X1 U867 ( .A(n4000), .Z(n4652) );
  INV_X1 U868 ( .A(pmp_addr_i[217]), .ZN(n733) );
  NAND2_X1 U869 ( .A1(n5337), .A2(pmp_addr_i[249]), .ZN(n348) );
  OAI21_X1 U870 ( .B1(n432), .B2(n733), .A(n348), .ZN(n7255) );
  NAND2_X1 U871 ( .A1(n4652), .A2(n7255), .ZN(n349) );
  NAND4_X1 U872 ( .A1(n381), .A2(n382), .A3(n370), .A4(n349), .ZN(n411) );
  INV_X1 U873 ( .A(pmp_addr_i[213]), .ZN(n704) );
  NAND2_X1 U874 ( .A1(n5337), .A2(pmp_addr_i[245]), .ZN(n350) );
  OAI21_X1 U875 ( .B1(n432), .B2(n704), .A(n350), .ZN(n7249) );
  INV_X1 U876 ( .A(instr_addr_i[25]), .ZN(n699) );
  INV_X1 U877 ( .A(pmp_addr_i[215]), .ZN(n701) );
  NAND2_X1 U878 ( .A1(n5337), .A2(pmp_addr_i[247]), .ZN(n351) );
  OAI21_X1 U879 ( .B1(n432), .B2(n701), .A(n351), .ZN(n7257) );
  INV_X1 U880 ( .A(n7257), .ZN(n391) );
  NOR2_X1 U881 ( .A1(n4644), .A2(n391), .ZN(n354) );
  INV_X1 U882 ( .A(pmp_addr_i[216]), .ZN(n697) );
  NAND2_X1 U883 ( .A1(n5337), .A2(pmp_addr_i[248]), .ZN(n352) );
  OAI21_X1 U884 ( .B1(n432), .B2(n697), .A(n352), .ZN(n7258) );
  INV_X1 U885 ( .A(n7258), .ZN(n353) );
  NOR2_X1 U886 ( .A1(instr_addr_o_26_), .A2(n353), .ZN(n393) );
  NOR2_X1 U887 ( .A1(n354), .A2(n393), .ZN(n396) );
  INV_X2 U888 ( .A(n3275), .ZN(n5330) );
  INV_X1 U889 ( .A(pmp_addr_i[214]), .ZN(n706) );
  NAND2_X1 U890 ( .A1(n5337), .A2(pmp_addr_i[246]), .ZN(n355) );
  OAI21_X1 U891 ( .B1(n432), .B2(n706), .A(n355), .ZN(n7250) );
  INV_X1 U892 ( .A(n7250), .ZN(n356) );
  OR2_X1 U893 ( .A1(n5330), .A2(n356), .ZN(n387) );
  OAI211_X1 U894 ( .C1(n5208), .C2(n7211), .A(n387), .B(n396), .ZN(n403) );
  OR2_X1 U895 ( .A1(n411), .A2(n403), .ZN(n386) );
  INV_X1 U896 ( .A(pmp_addr_i[212]), .ZN(n712) );
  NAND2_X1 U897 ( .A1(n5337), .A2(pmp_addr_i[244]), .ZN(n357) );
  OAI21_X1 U898 ( .B1(n432), .B2(n712), .A(n357), .ZN(n7289) );
  INV_X1 U899 ( .A(n7289), .ZN(n358) );
  NOR2_X1 U900 ( .A1(n5181), .A2(n358), .ZN(n367) );
  INV_X1 U901 ( .A(instr_addr_i[21]), .ZN(n3819) );
  INV_X1 U902 ( .A(pmp_addr_i[211]), .ZN(n710) );
  NAND2_X1 U903 ( .A1(n5337), .A2(pmp_addr_i[243]), .ZN(n359) );
  OAI21_X1 U904 ( .B1(n432), .B2(n710), .A(n359), .ZN(n7296) );
  INV_X1 U905 ( .A(n7296), .ZN(n365) );
  NOR2_X1 U906 ( .A1(n367), .A2(n360), .ZN(n404) );
  INV_X2 U907 ( .A(n3290), .ZN(n5187) );
  INV_X1 U908 ( .A(pmp_addr_i[210]), .ZN(n717) );
  NAND2_X1 U909 ( .A1(n5337), .A2(pmp_addr_i[242]), .ZN(n361) );
  OAI21_X1 U910 ( .B1(n432), .B2(n717), .A(n361), .ZN(n7256) );
  INV_X1 U911 ( .A(n7256), .ZN(n5347) );
  NOR2_X1 U912 ( .A1(n5187), .A2(n5347), .ZN(n405) );
  INV_X1 U913 ( .A(pmp_addr_i[209]), .ZN(n715) );
  NAND2_X1 U914 ( .A1(n5337), .A2(pmp_addr_i[241]), .ZN(n363) );
  OAI21_X1 U915 ( .B1(n432), .B2(n715), .A(n363), .ZN(n7248) );
  NAND2_X1 U916 ( .A1(n3793), .A2(n7201), .ZN(n364) );
  INV_X1 U917 ( .A(instr_addr_i[20]), .ZN(n1996) );
  BUF_X1 U918 ( .A(n1996), .Z(n2569) );
  OAI22_X1 U919 ( .A1(n405), .A2(n364), .B1(n2569), .B2(n7256), .ZN(n369) );
  INV_X2 U920 ( .A(n3984), .ZN(n3152) );
  NAND2_X1 U921 ( .A1(n3152), .A2(n365), .ZN(n366) );
  INV_X1 U922 ( .A(instr_addr_i[22]), .ZN(n2103) );
  OAI22_X1 U923 ( .A1(n367), .A2(n366), .B1(n5192), .B2(n7289), .ZN(n368) );
  AOI21_X1 U924 ( .B1(n404), .B2(n369), .A(n368), .ZN(n385) );
  INV_X1 U925 ( .A(n370), .ZN(n374) );
  INV_X1 U926 ( .A(n7255), .ZN(n371) );
  NAND2_X1 U927 ( .A1(instr_addr_o_27_), .A2(n371), .ZN(n373) );
  OAI22_X1 U929 ( .A1(n374), .A2(n373), .B1(n5111), .B2(n7295), .ZN(n380) );
  NAND2_X1 U930 ( .A1(n4900), .A2(n375), .ZN(n377) );
  OAI22_X1 U931 ( .A1(n378), .A2(n377), .B1(n4658), .B2(n7247), .ZN(n379) );
  AOI21_X1 U932 ( .B1(n381), .B2(n380), .A(n379), .ZN(n384) );
  INV_X1 U933 ( .A(n382), .ZN(n383) );
  OAI22_X1 U934 ( .A1(n386), .A2(n385), .B1(n384), .B2(n383), .ZN(n402) );
  INV_X1 U935 ( .A(n387), .ZN(n389) );
  NAND2_X1 U936 ( .A1(n5208), .A2(n7211), .ZN(n388) );
  INV_X1 U937 ( .A(instr_addr_i[24]), .ZN(n4135) );
  BUF_X1 U938 ( .A(n4135), .Z(n1269) );
  OAI22_X1 U939 ( .A1(n389), .A2(n388), .B1(n2580), .B2(n7250), .ZN(n395) );
  INV_X2 U940 ( .A(n699), .ZN(n5202) );
  NAND2_X1 U941 ( .A1(n5202), .A2(n391), .ZN(n392) );
  INV_X1 U942 ( .A(instr_addr_i[26]), .ZN(n1026) );
  BUF_X1 U943 ( .A(n1026), .Z(n1273) );
  OAI22_X1 U944 ( .A1(n393), .A2(n392), .B1(n1273), .B2(n7258), .ZN(n394) );
  AOI21_X1 U945 ( .B1(n12215), .B2(n395), .A(n394), .ZN(n400) );
  INV_X1 U946 ( .A(n7309), .ZN(n398) );
  NAND3_X1 U947 ( .A1(instr_addr_o_31_), .A2(n398), .A3(n10453), .ZN(n399) );
  OAI21_X1 U948 ( .B1(n400), .B2(n411), .A(n399), .ZN(n401) );
  NOR2_X1 U949 ( .A1(n402), .A2(n401), .ZN(n496) );
  INV_X1 U950 ( .A(n403), .ZN(n410) );
  INV_X1 U951 ( .A(n404), .ZN(n408) );
  INV_X1 U952 ( .A(n405), .ZN(n406) );
  OAI21_X1 U953 ( .B1(instr_addr_o_19_), .B2(n7201), .A(n406), .ZN(n407) );
  NOR2_X1 U954 ( .A1(n408), .A2(n407), .ZN(n409) );
  NOR2_X1 U955 ( .A1(n412), .A2(n411), .ZN(n493) );
  INV_X1 U956 ( .A(pmp_addr_i[204]), .ZN(n415) );
  NOR2_X1 U957 ( .A1(n5356), .A2(n471), .ZN(n481) );
  INV_X1 U958 ( .A(pmp_cfg_i[60]), .ZN(n454) );
  AOI21_X1 U959 ( .B1(n481), .B2(n413), .A(n454), .ZN(n436) );
  NAND2_X1 U960 ( .A1(n436), .A2(pmp_addr_i[236]), .ZN(n414) );
  OAI21_X1 U961 ( .B1(n432), .B2(n415), .A(n414), .ZN(n7302) );
  INV_X1 U962 ( .A(n7302), .ZN(n7281) );
  NOR2_X1 U963 ( .A1(instr_addr_o_14_), .A2(n7281), .ZN(n426) );
  NAND2_X1 U964 ( .A1(n481), .A2(pmp_addr_i[232]), .ZN(n421) );
  NAND2_X1 U965 ( .A1(pmp_addr_i[234]), .A2(pmp_addr_i[233]), .ZN(n416) );
  OAI21_X1 U966 ( .B1(n421), .B2(n416), .A(pmp_cfg_i[60]), .ZN(n420) );
  INV_X1 U967 ( .A(pmp_addr_i[235]), .ZN(n5390) );
  INV_X1 U968 ( .A(n432), .ZN(n7246) );
  NAND2_X1 U969 ( .A1(n7246), .A2(pmp_addr_i[203]), .ZN(n417) );
  OAI21_X1 U970 ( .B1(n420), .B2(n5390), .A(n417), .ZN(n7133) );
  INV_X1 U971 ( .A(n7133), .ZN(n425) );
  NOR2_X1 U972 ( .A1(n5997), .A2(n425), .ZN(n418) );
  INV_X1 U973 ( .A(pmp_addr_i[234]), .ZN(n5389) );
  NAND2_X1 U974 ( .A1(n7246), .A2(pmp_addr_i[202]), .ZN(n419) );
  OAI21_X1 U975 ( .B1(n420), .B2(n5389), .A(n419), .ZN(n7131) );
  INV_X1 U976 ( .A(n7131), .ZN(n7273) );
  OR2_X1 U977 ( .A1(n5245), .A2(n7273), .ZN(n447) );
  INV_X1 U978 ( .A(n447), .ZN(n424) );
  INV_X1 U979 ( .A(pmp_addr_i[201]), .ZN(n423) );
  NAND3_X1 U980 ( .A1(n421), .A2(pmp_cfg_i[60]), .A3(pmp_addr_i[233]), .ZN(
        n422) );
  OAI21_X1 U981 ( .B1(n432), .B2(n423), .A(n422), .ZN(n7130) );
  INV_X1 U982 ( .A(n7130), .ZN(n7266) );
  NAND2_X1 U983 ( .A1(instr_addr_o_11_), .A2(n7266), .ZN(n5374) );
  INV_X2 U984 ( .A(n679), .ZN(n5250) );
  NAND2_X1 U985 ( .A1(n5250), .A2(n7273), .ZN(n5355) );
  OAI21_X1 U986 ( .B1(n424), .B2(n5374), .A(n5355), .ZN(n428) );
  NAND2_X1 U987 ( .A1(n150), .A2(n425), .ZN(n5403) );
  INV_X2 U988 ( .A(n2739), .ZN(n5251) );
  NAND2_X1 U989 ( .A1(instr_addr_o_14_), .A2(n7281), .ZN(n5392) );
  OAI21_X1 U990 ( .B1(n426), .B2(n5403), .A(n5392), .ZN(n427) );
  AOI21_X1 U991 ( .B1(n448), .B2(n428), .A(n427), .ZN(n445) );
  INV_X1 U993 ( .A(pmp_addr_i[208]), .ZN(n627) );
  NAND2_X1 U994 ( .A1(n5337), .A2(pmp_addr_i[240]), .ZN(n429) );
  OAI21_X1 U995 ( .B1(n432), .B2(n627), .A(n429), .ZN(n7279) );
  INV_X1 U996 ( .A(n7279), .ZN(n430) );
  NOR2_X1 U997 ( .A1(n6019), .A2(n430), .ZN(n440) );
  INV_X1 U999 ( .A(pmp_addr_i[207]), .ZN(n630) );
  NAND2_X1 U1000 ( .A1(n5337), .A2(pmp_addr_i[239]), .ZN(n431) );
  OAI21_X1 U1001 ( .B1(n432), .B2(n630), .A(n431), .ZN(n7175) );
  INV_X1 U1002 ( .A(n7175), .ZN(n439) );
  NOR2_X1 U1003 ( .A1(n4069), .A2(n439), .ZN(n5385) );
  NOR2_X1 U1004 ( .A1(n440), .A2(n5385), .ZN(n443) );
  INV_X2 U1006 ( .A(n2896), .ZN(n5226) );
  INV_X1 U1007 ( .A(pmp_addr_i[206]), .ZN(n635) );
  NOR2_X1 U1008 ( .A1(n454), .A2(pmp_addr_i[237]), .ZN(n434) );
  OAI21_X1 U1009 ( .B1(n436), .B2(n434), .A(pmp_addr_i[238]), .ZN(n435) );
  OAI21_X1 U1010 ( .B1(n635), .B2(n432), .A(n435), .ZN(n11054) );
  INV_X1 U1011 ( .A(n11054), .ZN(n7301) );
  INV_X1 U1013 ( .A(pmp_addr_i[205]), .ZN(n633) );
  NAND2_X1 U1014 ( .A1(n436), .A2(pmp_addr_i[237]), .ZN(n437) );
  OAI21_X1 U1015 ( .B1(n432), .B2(n633), .A(n437), .ZN(n7126) );
  INV_X1 U1016 ( .A(n7126), .ZN(n7280) );
  OR2_X1 U1017 ( .A1(n12179), .A2(n7280), .ZN(n5396) );
  NAND3_X1 U1018 ( .A1(n443), .A2(n5387), .A3(n5396), .ZN(n449) );
  INV_X1 U1019 ( .A(n5387), .ZN(n438) );
  NAND2_X1 U1020 ( .A1(n208), .A2(n7280), .ZN(n5406) );
  NAND2_X1 U1021 ( .A1(n12203), .A2(n7301), .ZN(n5388) );
  OAI21_X1 U1022 ( .B1(n438), .B2(n5406), .A(n5388), .ZN(n442) );
  NAND2_X1 U1023 ( .A1(n12156), .A2(n439), .ZN(n5346) );
  OAI22_X1 U1024 ( .A1(n440), .A2(n5346), .B1(n2750), .B2(n7279), .ZN(n441) );
  AOI21_X1 U1025 ( .B1(n443), .B2(n442), .A(n441), .ZN(n444) );
  OAI21_X1 U1026 ( .B1(n445), .B2(n449), .A(n444), .ZN(n446) );
  INV_X1 U1027 ( .A(n537), .ZN(n6002) );
  NOR2_X1 U1028 ( .A1(n5364), .A2(n449), .ZN(n492) );
  AND2_X1 U1029 ( .A1(pmp_cfg_i[59]), .A2(pmp_addr_i[224]), .ZN(n459) );
  NAND3_X1 U1030 ( .A1(n450), .A2(n459), .A3(pmp_addr_i[225]), .ZN(n451) );
  NAND2_X1 U1031 ( .A1(n451), .A2(pmp_cfg_i[60]), .ZN(n474) );
  INV_X1 U1032 ( .A(pmp_addr_i[228]), .ZN(n453) );
  NAND2_X1 U1033 ( .A1(n7246), .A2(pmp_addr_i[196]), .ZN(n452) );
  OAI21_X1 U1034 ( .B1(n474), .B2(n453), .A(n452), .ZN(n7145) );
  INV_X1 U1035 ( .A(n7145), .ZN(n7137) );
  NOR2_X1 U1036 ( .A1(instr_addr_o_6_), .A2(n7137), .ZN(n468) );
  INV_X1 U1037 ( .A(pmp_addr_i[195]), .ZN(n611) );
  AND2_X1 U1038 ( .A1(pmp_addr_i[226]), .A2(pmp_addr_i[225]), .ZN(n455) );
  AOI21_X1 U1039 ( .B1(n459), .B2(n455), .A(n454), .ZN(n462) );
  NAND2_X1 U1040 ( .A1(n462), .A2(pmp_addr_i[227]), .ZN(n456) );
  OAI21_X1 U1041 ( .B1(n432), .B2(n611), .A(n456), .ZN(n7146) );
  INV_X1 U1042 ( .A(n7146), .ZN(n7136) );
  NOR2_X1 U1043 ( .A1(n5280), .A2(n7136), .ZN(n457) );
  OR2_X1 U1044 ( .A1(n468), .A2(n457), .ZN(n5336) );
  INV_X1 U1045 ( .A(pmp_addr_i[193]), .ZN(n653) );
  NAND2_X1 U1046 ( .A1(pmp_cfg_i[60]), .A2(pmp_addr_i[225]), .ZN(n458) );
  OAI22_X1 U1047 ( .A1(n432), .A2(n653), .B1(n459), .B2(n458), .ZN(n7267) );
  INV_X1 U1048 ( .A(pmp_addr_i[192]), .ZN(n461) );
  NAND2_X1 U1049 ( .A1(pmp_addr_i[224]), .A2(n471), .ZN(n460) );
  OAI21_X1 U1050 ( .B1(n432), .B2(n461), .A(n460), .ZN(n7304) );
  OR2_X1 U1051 ( .A1(n7267), .A2(n7304), .ZN(n464) );
  INV_X1 U1052 ( .A(pmp_addr_i[194]), .ZN(n657) );
  NAND2_X1 U1053 ( .A1(n462), .A2(pmp_addr_i[226]), .ZN(n463) );
  OAI21_X1 U1054 ( .B1(n432), .B2(n657), .A(n463), .ZN(n7142) );
  NAND2_X1 U1055 ( .A1(n464), .A2(n7142), .ZN(n465) );
  INV_X1 U1056 ( .A(n7142), .ZN(n7268) );
  INV_X1 U1057 ( .A(n464), .ZN(n5338) );
  AOI22_X1 U1058 ( .A1(n3836), .A2(n465), .B1(n7268), .B2(n5338), .ZN(n470) );
  NAND2_X1 U1060 ( .A1(instr_addr_o_6_), .A2(n7137), .ZN(n5377) );
  NAND2_X1 U1061 ( .A1(n5293), .A2(n7136), .ZN(n5327) );
  OR2_X1 U1062 ( .A1(n5327), .A2(n468), .ZN(n469) );
  OAI211_X1 U1063 ( .C1(n5336), .C2(n470), .A(n5377), .B(n469), .ZN(n476) );
  INV_X1 U1064 ( .A(instr_addr_i[8]), .ZN(n3894) );
  OAI21_X1 U1065 ( .B1(n11062), .B2(n471), .A(pmp_cfg_i[60]), .ZN(n483) );
  INV_X1 U1066 ( .A(pmp_addr_i[230]), .ZN(n1752) );
  NAND2_X1 U1067 ( .A1(n7246), .A2(pmp_addr_i[198]), .ZN(n472) );
  OAI21_X1 U1068 ( .B1(n483), .B2(n1752), .A(n472), .ZN(n7151) );
  INV_X1 U1069 ( .A(n7151), .ZN(n7274) );
  NOR2_X1 U1070 ( .A1(n5342), .A2(n7274), .ZN(n478) );
  INV_X1 U1071 ( .A(pmp_addr_i[229]), .ZN(n473) );
  INV_X1 U1072 ( .A(pmp_addr_i[197]), .ZN(n667) );
  OAI22_X1 U1073 ( .A1(n474), .A2(n473), .B1(n667), .B2(n432), .ZN(n7310) );
  INV_X1 U1074 ( .A(n7310), .ZN(n477) );
  NOR2_X1 U1075 ( .A1(n12267), .A2(n477), .ZN(n475) );
  NOR2_X1 U1076 ( .A1(n478), .A2(n475), .ZN(n5383) );
  NAND2_X1 U1077 ( .A1(n476), .A2(n5383), .ZN(n487) );
  BUF_X2 U1078 ( .A(n811), .Z(n4200) );
  INV_X2 U1079 ( .A(n4200), .ZN(n5740) );
  NAND2_X1 U1080 ( .A1(n5740), .A2(n477), .ZN(n5351) );
  INV_X2 U1081 ( .A(n3894), .ZN(n5269) );
  NAND2_X1 U1082 ( .A1(n205), .A2(n7274), .ZN(n5350) );
  OAI21_X1 U1083 ( .B1(n478), .B2(n5351), .A(n5350), .ZN(n485) );
  NAND2_X1 U1084 ( .A1(pmp_cfg_i[60]), .A2(pmp_addr_i[232]), .ZN(n480) );
  NAND2_X1 U1085 ( .A1(n7246), .A2(pmp_addr_i[200]), .ZN(n479) );
  OAI21_X1 U1086 ( .B1(n481), .B2(n480), .A(n479), .ZN(n7155) );
  INV_X1 U1087 ( .A(n7155), .ZN(n7265) );
  NOR2_X1 U1088 ( .A1(n12202), .A2(n7265), .ZN(n5329) );
  NAND2_X1 U1089 ( .A1(n7246), .A2(pmp_addr_i[199]), .ZN(n482) );
  OAI21_X1 U1090 ( .B1(n483), .B2(n1741), .A(n482), .ZN(n7154) );
  INV_X1 U1091 ( .A(n7154), .ZN(n7275) );
  NAND2_X1 U1092 ( .A1(instr_addr_o_9_), .A2(n7275), .ZN(n484) );
  NAND2_X1 U1093 ( .A1(instr_addr_o_10_), .A2(n7265), .ZN(n5328) );
  OAI21_X1 U1094 ( .B1(n5329), .B2(n484), .A(n5328), .ZN(n489) );
  NAND2_X1 U1095 ( .A1(n487), .A2(n486), .ZN(n491) );
  NOR2_X1 U1096 ( .A1(n4204), .A2(n7275), .ZN(n5398) );
  NOR2_X1 U1097 ( .A1(n5398), .A2(n5329), .ZN(n488) );
  NAND4_X1 U1098 ( .A1(n493), .A2(n492), .A3(n491), .A4(n490), .ZN(n494) );
  NAND2_X1 U1099 ( .A1(n5226), .A2(n1727), .ZN(n506) );
  INV_X1 U1100 ( .A(pmp_addr_i[237]), .ZN(n497) );
  NOR2_X1 U1101 ( .A1(n12179), .A2(n497), .ZN(n498) );
  BUF_X2 U1102 ( .A(n3228), .Z(n5058) );
  AOI22_X1 U1103 ( .A1(n506), .A2(n498), .B1(n5058), .B2(pmp_addr_i[238]), 
        .ZN(n505) );
  INV_X2 U1104 ( .A(n500), .ZN(n5047) );
  NAND2_X1 U1105 ( .A1(gte_x_382_A_16_), .A2(n1721), .ZN(n503) );
  OAI21_X1 U1106 ( .B1(n5048), .B2(pmp_addr_i[239]), .A(n503), .ZN(n508) );
  INV_X1 U1107 ( .A(pmp_addr_i[239]), .ZN(n501) );
  NOR2_X1 U1108 ( .A1(n12265), .A2(n501), .ZN(n502) );
  AOI22_X1 U1109 ( .A1(n503), .A2(n502), .B1(n2082), .B2(pmp_addr_i[240]), 
        .ZN(n504) );
  OAI21_X1 U1110 ( .B1(n505), .B2(n508), .A(n504), .ZN(n533) );
  OAI21_X1 U1112 ( .B1(n4578), .B2(pmp_addr_i[237]), .A(n506), .ZN(n507) );
  NOR2_X1 U1113 ( .A1(n508), .A2(n507), .ZN(n536) );
  OR2_X1 U1114 ( .A1(n533), .A2(n536), .ZN(n535) );
  INV_X1 U1115 ( .A(instr_addr_i[29]), .ZN(n3192) );
  BUF_X1 U1116 ( .A(n3192), .Z(n4656) );
  INV_X1 U1117 ( .A(pmp_addr_i[252]), .ZN(n509) );
  NAND2_X1 U1118 ( .A1(n12161), .A2(n509), .ZN(n586) );
  OAI21_X1 U1119 ( .B1(n4656), .B2(pmp_addr_i[251]), .A(n586), .ZN(n588) );
  BUF_X2 U1120 ( .A(n580), .Z(n5094) );
  INV_X1 U1121 ( .A(pmp_addr_i[250]), .ZN(n510) );
  NAND2_X1 U1122 ( .A1(n5368), .A2(n510), .ZN(n583) );
  INV_X1 U1124 ( .A(pmp_addr_i[253]), .ZN(n603) );
  NAND2_X1 U1125 ( .A1(n5154), .A2(n603), .ZN(n591) );
  OAI211_X1 U1126 ( .C1(n5094), .C2(pmp_addr_i[249]), .A(n583), .B(n591), .ZN(
        n512) );
  INV_X1 U1127 ( .A(pmp_addr_i[248]), .ZN(n513) );
  NAND2_X1 U1128 ( .A1(n210), .A2(n513), .ZN(n599) );
  INV_X1 U1129 ( .A(pmp_addr_i[247]), .ZN(n597) );
  NAND2_X1 U1130 ( .A1(n5202), .A2(n597), .ZN(n514) );
  NAND2_X1 U1131 ( .A1(n599), .A2(n514), .ZN(n602) );
  INV_X1 U1132 ( .A(pmp_addr_i[246]), .ZN(n515) );
  NAND2_X1 U1133 ( .A1(n5330), .A2(n515), .ZN(n596) );
  OAI21_X1 U1134 ( .B1(n5086), .B2(pmp_addr_i[245]), .A(n596), .ZN(n516) );
  NOR2_X1 U1135 ( .A1(n602), .A2(n516), .ZN(n568) );
  INV_X1 U1136 ( .A(pmp_addr_i[244]), .ZN(n517) );
  NAND2_X1 U1137 ( .A1(n12157), .A2(n517), .ZN(n575) );
  INV_X1 U1138 ( .A(pmp_addr_i[243]), .ZN(n574) );
  NAND2_X1 U1139 ( .A1(n3152), .A2(n574), .ZN(n518) );
  NAND2_X1 U1140 ( .A1(n575), .A2(n518), .ZN(n578) );
  INV_X1 U1141 ( .A(pmp_addr_i[242]), .ZN(n519) );
  NAND2_X1 U1142 ( .A1(instr_addr_o_20_), .A2(n519), .ZN(n572) );
  INV_X1 U1143 ( .A(pmp_addr_i[241]), .ZN(n571) );
  NAND2_X1 U1144 ( .A1(n3793), .A2(n571), .ZN(n520) );
  NAND2_X1 U1145 ( .A1(n572), .A2(n520), .ZN(n521) );
  NOR2_X1 U1146 ( .A1(n578), .A2(n521), .ZN(n522) );
  AND3_X1 U1147 ( .A1(n606), .A2(n568), .A3(n522), .ZN(n567) );
  NAND2_X1 U1148 ( .A1(n5250), .A2(n5389), .ZN(n539) );
  INV_X1 U1149 ( .A(pmp_addr_i[233]), .ZN(n523) );
  NOR2_X1 U1150 ( .A1(n5069), .A2(n523), .ZN(n525) );
  BUF_X1 U1151 ( .A(n679), .Z(n5070) );
  AOI22_X1 U1152 ( .A1(n525), .A2(n539), .B1(n5070), .B2(pmp_addr_i[234]), 
        .ZN(n531) );
  INV_X1 U1153 ( .A(pmp_addr_i[236]), .ZN(n526) );
  NAND2_X1 U1154 ( .A1(n4788), .A2(n526), .ZN(n529) );
  NAND2_X1 U1155 ( .A1(n150), .A2(n5390), .ZN(n527) );
  NAND2_X1 U1156 ( .A1(n529), .A2(n527), .ZN(n538) );
  NOR2_X1 U1157 ( .A1(n149), .A2(n5390), .ZN(n528) );
  AOI22_X1 U1158 ( .A1(n529), .A2(n528), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[236]), .ZN(n530) );
  OAI21_X1 U1159 ( .B1(n531), .B2(n538), .A(n530), .ZN(n532) );
  INV_X1 U1161 ( .A(n536), .ZN(n542) );
  INV_X1 U1162 ( .A(n538), .ZN(n540) );
  OAI211_X1 U1163 ( .C1(pmp_addr_i[233]), .C2(n5052), .A(n540), .B(n539), .ZN(
        n541) );
  NOR2_X1 U1164 ( .A1(n542), .A2(n541), .ZN(n566) );
  NOR2_X1 U1166 ( .A1(n155), .A2(n1741), .ZN(n546) );
  INV_X1 U1167 ( .A(pmp_addr_i[232]), .ZN(n544) );
  NAND2_X1 U1168 ( .A1(instr_addr_o_10_), .A2(n544), .ZN(n548) );
  BUF_X1 U1169 ( .A(n545), .Z(n5041) );
  AOI22_X1 U1170 ( .A1(n546), .A2(n548), .B1(n4602), .B2(pmp_addr_i[232]), 
        .ZN(n562) );
  NAND2_X1 U1171 ( .A1(instr_addr_o_9_), .A2(n1741), .ZN(n547) );
  NAND2_X1 U1172 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U1173 ( .A1(n562), .A2(n549), .ZN(n565) );
  BUF_X1 U1174 ( .A(n5031), .Z(n3839) );
  NAND2_X1 U1175 ( .A1(n12152), .A2(n453), .ZN(n554) );
  NOR2_X1 U1176 ( .A1(pmp_addr_i[225]), .A2(pmp_addr_i[224]), .ZN(n551) );
  INV_X1 U1177 ( .A(pmp_addr_i[226]), .ZN(n550) );
  AND2_X1 U1178 ( .A1(n551), .A2(n550), .ZN(n552) );
  OAI22_X1 U1179 ( .A1(n3836), .A2(n552), .B1(n551), .B2(n550), .ZN(n553) );
  NAND3_X1 U1180 ( .A1(n554), .A2(pmp_addr_i[227]), .A3(n3839), .ZN(n556) );
  NAND2_X1 U1182 ( .A1(n2611), .A2(pmp_addr_i[228]), .ZN(n555) );
  NAND2_X1 U1183 ( .A1(n205), .A2(n1752), .ZN(n560) );
  NAND2_X1 U1184 ( .A1(n5268), .A2(n473), .ZN(n557) );
  NAND3_X1 U1185 ( .A1(n558), .A2(n560), .A3(n557), .ZN(n563) );
  NOR2_X1 U1186 ( .A1(n5268), .A2(n473), .ZN(n559) );
  INV_X1 U1187 ( .A(n2623), .ZN(n4606) );
  AOI22_X1 U1188 ( .A1(n560), .A2(n559), .B1(n4606), .B2(pmp_addr_i[230]), 
        .ZN(n561) );
  NAND3_X1 U1189 ( .A1(n562), .A2(n563), .A3(n561), .ZN(n564) );
  INV_X1 U1190 ( .A(n568), .ZN(n570) );
  INV_X1 U1191 ( .A(n606), .ZN(n569) );
  NOR2_X1 U1192 ( .A1(n570), .A2(n569), .ZN(n593) );
  INV_X2 U1193 ( .A(n2339), .ZN(n5100) );
  NOR2_X1 U1194 ( .A1(n5100), .A2(n571), .ZN(n573) );
  BUF_X1 U1195 ( .A(n1996), .Z(n4631) );
  AOI22_X1 U1196 ( .A1(n573), .A2(n572), .B1(n4631), .B2(pmp_addr_i[242]), 
        .ZN(n579) );
  NOR2_X1 U1197 ( .A1(instr_addr_o_21_), .A2(n574), .ZN(n576) );
  AOI22_X1 U1199 ( .A1(n576), .A2(n575), .B1(n5192), .B2(pmp_addr_i[244]), 
        .ZN(n577) );
  OAI21_X1 U1200 ( .B1(n579), .B2(n578), .A(n577), .ZN(n592) );
  INV_X1 U1201 ( .A(n580), .ZN(n5162) );
  INV_X1 U1202 ( .A(pmp_addr_i[249]), .ZN(n581) );
  NOR2_X1 U1203 ( .A1(n5162), .A2(n581), .ZN(n582) );
  AOI22_X1 U1204 ( .A1(n583), .A2(n582), .B1(n4438), .B2(pmp_addr_i[250]), 
        .ZN(n589) );
  INV_X1 U1205 ( .A(pmp_addr_i[251]), .ZN(n584) );
  NOR2_X1 U1206 ( .A1(instr_addr_o_29_), .A2(n584), .ZN(n585) );
  AOI22_X1 U1208 ( .A1(n586), .A2(n585), .B1(n4658), .B2(pmp_addr_i[252]), 
        .ZN(n587) );
  OAI21_X1 U1209 ( .B1(n589), .B2(n588), .A(n587), .ZN(n590) );
  AOI22_X1 U1210 ( .A1(n593), .A2(n592), .B1(n591), .B2(n590), .ZN(n608) );
  INV_X1 U1211 ( .A(pmp_addr_i[245]), .ZN(n594) );
  NOR2_X1 U1212 ( .A1(n5208), .A2(n594), .ZN(n595) );
  BUF_X1 U1213 ( .A(n4135), .Z(n2580) );
  AOI22_X1 U1214 ( .A1(n596), .A2(n595), .B1(n2580), .B2(pmp_addr_i[246]), 
        .ZN(n601) );
  NOR2_X1 U1215 ( .A1(n137), .A2(n597), .ZN(n598) );
  BUF_X1 U1216 ( .A(n1026), .Z(n3806) );
  AOI22_X1 U1217 ( .A1(n599), .A2(n598), .B1(n3806), .B2(pmp_addr_i[248]), 
        .ZN(n600) );
  OAI21_X1 U1218 ( .B1(n602), .B2(n601), .A(n600), .ZN(n605) );
  INV_X1 U1219 ( .A(instr_addr_i[31]), .ZN(n3295) );
  NOR2_X1 U1220 ( .A1(pmp_addr_i[254]), .A2(pmp_addr_i[255]), .ZN(n7116) );
  OAI21_X1 U1221 ( .B1(n6018), .B2(n603), .A(n7116), .ZN(n604) );
  AOI21_X1 U1222 ( .B1(n606), .B2(n605), .A(n604), .ZN(n607) );
  INV_X1 U1223 ( .A(pmp_addr_i[171]), .ZN(n5239) );
  INV_X1 U1224 ( .A(pmp_cfg_i[51]), .ZN(n663) );
  NAND2_X1 U1225 ( .A1(pmp_addr_i[192]), .A2(pmp_addr_i[193]), .ZN(n651) );
  OR2_X1 U1226 ( .A1(n651), .A2(n657), .ZN(n4891) );
  NAND2_X1 U1227 ( .A1(n4842), .A2(pmp_addr_i[196]), .ZN(n11543) );
  OR2_X1 U1228 ( .A1(n11543), .A2(n667), .ZN(n11533) );
  INV_X1 U1229 ( .A(pmp_addr_i[198]), .ZN(n665) );
  OR2_X1 U1230 ( .A1(n11533), .A2(n665), .ZN(n11526) );
  AND2_X1 U1231 ( .A1(pmp_addr_i[199]), .A2(pmp_addr_i[200]), .ZN(n623) );
  NAND2_X1 U1232 ( .A1(n623), .A2(pmp_addr_i[201]), .ZN(n612) );
  NOR2_X1 U1233 ( .A1(n11526), .A2(n612), .ZN(n11521) );
  INV_X1 U1234 ( .A(pmp_cfg_i[52]), .ZN(n10596) );
  AOI21_X1 U1235 ( .B1(n11521), .B2(pmp_cfg_i[51]), .A(n10596), .ZN(n620) );
  NAND2_X1 U1236 ( .A1(pmp_addr_i[203]), .A2(pmp_addr_i[202]), .ZN(n613) );
  AND2_X1 U1237 ( .A1(n613), .A2(pmp_cfg_i[52]), .ZN(n614) );
  OR2_X1 U1238 ( .A1(n620), .A2(n614), .ZN(n617) );
  NAND2_X1 U1239 ( .A1(n617), .A2(pmp_addr_i[203]), .ZN(n615) );
  OAI21_X1 U1240 ( .B1(n5239), .B2(n4892), .A(n615), .ZN(n10517) );
  INV_X1 U1241 ( .A(n10517), .ZN(n4849) );
  NOR2_X1 U1242 ( .A1(n150), .A2(n4849), .ZN(n4871) );
  INV_X1 U1243 ( .A(pmp_addr_i[172]), .ZN(n5235) );
  NAND2_X1 U1244 ( .A1(n617), .A2(pmp_addr_i[204]), .ZN(n618) );
  OAI21_X1 U1245 ( .B1(n5235), .B2(n4892), .A(n618), .ZN(n10519) );
  NOR2_X1 U1246 ( .A1(n206), .A2(n10516), .ZN(n4865) );
  NOR2_X1 U1247 ( .A1(n4871), .A2(n4865), .ZN(n685) );
  INV_X1 U1248 ( .A(pmp_addr_i[170]), .ZN(n5243) );
  NAND2_X1 U1249 ( .A1(n620), .A2(pmp_addr_i[202]), .ZN(n619) );
  OAI21_X1 U1250 ( .B1(n5243), .B2(n4892), .A(n619), .ZN(n10506) );
  INV_X1 U1251 ( .A(n10506), .ZN(n10500) );
  OR2_X1 U1252 ( .A1(n5245), .A2(n10500), .ZN(n4861) );
  INV_X1 U1253 ( .A(pmp_addr_i[169]), .ZN(n5868) );
  NAND2_X1 U1254 ( .A1(n620), .A2(pmp_addr_i[201]), .ZN(n621) );
  OAI21_X1 U1255 ( .B1(n5868), .B2(n4892), .A(n621), .ZN(n10507) );
  INV_X1 U1256 ( .A(n10507), .ZN(n10498) );
  OR2_X1 U1257 ( .A1(instr_addr_o_11_), .A2(n10498), .ZN(n4869) );
  AND4_X1 U1258 ( .A1(pmp_addr_i[196]), .A2(pmp_addr_i[201]), .A3(
        pmp_addr_i[202]), .A4(pmp_addr_i[198]), .ZN(n622) );
  NAND4_X1 U1259 ( .A1(n4842), .A2(pmp_addr_i[197]), .A3(n623), .A4(n622), 
        .ZN(n11570) );
  INV_X1 U1260 ( .A(pmp_addr_i[203]), .ZN(n624) );
  NOR2_X1 U1261 ( .A1(n11570), .A2(n624), .ZN(n11561) );
  NAND2_X1 U1262 ( .A1(n11561), .A2(pmp_addr_i[204]), .ZN(n11522) );
  OR2_X1 U1263 ( .A1(n11522), .A2(n633), .ZN(n4883) );
  OR2_X1 U1264 ( .A1(n4883), .A2(n635), .ZN(n11564) );
  NAND2_X1 U1265 ( .A1(pmp_cfg_i[51]), .A2(pmp_addr_i[207]), .ZN(n625) );
  NAND2_X1 U1266 ( .A1(n878), .A2(pmp_addr_i[176]), .ZN(n626) );
  OAI21_X1 U1267 ( .B1(n4893), .B2(n627), .A(n626), .ZN(n10625) );
  INV_X1 U1268 ( .A(n10625), .ZN(n628) );
  NOR2_X1 U1269 ( .A1(n6019), .A2(n628), .ZN(n689) );
  NAND2_X1 U1270 ( .A1(n878), .A2(pmp_addr_i[175]), .ZN(n629) );
  OAI21_X1 U1271 ( .B1(n4893), .B2(n630), .A(n629), .ZN(n10527) );
  INV_X1 U1272 ( .A(n10527), .ZN(n4857) );
  NOR2_X1 U1273 ( .A1(n4069), .A2(n4857), .ZN(n631) );
  NOR2_X1 U1274 ( .A1(n689), .A2(n631), .ZN(n692) );
  OAI21_X1 U1275 ( .B1(n4883), .B2(n663), .A(pmp_cfg_i[52]), .ZN(n636) );
  NAND2_X1 U1276 ( .A1(n878), .A2(pmp_addr_i[173]), .ZN(n632) );
  OAI21_X1 U1277 ( .B1(n636), .B2(n633), .A(n632), .ZN(n10464) );
  INV_X1 U1278 ( .A(n10464), .ZN(n10658) );
  NOR2_X1 U1279 ( .A1(instr_addr_o_15_), .A2(n10658), .ZN(n4870) );
  NAND2_X1 U1280 ( .A1(n878), .A2(pmp_addr_i[174]), .ZN(n634) );
  OAI21_X1 U1281 ( .B1(n636), .B2(n635), .A(n634), .ZN(n11568) );
  INV_X1 U1282 ( .A(n11568), .ZN(n637) );
  NOR2_X1 U1283 ( .A1(n3100), .A2(n637), .ZN(n4860) );
  NOR2_X1 U1284 ( .A1(n4870), .A2(n4860), .ZN(n638) );
  NAND2_X1 U1285 ( .A1(n692), .A2(n638), .ZN(n694) );
  INV_X1 U1286 ( .A(pmp_addr_i[167]), .ZN(n5258) );
  INV_X1 U1287 ( .A(pmp_addr_i[199]), .ZN(n639) );
  NOR2_X1 U1288 ( .A1(n11526), .A2(n639), .ZN(n11530) );
  AOI21_X1 U1289 ( .B1(n11530), .B2(pmp_cfg_i[51]), .A(n10596), .ZN(n641) );
  NAND2_X1 U1290 ( .A1(n641), .A2(pmp_addr_i[199]), .ZN(n640) );
  OAI21_X1 U1291 ( .B1(n4892), .B2(n5258), .A(n640), .ZN(n10503) );
  INV_X1 U1292 ( .A(n10503), .ZN(n4848) );
  AND2_X1 U1293 ( .A1(n155), .A2(n4848), .ZN(n644) );
  INV_X1 U1294 ( .A(pmp_addr_i[168]), .ZN(n5867) );
  NAND2_X1 U1295 ( .A1(n641), .A2(pmp_addr_i[200]), .ZN(n642) );
  OAI21_X1 U1296 ( .B1(n4892), .B2(n5867), .A(n642), .ZN(n10502) );
  INV_X1 U1297 ( .A(n10502), .ZN(n643) );
  OR2_X1 U1298 ( .A1(n5262), .A2(n643), .ZN(n4853) );
  AOI22_X1 U1299 ( .A1(n644), .A2(n4853), .B1(n12202), .B2(n643), .ZN(n676) );
  NAND2_X1 U1300 ( .A1(n320), .A2(n4853), .ZN(n645) );
  NOR2_X1 U1301 ( .A1(n694), .A2(n646), .ZN(n678) );
  INV_X1 U1302 ( .A(pmp_addr_i[164]), .ZN(n648) );
  AOI21_X1 U1303 ( .B1(n4842), .B2(pmp_cfg_i[51]), .A(n10596), .ZN(n649) );
  NAND2_X1 U1304 ( .A1(n649), .A2(pmp_addr_i[196]), .ZN(n647) );
  OAI21_X1 U1305 ( .B1(n4892), .B2(n648), .A(n647), .ZN(n10484) );
  INV_X1 U1306 ( .A(n10484), .ZN(n10654) );
  NOR2_X1 U1307 ( .A1(n12152), .A2(n10654), .ZN(n4872) );
  INV_X1 U1308 ( .A(pmp_addr_i[163]), .ZN(n5859) );
  NAND2_X1 U1309 ( .A1(n649), .A2(pmp_addr_i[195]), .ZN(n650) );
  OAI21_X1 U1310 ( .B1(n4892), .B2(n5859), .A(n650), .ZN(n10485) );
  INV_X1 U1311 ( .A(n10485), .ZN(n10483) );
  NOR2_X1 U1312 ( .A1(n4596), .A2(n10483), .ZN(n4841) );
  OAI21_X1 U1313 ( .B1(n651), .B2(n663), .A(pmp_cfg_i[52]), .ZN(n658) );
  NAND2_X1 U1314 ( .A1(n878), .A2(pmp_addr_i[161]), .ZN(n652) );
  OAI21_X1 U1315 ( .B1(n658), .B2(n653), .A(n652), .ZN(n10474) );
  NAND2_X1 U1316 ( .A1(n878), .A2(pmp_addr_i[160]), .ZN(n655) );
  NAND2_X1 U1317 ( .A1(n663), .A2(pmp_addr_i[192]), .ZN(n654) );
  NAND2_X1 U1318 ( .A1(n655), .A2(n654), .ZN(n10652) );
  OR2_X1 U1319 ( .A1(n10474), .A2(n10652), .ZN(n659) );
  NAND2_X1 U1320 ( .A1(n878), .A2(pmp_addr_i[162]), .ZN(n656) );
  OAI21_X1 U1321 ( .B1(n658), .B2(n657), .A(n656), .ZN(n10478) );
  NAND2_X1 U1322 ( .A1(n659), .A2(n10478), .ZN(n660) );
  INV_X1 U1323 ( .A(n659), .ZN(n4894) );
  INV_X1 U1324 ( .A(n10478), .ZN(n10650) );
  AOI22_X1 U1325 ( .A1(n3836), .A2(n660), .B1(n4894), .B2(n10650), .ZN(n661)
         );
  NOR3_X1 U1326 ( .A1(n4872), .A2(n4841), .A3(n661), .ZN(n671) );
  NAND2_X1 U1327 ( .A1(n5293), .A2(n10483), .ZN(n662) );
  OAI22_X1 U1328 ( .A1(n4872), .A2(n662), .B1(n2611), .B2(n10484), .ZN(n670)
         );
  OAI21_X1 U1329 ( .B1(n11533), .B2(n663), .A(pmp_cfg_i[52]), .ZN(n668) );
  NAND2_X1 U1330 ( .A1(n878), .A2(pmp_addr_i[166]), .ZN(n664) );
  OAI21_X1 U1331 ( .B1(n668), .B2(n665), .A(n664), .ZN(n10491) );
  INV_X1 U1332 ( .A(n10491), .ZN(n672) );
  NOR2_X1 U1333 ( .A1(n5342), .A2(n672), .ZN(n673) );
  NAND2_X1 U1334 ( .A1(n878), .A2(pmp_addr_i[165]), .ZN(n666) );
  OAI21_X1 U1335 ( .B1(n668), .B2(n667), .A(n666), .ZN(n10492) );
  INV_X1 U1336 ( .A(n10492), .ZN(n4843) );
  NOR2_X1 U1337 ( .A1(n5268), .A2(n4843), .ZN(n669) );
  NOR2_X1 U1338 ( .A1(n673), .A2(n669), .ZN(n4886) );
  OAI21_X1 U1339 ( .B1(n671), .B2(n670), .A(n4886), .ZN(n677) );
  NAND2_X1 U1340 ( .A1(instr_addr_o_8_), .A2(n672), .ZN(n4833) );
  INV_X1 U1341 ( .A(n673), .ZN(n674) );
  NAND3_X1 U1342 ( .A1(n674), .A2(n5268), .A3(n4843), .ZN(n675) );
  INV_X1 U1343 ( .A(n4861), .ZN(n681) );
  NAND2_X1 U1344 ( .A1(instr_addr_o_11_), .A2(n10498), .ZN(n680) );
  OAI22_X1 U1345 ( .A1(n681), .A2(n680), .B1(n2733), .B2(n10506), .ZN(n684) );
  NAND2_X1 U1346 ( .A1(n149), .A2(n4849), .ZN(n682) );
  OAI22_X1 U1347 ( .A1(n4865), .A2(n682), .B1(instr_addr_o_14__BAR), .B2(
        n10519), .ZN(n683) );
  AOI21_X1 U1348 ( .B1(n685), .B2(n684), .A(n683), .ZN(n695) );
  NAND2_X1 U1349 ( .A1(n12179), .A2(n10658), .ZN(n686) );
  OAI22_X1 U1350 ( .A1(n4860), .A2(n686), .B1(n5058), .B2(n11568), .ZN(n691)
         );
  INV_X2 U1351 ( .A(n12228), .ZN(n5974) );
  NAND2_X1 U1352 ( .A1(n12265), .A2(n4857), .ZN(n688) );
  OAI22_X1 U1353 ( .A1(n689), .A2(n688), .B1(n1922), .B2(n10625), .ZN(n690) );
  AOI21_X1 U1354 ( .B1(n692), .B2(n691), .A(n690), .ZN(n693) );
  OAI21_X1 U1355 ( .B1(n695), .B2(n694), .A(n693), .ZN(n737) );
  NAND2_X1 U1356 ( .A1(n878), .A2(pmp_addr_i[184]), .ZN(n696) );
  OAI21_X1 U1357 ( .B1(n4893), .B2(n697), .A(n696), .ZN(n10605) );
  INV_X1 U1358 ( .A(n10605), .ZN(n698) );
  NOR2_X1 U1359 ( .A1(n210), .A2(n698), .ZN(n773) );
  NAND2_X1 U1360 ( .A1(n878), .A2(pmp_addr_i[183]), .ZN(n700) );
  OAI21_X1 U1361 ( .B1(n4893), .B2(n701), .A(n700), .ZN(n10613) );
  INV_X1 U1362 ( .A(n10613), .ZN(n771) );
  NOR2_X1 U1363 ( .A1(n5365), .A2(n771), .ZN(n702) );
  NAND2_X1 U1364 ( .A1(n878), .A2(pmp_addr_i[181]), .ZN(n703) );
  OAI21_X1 U1365 ( .B1(n4893), .B2(n704), .A(n703), .ZN(n10639) );
  INV_X1 U1366 ( .A(n10639), .ZN(n768) );
  NAND2_X1 U1367 ( .A1(n878), .A2(pmp_addr_i[182]), .ZN(n705) );
  OAI21_X1 U1368 ( .B1(n4893), .B2(n706), .A(n705), .ZN(n10628) );
  OR2_X1 U1369 ( .A1(n5330), .A2(n10558), .ZN(n767) );
  OAI21_X1 U1370 ( .B1(n5208), .B2(n768), .A(n767), .ZN(n707) );
  INV_X1 U1371 ( .A(n707), .ZN(n708) );
  INV_X1 U1373 ( .A(n739), .ZN(n721) );
  NAND2_X1 U1374 ( .A1(n878), .A2(pmp_addr_i[179]), .ZN(n709) );
  OAI21_X1 U1375 ( .B1(n4893), .B2(n710), .A(n709), .ZN(n10611) );
  INV_X1 U1376 ( .A(n10611), .ZN(n746) );
  NAND2_X1 U1377 ( .A1(n878), .A2(pmp_addr_i[180]), .ZN(n711) );
  OAI21_X1 U1378 ( .B1(n4893), .B2(n712), .A(n711), .ZN(n10637) );
  INV_X1 U1379 ( .A(n10637), .ZN(n713) );
  OR2_X1 U1380 ( .A1(n5181), .A2(n713), .ZN(n745) );
  OAI21_X1 U1381 ( .B1(n3152), .B2(n746), .A(n745), .ZN(n740) );
  NAND2_X1 U1382 ( .A1(n878), .A2(pmp_addr_i[177]), .ZN(n714) );
  OAI21_X1 U1383 ( .B1(n4893), .B2(n715), .A(n714), .ZN(n10626) );
  INV_X1 U1384 ( .A(n10626), .ZN(n742) );
  NAND2_X1 U1385 ( .A1(n878), .A2(pmp_addr_i[178]), .ZN(n716) );
  OAI21_X1 U1386 ( .B1(n4893), .B2(n717), .A(n716), .ZN(n10636) );
  INV_X1 U1387 ( .A(n10636), .ZN(n718) );
  OR2_X1 U1388 ( .A1(n5187), .A2(n718), .ZN(n741) );
  OAI21_X1 U1389 ( .B1(instr_addr_o_19_), .B2(n742), .A(n741), .ZN(n719) );
  NOR2_X1 U1390 ( .A1(n740), .A2(n719), .ZN(n720) );
  NAND2_X1 U1391 ( .A1(n721), .A2(n720), .ZN(n735) );
  NAND2_X1 U1392 ( .A1(n878), .A2(pmp_addr_i[188]), .ZN(n722) );
  OAI21_X1 U1393 ( .B1(n4893), .B2(n723), .A(n722), .ZN(n10623) );
  INV_X1 U1394 ( .A(n10623), .ZN(n724) );
  NOR2_X1 U1395 ( .A1(n4753), .A2(n724), .ZN(n758) );
  NAND2_X1 U1396 ( .A1(n878), .A2(pmp_addr_i[187]), .ZN(n725) );
  OAI21_X1 U1397 ( .B1(n4893), .B2(n726), .A(n725), .ZN(n10648) );
  INV_X1 U1398 ( .A(n10648), .ZN(n756) );
  NOR2_X1 U1399 ( .A1(instr_addr_o_29_), .A2(n756), .ZN(n727) );
  NOR2_X1 U1400 ( .A1(n758), .A2(n727), .ZN(n761) );
  INV_X1 U1401 ( .A(pmp_addr_i[189]), .ZN(n12073) );
  OR2_X1 U1402 ( .A1(n4893), .A2(n728), .ZN(n12092) );
  OAI21_X1 U1403 ( .B1(n4892), .B2(n12073), .A(n12092), .ZN(n10661) );
  NOR2_X1 U1404 ( .A1(pmp_addr_i[190]), .A2(pmp_addr_i[191]), .ZN(n5135) );
  INV_X1 U1405 ( .A(n5135), .ZN(n776) );
  AOI21_X1 U1406 ( .B1(n4660), .B2(n10661), .A(n776), .ZN(n762) );
  NAND2_X1 U1407 ( .A1(n878), .A2(pmp_addr_i[186]), .ZN(n729) );
  OAI21_X1 U1408 ( .B1(n4893), .B2(n730), .A(n729), .ZN(n10634) );
  INV_X1 U1409 ( .A(n10634), .ZN(n731) );
  OR2_X1 U1410 ( .A1(n5368), .A2(n731), .ZN(n752) );
  NAND2_X1 U1411 ( .A1(n878), .A2(pmp_addr_i[185]), .ZN(n732) );
  OAI21_X1 U1412 ( .B1(n4893), .B2(n733), .A(n732), .ZN(n10615) );
  NAND2_X1 U1413 ( .A1(n4652), .A2(n10615), .ZN(n734) );
  NAND4_X1 U1414 ( .A1(n761), .A2(n762), .A3(n752), .A4(n734), .ZN(n778) );
  NOR2_X1 U1415 ( .A1(n735), .A2(n778), .ZN(n736) );
  OAI21_X1 U1416 ( .B1(n738), .B2(n737), .A(n736), .ZN(n783) );
  OR2_X1 U1417 ( .A1(n778), .A2(n739), .ZN(n766) );
  INV_X1 U1418 ( .A(n740), .ZN(n751) );
  INV_X1 U1419 ( .A(n741), .ZN(n744) );
  NAND2_X1 U1420 ( .A1(instr_addr_o_19_), .A2(n742), .ZN(n743) );
  OAI22_X1 U1421 ( .A1(n744), .A2(n743), .B1(n2569), .B2(n10636), .ZN(n750) );
  INV_X1 U1422 ( .A(n745), .ZN(n748) );
  NAND2_X1 U1423 ( .A1(n3152), .A2(n746), .ZN(n747) );
  OAI22_X1 U1424 ( .A1(n748), .A2(n747), .B1(n999), .B2(n10637), .ZN(n749) );
  AOI21_X1 U1425 ( .B1(n751), .B2(n750), .A(n749), .ZN(n765) );
  INV_X1 U1426 ( .A(n752), .ZN(n755) );
  INV_X1 U1427 ( .A(n10615), .ZN(n753) );
  NAND2_X1 U1428 ( .A1(instr_addr_o_27_), .A2(n753), .ZN(n754) );
  OAI22_X1 U1429 ( .A1(n755), .A2(n754), .B1(n4438), .B2(n10634), .ZN(n760) );
  NAND2_X1 U1430 ( .A1(n5550), .A2(n756), .ZN(n757) );
  OAI22_X1 U1431 ( .A1(n758), .A2(n757), .B1(n5115), .B2(n10623), .ZN(n759) );
  AOI21_X1 U1432 ( .B1(n761), .B2(n760), .A(n759), .ZN(n764) );
  INV_X1 U1433 ( .A(n762), .ZN(n763) );
  OAI22_X1 U1434 ( .A1(n766), .A2(n765), .B1(n764), .B2(n763), .ZN(n781) );
  INV_X1 U1435 ( .A(n767), .ZN(n770) );
  NAND2_X1 U1436 ( .A1(n5208), .A2(n768), .ZN(n769) );
  OAI22_X1 U1437 ( .A1(n770), .A2(n769), .B1(n1269), .B2(n10628), .ZN(n775) );
  NAND2_X1 U1438 ( .A1(n12226), .A2(n771), .ZN(n772) );
  OAI22_X1 U1439 ( .A1(n773), .A2(n772), .B1(n1273), .B2(n10605), .ZN(n774) );
  AOI21_X1 U1440 ( .B1(n169), .B2(n775), .A(n774), .ZN(n779) );
  NAND3_X1 U1441 ( .A1(n4866), .A2(n10580), .A3(n5135), .ZN(n777) );
  OAI21_X1 U1442 ( .B1(n779), .B2(n778), .A(n777), .ZN(n780) );
  NOR2_X1 U1443 ( .A1(n781), .A2(n780), .ZN(n782) );
  BUF_X1 U1444 ( .A(n207), .Z(n6017) );
  NAND2_X1 U1445 ( .A1(n5047), .A2(n627), .ZN(n797) );
  NAND2_X1 U1446 ( .A1(n5974), .A2(n630), .ZN(n784) );
  AND2_X1 U1447 ( .A1(n797), .A2(n784), .ZN(n795) );
  NAND2_X1 U1448 ( .A1(n5226), .A2(n635), .ZN(n794) );
  OAI211_X1 U1449 ( .C1(pmp_addr_i[205]), .C2(n6017), .A(n795), .B(n794), .ZN(
        n823) );
  INV_X1 U1450 ( .A(n823), .ZN(n803) );
  INV_X1 U1451 ( .A(pmp_addr_i[202]), .ZN(n785) );
  NAND2_X1 U1452 ( .A1(n5250), .A2(n785), .ZN(n820) );
  NOR2_X1 U1453 ( .A1(n5069), .A2(n423), .ZN(n786) );
  AOI22_X1 U1454 ( .A1(n820), .A2(n786), .B1(n5070), .B2(pmp_addr_i[202]), 
        .ZN(n792) );
  NAND2_X1 U1455 ( .A1(n5251), .A2(n415), .ZN(n789) );
  NAND2_X1 U1456 ( .A1(n150), .A2(n624), .ZN(n787) );
  AND2_X1 U1457 ( .A1(n789), .A2(n787), .ZN(n821) );
  INV_X1 U1458 ( .A(n821), .ZN(n791) );
  NOR2_X1 U1459 ( .A1(n150), .A2(n624), .ZN(n788) );
  AOI22_X1 U1460 ( .A1(n789), .A2(n788), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[204]), .ZN(n790) );
  OAI21_X1 U1461 ( .B1(n792), .B2(n791), .A(n790), .ZN(n802) );
  NOR2_X1 U1462 ( .A1(instr_addr_o_15_), .A2(n633), .ZN(n793) );
  AOI22_X1 U1463 ( .A1(n794), .A2(n793), .B1(n5058), .B2(pmp_addr_i[206]), 
        .ZN(n800) );
  INV_X1 U1464 ( .A(n795), .ZN(n799) );
  NOR2_X1 U1465 ( .A1(n5062), .A2(n630), .ZN(n796) );
  AOI22_X1 U1466 ( .A1(n797), .A2(n796), .B1(n2082), .B2(pmp_addr_i[208]), 
        .ZN(n798) );
  OAI21_X1 U1467 ( .B1(n800), .B2(n799), .A(n798), .ZN(n801) );
  AOI21_X1 U1468 ( .B1(n803), .B2(n802), .A(n801), .ZN(n842) );
  INV_X1 U1469 ( .A(pmp_addr_i[196]), .ZN(n804) );
  NAND2_X1 U1470 ( .A1(instr_addr_o_6_), .A2(n804), .ZN(n810) );
  NOR2_X1 U1471 ( .A1(n4596), .A2(n611), .ZN(n805) );
  AOI22_X1 U1472 ( .A1(n810), .A2(n805), .B1(n2611), .B2(pmp_addr_i[196]), 
        .ZN(n814) );
  OR2_X1 U1473 ( .A1(pmp_addr_i[193]), .A2(pmp_addr_i[192]), .ZN(n806) );
  NOR2_X1 U1474 ( .A1(n806), .A2(pmp_addr_i[194]), .ZN(n808) );
  INV_X1 U1475 ( .A(n806), .ZN(n807) );
  OAI22_X1 U1476 ( .A1(n5899), .A2(n808), .B1(n807), .B2(n657), .ZN(n809) );
  OAI211_X1 U1477 ( .C1(pmp_addr_i[195]), .C2(n5031), .A(n810), .B(n809), .ZN(
        n813) );
  BUF_X1 U1478 ( .A(n2424), .Z(n3844) );
  NAND2_X1 U1479 ( .A1(n205), .A2(n665), .ZN(n817) );
  OAI21_X1 U1480 ( .B1(n3844), .B2(pmp_addr_i[197]), .A(n817), .ZN(n812) );
  AOI21_X1 U1481 ( .B1(n814), .B2(n813), .A(n812), .ZN(n831) );
  NOR2_X1 U1482 ( .A1(n154), .A2(n639), .ZN(n816) );
  INV_X1 U1483 ( .A(pmp_addr_i[200]), .ZN(n815) );
  NAND2_X1 U1484 ( .A1(n5270), .A2(n815), .ZN(n825) );
  AOI22_X1 U1485 ( .A1(n816), .A2(n825), .B1(n4602), .B2(pmp_addr_i[200]), 
        .ZN(n827) );
  NAND3_X1 U1486 ( .A1(n817), .A2(n3844), .A3(pmp_addr_i[197]), .ZN(n819) );
  NAND2_X1 U1487 ( .A1(n3894), .A2(pmp_addr_i[198]), .ZN(n818) );
  NAND3_X1 U1488 ( .A1(n827), .A2(n819), .A3(n818), .ZN(n830) );
  OAI211_X1 U1489 ( .C1(pmp_addr_i[201]), .C2(n5052), .A(n821), .B(n820), .ZN(
        n822) );
  NOR2_X1 U1490 ( .A1(n823), .A2(n822), .ZN(n829) );
  NAND2_X1 U1491 ( .A1(n154), .A2(n639), .ZN(n824) );
  NAND2_X1 U1492 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U1493 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U1495 ( .A1(n12161), .A2(n723), .ZN(n864) );
  OAI21_X1 U1496 ( .B1(n4656), .B2(pmp_addr_i[219]), .A(n864), .ZN(n866) );
  NAND2_X1 U1497 ( .A1(instr_addr_o_28_), .A2(n730), .ZN(n862) );
  NOR2_X1 U1500 ( .A1(n866), .A2(n832), .ZN(n860) );
  NAND2_X1 U1501 ( .A1(n4802), .A2(n717), .ZN(n843) );
  NAND2_X1 U1502 ( .A1(n3793), .A2(n715), .ZN(n833) );
  AND2_X1 U1503 ( .A1(n843), .A2(n833), .ZN(n839) );
  NAND2_X1 U1504 ( .A1(n210), .A2(n697), .ZN(n855) );
  NAND2_X1 U1505 ( .A1(n5202), .A2(n701), .ZN(n834) );
  NAND2_X1 U1506 ( .A1(n855), .A2(n834), .ZN(n858) );
  NAND2_X1 U1507 ( .A1(n6028), .A2(n706), .ZN(n853) );
  OAI21_X1 U1508 ( .B1(n5086), .B2(pmp_addr_i[213]), .A(n853), .ZN(n835) );
  NOR2_X1 U1509 ( .A1(n858), .A2(n835), .ZN(n851) );
  NAND2_X1 U1510 ( .A1(n3152), .A2(n710), .ZN(n836) );
  NAND2_X1 U1511 ( .A1(n12157), .A2(n712), .ZN(n845) );
  NAND2_X1 U1512 ( .A1(n836), .A2(n845), .ZN(n848) );
  INV_X1 U1513 ( .A(n848), .ZN(n837) );
  NAND3_X1 U1514 ( .A1(n860), .A2(n839), .A3(n838), .ZN(n840) );
  NOR2_X1 U1516 ( .A1(n5100), .A2(n715), .ZN(n844) );
  AOI22_X1 U1517 ( .A1(n844), .A2(n843), .B1(n2569), .B2(pmp_addr_i[210]), 
        .ZN(n849) );
  NOR2_X1 U1518 ( .A1(n5842), .A2(n710), .ZN(n846) );
  AOI22_X1 U1519 ( .A1(n846), .A2(n845), .B1(n5192), .B2(pmp_addr_i[212]), 
        .ZN(n847) );
  OAI21_X1 U1520 ( .B1(n849), .B2(n848), .A(n847), .ZN(n850) );
  NAND3_X1 U1521 ( .A1(n860), .A2(n851), .A3(n850), .ZN(n874) );
  NOR2_X1 U1522 ( .A1(n5208), .A2(n704), .ZN(n852) );
  AOI22_X1 U1523 ( .A1(n853), .A2(n852), .B1(n1269), .B2(pmp_addr_i[214]), 
        .ZN(n857) );
  NOR2_X1 U1524 ( .A1(n5365), .A2(n701), .ZN(n854) );
  AOI22_X1 U1525 ( .A1(n855), .A2(n854), .B1(n1273), .B2(pmp_addr_i[216]), 
        .ZN(n856) );
  OAI21_X1 U1526 ( .B1(n858), .B2(n857), .A(n856), .ZN(n859) );
  NAND2_X1 U1527 ( .A1(n860), .A2(n859), .ZN(n873) );
  NOR2_X1 U1528 ( .A1(n5162), .A2(n733), .ZN(n861) );
  AOI22_X1 U1529 ( .A1(n862), .A2(n861), .B1(n4438), .B2(pmp_addr_i[218]), 
        .ZN(n867) );
  NOR2_X1 U1530 ( .A1(instr_addr_o_29_), .A2(n726), .ZN(n863) );
  AOI22_X1 U1531 ( .A1(n864), .A2(n863), .B1(n5115), .B2(pmp_addr_i[220]), 
        .ZN(n865) );
  OAI21_X1 U1532 ( .B1(n867), .B2(n866), .A(n865), .ZN(n869) );
  NAND2_X1 U1533 ( .A1(n869), .A2(n868), .ZN(n872) );
  OAI21_X1 U1534 ( .B1(n6018), .B2(n728), .A(n10453), .ZN(n870) );
  INV_X1 U1535 ( .A(n870), .ZN(n871) );
  NAND4_X1 U1536 ( .A1(n874), .A2(n873), .A3(n872), .A4(n871), .ZN(n875) );
  OR2_X1 U1537 ( .A1(n876), .A2(n875), .ZN(n877) );
  INV_X1 U1538 ( .A(pmp_cfg_i[83]), .ZN(n11659) );
  INV_X1 U1539 ( .A(n9329), .ZN(n984) );
  INV_X1 U1540 ( .A(pmp_addr_i[304]), .ZN(n883) );
  NAND2_X1 U1541 ( .A1(pmp_addr_i[323]), .A2(pmp_addr_i[324]), .ZN(n911) );
  NAND2_X1 U1542 ( .A1(pmp_addr_i[326]), .A2(pmp_addr_i[325]), .ZN(n879) );
  OR2_X1 U1543 ( .A1(n911), .A2(n879), .ZN(n11642) );
  INV_X1 U1544 ( .A(pmp_addr_i[327]), .ZN(n2963) );
  NOR2_X1 U1545 ( .A1(n11642), .A2(n2963), .ZN(n3350) );
  AND2_X1 U1546 ( .A1(pmp_addr_i[330]), .A2(pmp_addr_i[329]), .ZN(n3351) );
  NAND3_X1 U1547 ( .A1(n3350), .A2(pmp_addr_i[328]), .A3(n3351), .ZN(n896) );
  AND2_X1 U1548 ( .A1(pmp_addr_i[320]), .A2(pmp_addr_i[321]), .ZN(n3373) );
  NAND4_X1 U1549 ( .A1(n3373), .A2(pmp_addr_i[322]), .A3(pmp_addr_i[332]), 
        .A4(pmp_addr_i[331]), .ZN(n880) );
  OR2_X1 U1550 ( .A1(n896), .A2(n880), .ZN(n11648) );
  INV_X1 U1551 ( .A(pmp_addr_i[333]), .ZN(n887) );
  NOR2_X1 U1552 ( .A1(n11648), .A2(n887), .ZN(n3366) );
  NAND2_X1 U1553 ( .A1(n3366), .A2(pmp_addr_i[334]), .ZN(n11689) );
  INV_X1 U1554 ( .A(pmp_addr_i[335]), .ZN(n2999) );
  OAI21_X1 U1555 ( .B1(n11689), .B2(n2999), .A(pmp_cfg_i[84]), .ZN(n881) );
  NAND2_X1 U1556 ( .A1(n881), .A2(pmp_cfg_i[83]), .ZN(n3374) );
  NAND2_X1 U1557 ( .A1(n3374), .A2(pmp_addr_i[336]), .ZN(n882) );
  OAI21_X1 U1558 ( .B1(n984), .B2(n883), .A(n882), .ZN(n9199) );
  INV_X1 U1559 ( .A(n9199), .ZN(n884) );
  INV_X1 U1560 ( .A(pmp_addr_i[303]), .ZN(n886) );
  NAND2_X1 U1561 ( .A1(n3374), .A2(pmp_addr_i[335]), .ZN(n885) );
  OAI21_X1 U1562 ( .B1(n984), .B2(n886), .A(n885), .ZN(n9045) );
  INV_X1 U1563 ( .A(n9045), .ZN(n9077) );
  OR2_X1 U1564 ( .A1(n943), .A2(n3322), .ZN(n942) );
  OAI21_X1 U1565 ( .B1(n11648), .B2(n11659), .A(pmp_cfg_i[84]), .ZN(n900) );
  INV_X1 U1566 ( .A(pmp_addr_i[301]), .ZN(n5434) );
  OAI22_X1 U1567 ( .A1(n900), .A2(n887), .B1(n5434), .B2(n984), .ZN(n9197) );
  INV_X1 U1568 ( .A(n9197), .ZN(n9062) );
  NOR2_X1 U1569 ( .A1(n5057), .A2(n9062), .ZN(n3313) );
  NAND2_X1 U1570 ( .A1(pmp_cfg_i[84]), .A2(pmp_addr_i[334]), .ZN(n888) );
  AOI21_X1 U1571 ( .B1(n3366), .B2(pmp_cfg_i[83]), .A(n888), .ZN(n890) );
  AND2_X1 U1572 ( .A1(n9329), .A2(pmp_addr_i[302]), .ZN(n889) );
  OR2_X1 U1573 ( .A1(n890), .A2(n889), .ZN(n11681) );
  INV_X1 U1574 ( .A(n11681), .ZN(n9057) );
  OR2_X1 U1575 ( .A1(n3313), .A2(n3320), .ZN(n891) );
  NOR2_X1 U1576 ( .A1(n942), .A2(n891), .ZN(n941) );
  NAND3_X1 U1577 ( .A1(n3373), .A2(pmp_addr_i[322]), .A3(pmp_cfg_i[83]), .ZN(
        n925) );
  OAI21_X1 U1578 ( .B1(n925), .B2(n11642), .A(pmp_cfg_i[84]), .ZN(n910) );
  NAND2_X1 U1579 ( .A1(n9329), .A2(pmp_addr_i[295]), .ZN(n892) );
  OAI21_X1 U1580 ( .B1(n910), .B2(n2963), .A(n892), .ZN(n9229) );
  INV_X1 U1581 ( .A(n9229), .ZN(n9070) );
  NAND2_X1 U1582 ( .A1(instr_addr_o_9_), .A2(n9070), .ZN(n3383) );
  INV_X1 U1583 ( .A(pmp_addr_i[296]), .ZN(n894) );
  INV_X1 U1584 ( .A(pmp_cfg_i[84]), .ZN(n901) );
  OAI21_X1 U1585 ( .B1(pmp_addr_i[327]), .B2(n901), .A(n910), .ZN(n903) );
  NAND2_X1 U1586 ( .A1(n903), .A2(pmp_addr_i[328]), .ZN(n893) );
  OAI21_X1 U1587 ( .B1(n984), .B2(n894), .A(n893), .ZN(n9230) );
  INV_X1 U1588 ( .A(n9230), .ZN(n9074) );
  NOR2_X1 U1589 ( .A1(n214), .A2(n9074), .ZN(n3329) );
  NAND2_X1 U1590 ( .A1(n5270), .A2(n9074), .ZN(n3387) );
  OAI21_X1 U1591 ( .B1(n3383), .B2(n3329), .A(n3387), .ZN(n915) );
  NOR2_X1 U1592 ( .A1(n5040), .A2(n9070), .ZN(n3315) );
  NOR2_X1 U1593 ( .A1(n3315), .A2(n3329), .ZN(n895) );
  OAI21_X1 U1594 ( .B1(n896), .B2(n925), .A(pmp_cfg_i[84]), .ZN(n907) );
  INV_X1 U1595 ( .A(pmp_addr_i[331]), .ZN(n897) );
  INV_X1 U1596 ( .A(pmp_addr_i[299]), .ZN(n2229) );
  OAI22_X1 U1597 ( .A1(n907), .A2(n897), .B1(n2229), .B2(n984), .ZN(n9206) );
  INV_X1 U1598 ( .A(n9206), .ZN(n9063) );
  NOR2_X1 U1599 ( .A1(n150), .A2(n9063), .ZN(n3342) );
  INV_X1 U1600 ( .A(pmp_addr_i[332]), .ZN(n899) );
  NAND2_X1 U1601 ( .A1(n9329), .A2(pmp_addr_i[300]), .ZN(n898) );
  OAI21_X1 U1602 ( .B1(n900), .B2(n899), .A(n898), .ZN(n9207) );
  INV_X1 U1603 ( .A(n9207), .ZN(n9065) );
  NOR2_X1 U1604 ( .A1(n206), .A2(n9065), .ZN(n3309) );
  NOR2_X1 U1605 ( .A1(n3342), .A2(n3309), .ZN(n940) );
  INV_X1 U1606 ( .A(pmp_addr_i[297]), .ZN(n2139) );
  NOR2_X1 U1607 ( .A1(n901), .A2(pmp_addr_i[328]), .ZN(n902) );
  OAI21_X1 U1608 ( .B1(n903), .B2(n902), .A(pmp_addr_i[329]), .ZN(n904) );
  OAI21_X1 U1609 ( .B1(n984), .B2(n2139), .A(n904), .ZN(n9203) );
  INV_X1 U1610 ( .A(n9203), .ZN(n9073) );
  NOR2_X1 U1611 ( .A1(n4493), .A2(n9073), .ZN(n3308) );
  INV_X1 U1612 ( .A(pmp_addr_i[330]), .ZN(n906) );
  NAND2_X1 U1613 ( .A1(n9329), .A2(pmp_addr_i[298]), .ZN(n905) );
  OAI21_X1 U1614 ( .B1(n907), .B2(n906), .A(n905), .ZN(n9204) );
  INV_X1 U1615 ( .A(n9204), .ZN(n9072) );
  NOR2_X1 U1616 ( .A1(n3308), .A2(n3321), .ZN(n908) );
  INV_X1 U1617 ( .A(pmp_addr_i[326]), .ZN(n2954) );
  NAND2_X1 U1618 ( .A1(n9329), .A2(pmp_addr_i[294]), .ZN(n909) );
  OAI21_X1 U1619 ( .B1(n910), .B2(n2954), .A(n909), .ZN(n9226) );
  INV_X1 U1620 ( .A(n9226), .ZN(n9075) );
  OR2_X1 U1621 ( .A1(n5342), .A2(n9075), .ZN(n3323) );
  INV_X1 U1622 ( .A(n3323), .ZN(n913) );
  OAI21_X1 U1623 ( .B1(n925), .B2(n911), .A(pmp_cfg_i[84]), .ZN(n917) );
  INV_X1 U1624 ( .A(pmp_addr_i[325]), .ZN(n2957) );
  NAND2_X1 U1625 ( .A1(n9329), .A2(pmp_addr_i[293]), .ZN(n912) );
  OAI21_X1 U1626 ( .B1(n917), .B2(n2957), .A(n912), .ZN(n9227) );
  INV_X1 U1627 ( .A(n9227), .ZN(n9058) );
  NAND2_X1 U1628 ( .A1(n5740), .A2(n9058), .ZN(n3381) );
  NAND2_X1 U1629 ( .A1(n5342), .A2(n9075), .ZN(n3395) );
  OAI21_X1 U1630 ( .B1(n913), .B2(n3381), .A(n3395), .ZN(n914) );
  NOR2_X1 U1631 ( .A1(n915), .A2(n914), .ZN(n934) );
  INV_X1 U1632 ( .A(pmp_addr_i[324]), .ZN(n2933) );
  NAND2_X1 U1633 ( .A1(n9329), .A2(pmp_addr_i[292]), .ZN(n916) );
  OAI21_X1 U1634 ( .B1(n917), .B2(n2933), .A(n916), .ZN(n9220) );
  INV_X1 U1635 ( .A(n9220), .ZN(n9071) );
  NOR2_X1 U1636 ( .A1(n12152), .A2(n9071), .ZN(n3314) );
  NAND3_X1 U1637 ( .A1(n925), .A2(pmp_cfg_i[84]), .A3(pmp_addr_i[323]), .ZN(
        n919) );
  NAND2_X1 U1638 ( .A1(n9329), .A2(pmp_addr_i[291]), .ZN(n918) );
  NAND2_X1 U1639 ( .A1(n919), .A2(n918), .ZN(n9221) );
  INV_X1 U1640 ( .A(n9221), .ZN(n9034) );
  NOR2_X1 U1641 ( .A1(n4596), .A2(n9034), .ZN(n3330) );
  AND2_X1 U1642 ( .A1(pmp_cfg_i[83]), .A2(pmp_addr_i[320]), .ZN(n922) );
  NAND2_X1 U1643 ( .A1(pmp_cfg_i[84]), .A2(pmp_addr_i[321]), .ZN(n921) );
  NAND2_X1 U1644 ( .A1(n9329), .A2(pmp_addr_i[289]), .ZN(n920) );
  OAI21_X1 U1645 ( .B1(n922), .B2(n921), .A(n920), .ZN(n9213) );
  NAND2_X1 U1646 ( .A1(n9329), .A2(pmp_addr_i[288]), .ZN(n924) );
  NAND2_X1 U1647 ( .A1(n11659), .A2(pmp_addr_i[320]), .ZN(n923) );
  NAND2_X1 U1648 ( .A1(n924), .A2(n923), .ZN(n9212) );
  OR2_X1 U1649 ( .A1(n9213), .A2(n9212), .ZN(n928) );
  NAND3_X1 U1650 ( .A1(n925), .A2(pmp_cfg_i[84]), .A3(pmp_addr_i[322]), .ZN(
        n927) );
  NAND2_X1 U1651 ( .A1(n9329), .A2(pmp_addr_i[290]), .ZN(n926) );
  NAND2_X1 U1652 ( .A1(n927), .A2(n926), .ZN(n9217) );
  NAND2_X1 U1653 ( .A1(n928), .A2(n9217), .ZN(n929) );
  INV_X1 U1654 ( .A(n9217), .ZN(n9059) );
  INV_X1 U1655 ( .A(n928), .ZN(n3340) );
  AOI22_X1 U1656 ( .A1(n3836), .A2(n929), .B1(n9059), .B2(n3340), .ZN(n930) );
  NOR3_X1 U1657 ( .A1(n3314), .A2(n3330), .A3(n930), .ZN(n932) );
  NAND2_X1 U1658 ( .A1(n5293), .A2(n9034), .ZN(n3386) );
  NAND2_X1 U1659 ( .A1(n5277), .A2(n9071), .ZN(n3382) );
  OAI21_X1 U1660 ( .B1(n3314), .B2(n3386), .A(n3382), .ZN(n931) );
  OR2_X1 U1661 ( .A1(n12267), .A2(n9058), .ZN(n3316) );
  OAI211_X1 U1662 ( .C1(n932), .C2(n931), .A(n3316), .B(n3323), .ZN(n933) );
  AND2_X1 U1663 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1664 ( .A1(n936), .A2(n935), .ZN(n990) );
  NAND2_X1 U1665 ( .A1(instr_addr_o_11_), .A2(n9073), .ZN(n3397) );
  NAND2_X1 U1666 ( .A1(n5250), .A2(n9072), .ZN(n3389) );
  OAI21_X1 U1667 ( .B1(n3321), .B2(n3397), .A(n3389), .ZN(n939) );
  NAND2_X1 U1668 ( .A1(n4061), .A2(n9063), .ZN(n3390) );
  NAND2_X1 U1669 ( .A1(n4788), .A2(n9065), .ZN(n3396) );
  OAI21_X1 U1670 ( .B1(n3309), .B2(n3390), .A(n3396), .ZN(n938) );
  AOI21_X1 U1671 ( .B1(n940), .B2(n939), .A(n938), .ZN(n949) );
  INV_X1 U1672 ( .A(n941), .ZN(n948) );
  INV_X1 U1673 ( .A(n942), .ZN(n946) );
  NAND2_X1 U1674 ( .A1(n208), .A2(n9062), .ZN(n3384) );
  NAND2_X1 U1675 ( .A1(n5226), .A2(n9057), .ZN(n3394) );
  OAI21_X1 U1676 ( .B1(n3384), .B2(n3320), .A(n3394), .ZN(n945) );
  NAND2_X1 U1677 ( .A1(n5974), .A2(n9077), .ZN(n3388) );
  OAI22_X1 U1678 ( .A1(n943), .A2(n3388), .B1(n1922), .B2(n9199), .ZN(n944) );
  AOI21_X1 U1679 ( .B1(n946), .B2(n945), .A(n944), .ZN(n947) );
  OAI21_X1 U1680 ( .B1(n949), .B2(n948), .A(n947), .ZN(n989) );
  NAND2_X1 U1681 ( .A1(n3374), .A2(pmp_addr_i[344]), .ZN(n950) );
  OAI21_X1 U1682 ( .B1(n984), .B2(n2341), .A(n950), .ZN(n9264) );
  INV_X1 U1683 ( .A(n9264), .ZN(n951) );
  NOR2_X1 U1684 ( .A1(n12158), .A2(n951), .ZN(n1028) );
  NAND2_X1 U1685 ( .A1(n3374), .A2(pmp_addr_i[343]), .ZN(n952) );
  OAI21_X1 U1686 ( .B1(n984), .B2(n2374), .A(n952), .ZN(n9263) );
  INV_X1 U1687 ( .A(n9263), .ZN(n1025) );
  NOR2_X1 U1688 ( .A1(n5202), .A2(n1025), .ZN(n953) );
  OR2_X1 U1689 ( .A1(n1028), .A2(n953), .ZN(n1020) );
  INV_X1 U1690 ( .A(pmp_addr_i[309]), .ZN(n955) );
  NAND2_X1 U1691 ( .A1(n3374), .A2(pmp_addr_i[341]), .ZN(n954) );
  OAI21_X1 U1692 ( .B1(n984), .B2(n955), .A(n954), .ZN(n9260) );
  INV_X1 U1693 ( .A(n9260), .ZN(n1022) );
  INV_X1 U1694 ( .A(pmp_addr_i[310]), .ZN(n957) );
  NAND2_X1 U1695 ( .A1(n3374), .A2(pmp_addr_i[342]), .ZN(n956) );
  OAI21_X1 U1696 ( .B1(n984), .B2(n957), .A(n956), .ZN(n9261) );
  INV_X1 U1697 ( .A(n9261), .ZN(n958) );
  OR2_X1 U1698 ( .A1(n5330), .A2(n958), .ZN(n1021) );
  OAI21_X1 U1699 ( .B1(instr_addr_o_23_), .B2(n1022), .A(n1021), .ZN(n959) );
  NOR2_X1 U1700 ( .A1(n1020), .A2(n959), .ZN(n991) );
  INV_X1 U1701 ( .A(pmp_addr_i[307]), .ZN(n961) );
  NAND2_X1 U1702 ( .A1(n3374), .A2(pmp_addr_i[339]), .ZN(n960) );
  OAI21_X1 U1703 ( .B1(n984), .B2(n961), .A(n960), .ZN(n9267) );
  INV_X1 U1704 ( .A(n9267), .ZN(n998) );
  INV_X1 U1705 ( .A(pmp_addr_i[308]), .ZN(n963) );
  NAND2_X1 U1706 ( .A1(n3374), .A2(pmp_addr_i[340]), .ZN(n962) );
  OAI21_X1 U1707 ( .B1(n984), .B2(n963), .A(n962), .ZN(n9268) );
  INV_X1 U1708 ( .A(n9268), .ZN(n964) );
  OR2_X1 U1709 ( .A1(n5181), .A2(n964), .ZN(n997) );
  OAI21_X1 U1710 ( .B1(n3152), .B2(n998), .A(n997), .ZN(n992) );
  INV_X1 U1711 ( .A(pmp_addr_i[305]), .ZN(n966) );
  NAND2_X1 U1712 ( .A1(n3374), .A2(pmp_addr_i[337]), .ZN(n965) );
  OAI21_X1 U1713 ( .B1(n984), .B2(n966), .A(n965), .ZN(n9270) );
  INV_X1 U1714 ( .A(n9270), .ZN(n994) );
  INV_X1 U1715 ( .A(pmp_addr_i[306]), .ZN(n968) );
  NAND2_X1 U1716 ( .A1(n3374), .A2(pmp_addr_i[338]), .ZN(n967) );
  OAI21_X1 U1717 ( .B1(n984), .B2(n968), .A(n967), .ZN(n9271) );
  INV_X1 U1718 ( .A(n9271), .ZN(n969) );
  OR2_X1 U1719 ( .A1(n5187), .A2(n969), .ZN(n993) );
  OAI21_X1 U1720 ( .B1(n5100), .B2(n994), .A(n993), .ZN(n970) );
  NOR2_X1 U1721 ( .A1(n992), .A2(n970), .ZN(n971) );
  NAND2_X1 U1722 ( .A1(n991), .A2(n971), .ZN(n987) );
  INV_X1 U1723 ( .A(pmp_addr_i[316]), .ZN(n973) );
  NAND2_X1 U1724 ( .A1(n3374), .A2(pmp_addr_i[348]), .ZN(n972) );
  OAI21_X1 U1725 ( .B1(n984), .B2(n973), .A(n972), .ZN(n9279) );
  INV_X1 U1726 ( .A(n9279), .ZN(n974) );
  NOR2_X1 U1727 ( .A1(n4560), .A2(n974), .ZN(n1011) );
  INV_X1 U1728 ( .A(pmp_addr_i[315]), .ZN(n976) );
  NAND2_X1 U1729 ( .A1(n3374), .A2(pmp_addr_i[347]), .ZN(n975) );
  OAI21_X1 U1730 ( .B1(n984), .B2(n976), .A(n975), .ZN(n9278) );
  INV_X1 U1731 ( .A(n9278), .ZN(n1009) );
  NOR2_X1 U1732 ( .A1(instr_addr_o_29_), .A2(n1009), .ZN(n977) );
  NOR2_X1 U1733 ( .A1(n1011), .A2(n977), .ZN(n1014) );
  INV_X1 U1734 ( .A(pmp_addr_i[314]), .ZN(n979) );
  NAND2_X1 U1735 ( .A1(n3374), .A2(pmp_addr_i[346]), .ZN(n978) );
  OAI21_X1 U1736 ( .B1(n984), .B2(n979), .A(n978), .ZN(n9276) );
  INV_X1 U1737 ( .A(n9276), .ZN(n980) );
  OR2_X1 U1738 ( .A1(n5368), .A2(n980), .ZN(n1005) );
  INV_X1 U1739 ( .A(pmp_addr_i[313]), .ZN(n982) );
  NAND2_X1 U1740 ( .A1(n3374), .A2(pmp_addr_i[345]), .ZN(n981) );
  OAI21_X1 U1741 ( .B1(n984), .B2(n982), .A(n981), .ZN(n9275) );
  NAND2_X1 U1742 ( .A1(n4652), .A2(n9275), .ZN(n986) );
  INV_X1 U1743 ( .A(pmp_addr_i[317]), .ZN(n983) );
  NAND2_X1 U1744 ( .A1(n3374), .A2(pmp_addr_i[349]), .ZN(n12099) );
  OAI21_X1 U1745 ( .B1(n984), .B2(n983), .A(n12099), .ZN(n9282) );
  INV_X1 U1746 ( .A(pmp_addr_i[319]), .ZN(n985) );
  OR2_X1 U1747 ( .A1(pmp_addr_i[319]), .A2(pmp_addr_i[318]), .ZN(n1032) );
  AOI21_X1 U1748 ( .B1(n4005), .B2(n9282), .A(n1032), .ZN(n1015) );
  NAND2_X1 U1749 ( .A1(n1014), .A2(n333), .ZN(n1036) );
  NOR2_X1 U1750 ( .A1(n987), .A2(n1036), .ZN(n988) );
  NAND2_X1 U1751 ( .A1(n202), .A2(n991), .ZN(n1019) );
  INV_X1 U1752 ( .A(n992), .ZN(n1004) );
  INV_X1 U1753 ( .A(n993), .ZN(n996) );
  NAND2_X1 U1754 ( .A1(n3793), .A2(n994), .ZN(n995) );
  OAI22_X1 U1755 ( .A1(n996), .A2(n995), .B1(n2569), .B2(n9271), .ZN(n1003) );
  INV_X1 U1756 ( .A(n997), .ZN(n1001) );
  NAND2_X1 U1757 ( .A1(n3152), .A2(n998), .ZN(n1000) );
  OAI22_X1 U1758 ( .A1(n1001), .A2(n1000), .B1(n999), .B2(n9268), .ZN(n1002)
         );
  AOI21_X1 U1759 ( .B1(n1004), .B2(n1003), .A(n1002), .ZN(n1018) );
  INV_X1 U1760 ( .A(n1005), .ZN(n1008) );
  INV_X1 U1761 ( .A(n9275), .ZN(n1006) );
  NAND2_X1 U1762 ( .A1(instr_addr_o_27_), .A2(n1006), .ZN(n1007) );
  OAI22_X1 U1763 ( .A1(n1008), .A2(n1007), .B1(n4438), .B2(n9276), .ZN(n1013)
         );
  NAND2_X1 U1764 ( .A1(instr_addr_o_29_), .A2(n1009), .ZN(n1010) );
  OAI22_X1 U1765 ( .A1(n1011), .A2(n1010), .B1(n4658), .B2(n9279), .ZN(n1012)
         );
  AOI21_X1 U1766 ( .B1(n1014), .B2(n1013), .A(n1012), .ZN(n1017) );
  INV_X1 U1767 ( .A(n1015), .ZN(n1016) );
  OAI22_X1 U1768 ( .A1(n1018), .A2(n1019), .B1(n1017), .B2(n1016), .ZN(n1039)
         );
  INV_X1 U1769 ( .A(n1020), .ZN(n1031) );
  INV_X1 U1770 ( .A(n1021), .ZN(n1024) );
  NAND2_X1 U1771 ( .A1(n5208), .A2(n1022), .ZN(n1023) );
  OAI22_X1 U1772 ( .A1(n1024), .A2(n1023), .B1(n1269), .B2(n9261), .ZN(n1030)
         );
  NAND2_X1 U1773 ( .A1(n5202), .A2(n1025), .ZN(n1027) );
  OAI22_X1 U1774 ( .A1(n1028), .A2(n1027), .B1(n1273), .B2(n9264), .ZN(n1029)
         );
  AOI21_X1 U1775 ( .B1(n1031), .B2(n1030), .A(n1029), .ZN(n1037) );
  INV_X1 U1776 ( .A(n9282), .ZN(n1034) );
  INV_X1 U1777 ( .A(n1032), .ZN(n1033) );
  NAND3_X1 U1778 ( .A1(n6018), .A2(n1034), .A3(n1033), .ZN(n1035) );
  OAI21_X1 U1779 ( .B1(n1037), .B2(n1036), .A(n1035), .ZN(n1038) );
  NOR2_X1 U1780 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NAND2_X1 U1781 ( .A1(n5245), .A2(n906), .ZN(n1073) );
  INV_X1 U1782 ( .A(pmp_addr_i[329]), .ZN(n1041) );
  NOR2_X1 U1783 ( .A1(n5069), .A2(n1041), .ZN(n1042) );
  AOI22_X1 U1784 ( .A1(n1073), .A2(n1042), .B1(n5070), .B2(pmp_addr_i[330]), 
        .ZN(n1047) );
  NAND2_X1 U1785 ( .A1(n4788), .A2(n899), .ZN(n1045) );
  NAND2_X1 U1786 ( .A1(n4061), .A2(n897), .ZN(n1043) );
  NAND2_X1 U1787 ( .A1(n1045), .A2(n1043), .ZN(n1072) );
  NOR2_X1 U1788 ( .A1(n149), .A2(n897), .ZN(n1044) );
  AOI22_X1 U1789 ( .A1(n1045), .A2(n1044), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[332]), .ZN(n1046) );
  OAI21_X1 U1790 ( .B1(n1047), .B2(n1072), .A(n1046), .ZN(n1070) );
  INV_X1 U1791 ( .A(pmp_addr_i[334]), .ZN(n1048) );
  NAND2_X1 U1792 ( .A1(n5226), .A2(n1048), .ZN(n1067) );
  NOR2_X1 U1793 ( .A1(n208), .A2(n887), .ZN(n1049) );
  AOI22_X1 U1794 ( .A1(n1067), .A2(n1049), .B1(n5058), .B2(pmp_addr_i[334]), 
        .ZN(n1054) );
  INV_X1 U1795 ( .A(pmp_addr_i[336]), .ZN(n1050) );
  NAND2_X1 U1796 ( .A1(n6019), .A2(n1050), .ZN(n1052) );
  OAI21_X1 U1797 ( .B1(n5048), .B2(pmp_addr_i[335]), .A(n1052), .ZN(n1069) );
  NOR2_X1 U1798 ( .A1(n12156), .A2(n2999), .ZN(n1051) );
  AOI22_X1 U1799 ( .A1(n1052), .A2(n1051), .B1(n2750), .B2(pmp_addr_i[336]), 
        .ZN(n1053) );
  INV_X1 U1800 ( .A(pmp_addr_i[348]), .ZN(n1055) );
  NAND2_X1 U1801 ( .A1(n12161), .A2(n1055), .ZN(n1119) );
  OAI21_X1 U1802 ( .B1(n4656), .B2(pmp_addr_i[347]), .A(n1119), .ZN(n1121) );
  BUF_X1 U1803 ( .A(n4000), .Z(n4147) );
  INV_X1 U1804 ( .A(pmp_addr_i[349]), .ZN(n1138) );
  NAND2_X1 U1805 ( .A1(n5154), .A2(n1138), .ZN(n1124) );
  INV_X1 U1806 ( .A(pmp_addr_i[344]), .ZN(n1057) );
  NAND2_X1 U1807 ( .A1(n12158), .A2(n1057), .ZN(n1133) );
  INV_X1 U1808 ( .A(pmp_addr_i[343]), .ZN(n1130) );
  NAND2_X1 U1809 ( .A1(n5202), .A2(n1130), .ZN(n1058) );
  NAND2_X1 U1810 ( .A1(n1133), .A2(n1058), .ZN(n1136) );
  INV_X1 U1811 ( .A(pmp_addr_i[342]), .ZN(n1059) );
  NAND2_X1 U1812 ( .A1(n4835), .A2(n1059), .ZN(n1129) );
  OAI21_X1 U1813 ( .B1(n5086), .B2(pmp_addr_i[341]), .A(n1129), .ZN(n1060) );
  NOR2_X1 U1814 ( .A1(n1136), .A2(n1060), .ZN(n1102) );
  INV_X1 U1815 ( .A(pmp_addr_i[340]), .ZN(n1061) );
  NAND2_X1 U1816 ( .A1(n12157), .A2(n1061), .ZN(n1109) );
  INV_X1 U1817 ( .A(pmp_addr_i[339]), .ZN(n1108) );
  NAND2_X1 U1818 ( .A1(n3152), .A2(n1108), .ZN(n1062) );
  NAND2_X1 U1819 ( .A1(n1109), .A2(n1062), .ZN(n1112) );
  INV_X1 U1820 ( .A(pmp_addr_i[338]), .ZN(n1063) );
  NAND2_X1 U1821 ( .A1(n6027), .A2(n1063), .ZN(n1106) );
  INV_X1 U1822 ( .A(pmp_addr_i[337]), .ZN(n1105) );
  NAND2_X1 U1823 ( .A1(n3793), .A2(n1105), .ZN(n1064) );
  NAND2_X1 U1824 ( .A1(n1106), .A2(n1064), .ZN(n1065) );
  NOR2_X1 U1825 ( .A1(n1112), .A2(n1065), .ZN(n1066) );
  AND3_X1 U1826 ( .A1(n1102), .A2(n1141), .A3(n1066), .ZN(n1101) );
  OAI21_X1 U1827 ( .B1(n4578), .B2(pmp_addr_i[333]), .A(n1067), .ZN(n1068) );
  NOR2_X1 U1828 ( .A1(n1069), .A2(n1068), .ZN(n1071) );
  INV_X1 U1829 ( .A(n1071), .ZN(n1076) );
  INV_X1 U1830 ( .A(n1072), .ZN(n1074) );
  OAI211_X1 U1831 ( .C1(pmp_addr_i[329]), .C2(n5052), .A(n1074), .B(n1073), 
        .ZN(n1075) );
  NOR2_X1 U1832 ( .A1(n1076), .A2(n1075), .ZN(n1100) );
  NOR2_X1 U1833 ( .A1(n154), .A2(n2963), .ZN(n1078) );
  INV_X1 U1834 ( .A(pmp_addr_i[328]), .ZN(n1077) );
  NAND2_X1 U1835 ( .A1(instr_addr_o_10_), .A2(n1077), .ZN(n1080) );
  AOI22_X1 U1836 ( .A1(n1078), .A2(n1080), .B1(n4602), .B2(pmp_addr_i[328]), 
        .ZN(n1096) );
  NAND2_X1 U1837 ( .A1(instr_addr_o_9_), .A2(n2963), .ZN(n1079) );
  NAND2_X1 U1838 ( .A1(n1080), .A2(n1079), .ZN(n1081) );
  NAND2_X1 U1839 ( .A1(n1096), .A2(n1081), .ZN(n1099) );
  NAND2_X1 U1840 ( .A1(n12152), .A2(n2933), .ZN(n1087) );
  OR2_X1 U1841 ( .A1(pmp_addr_i[321]), .A2(pmp_addr_i[320]), .ZN(n1082) );
  NOR2_X1 U1842 ( .A1(n1082), .A2(pmp_addr_i[322]), .ZN(n1085) );
  INV_X1 U1843 ( .A(n1082), .ZN(n1084) );
  INV_X1 U1844 ( .A(pmp_addr_i[322]), .ZN(n1083) );
  OAI22_X1 U1845 ( .A1(n3836), .A2(n1085), .B1(n1084), .B2(n1083), .ZN(n1086)
         );
  OAI211_X1 U1846 ( .C1(pmp_addr_i[323]), .C2(n3839), .A(n1087), .B(n1086), 
        .ZN(n1090) );
  NAND3_X1 U1847 ( .A1(n1087), .A2(pmp_addr_i[323]), .A3(n3839), .ZN(n1089) );
  NAND2_X1 U1848 ( .A1(n2611), .A2(pmp_addr_i[324]), .ZN(n1088) );
  NAND3_X1 U1849 ( .A1(n1090), .A2(n1089), .A3(n1088), .ZN(n1092) );
  NAND2_X1 U1850 ( .A1(n5342), .A2(n2954), .ZN(n1094) );
  NAND2_X1 U1851 ( .A1(n5268), .A2(n2957), .ZN(n1091) );
  NAND3_X1 U1852 ( .A1(n1092), .A2(n1094), .A3(n1091), .ZN(n1097) );
  NOR2_X1 U1853 ( .A1(n5268), .A2(n2957), .ZN(n1093) );
  AOI22_X1 U1854 ( .A1(n1094), .A2(n1093), .B1(n4606), .B2(pmp_addr_i[326]), 
        .ZN(n1095) );
  NAND3_X1 U1855 ( .A1(n1097), .A2(n1096), .A3(n1095), .ZN(n1098) );
  NAND4_X1 U1856 ( .A1(n1101), .A2(n1100), .A3(n1099), .A4(n1098), .ZN(n1144)
         );
  INV_X1 U1857 ( .A(n1102), .ZN(n1104) );
  INV_X1 U1858 ( .A(n1141), .ZN(n1103) );
  NOR2_X1 U1859 ( .A1(n1104), .A2(n1103), .ZN(n1126) );
  NOR2_X1 U1860 ( .A1(n5100), .A2(n1105), .ZN(n1107) );
  AOI22_X1 U1861 ( .A1(n1107), .A2(n1106), .B1(n4631), .B2(pmp_addr_i[338]), 
        .ZN(n1113) );
  NOR2_X1 U1862 ( .A1(instr_addr_o_21_), .A2(n1108), .ZN(n1110) );
  AOI22_X1 U1863 ( .A1(n1110), .A2(n1109), .B1(n999), .B2(pmp_addr_i[340]), 
        .ZN(n1111) );
  OAI21_X1 U1864 ( .B1(n1113), .B2(n1112), .A(n1111), .ZN(n1125) );
  INV_X1 U1865 ( .A(pmp_addr_i[345]), .ZN(n1114) );
  NOR2_X1 U1866 ( .A1(n5162), .A2(n1114), .ZN(n1115) );
  AOI22_X1 U1867 ( .A1(n1116), .A2(n1115), .B1(n5111), .B2(pmp_addr_i[346]), 
        .ZN(n1122) );
  INV_X1 U1868 ( .A(pmp_addr_i[347]), .ZN(n1117) );
  NOR2_X1 U1869 ( .A1(instr_addr_o_29_), .A2(n1117), .ZN(n1118) );
  AOI22_X1 U1870 ( .A1(n1119), .A2(n1118), .B1(n5115), .B2(pmp_addr_i[348]), 
        .ZN(n1120) );
  OAI21_X1 U1871 ( .B1(n1122), .B2(n1121), .A(n1120), .ZN(n1123) );
  AOI22_X1 U1872 ( .A1(n1126), .A2(n1125), .B1(n1124), .B2(n1123), .ZN(n1143)
         );
  INV_X1 U1873 ( .A(pmp_addr_i[341]), .ZN(n1127) );
  NOR2_X1 U1874 ( .A1(n5208), .A2(n1127), .ZN(n1128) );
  AOI22_X1 U1875 ( .A1(n1129), .A2(n1128), .B1(n2580), .B2(pmp_addr_i[342]), 
        .ZN(n1135) );
  NOR2_X1 U1876 ( .A1(n5365), .A2(n1130), .ZN(n1132) );
  AOI22_X1 U1877 ( .A1(n1133), .A2(n1132), .B1(n3806), .B2(pmp_addr_i[344]), 
        .ZN(n1134) );
  OAI21_X1 U1878 ( .B1(n1136), .B2(n1135), .A(n1134), .ZN(n1140) );
  NOR2_X1 U1879 ( .A1(pmp_addr_i[350]), .A2(pmp_addr_i[351]), .ZN(n1137) );
  OAI21_X1 U1880 ( .B1(n4866), .B2(n1138), .A(n1137), .ZN(n1139) );
  AOI21_X1 U1881 ( .B1(n1141), .B2(n1140), .A(n1139), .ZN(n1142) );
  NAND4_X1 U1882 ( .A1(n1145), .A2(n1144), .A3(n1143), .A4(n1142), .ZN(n1146)
         );
  INV_X1 U1883 ( .A(pmp_cfg_i[35]), .ZN(n1215) );
  INV_X1 U1884 ( .A(pmp_addr_i[103]), .ZN(n4782) );
  NAND2_X1 U1885 ( .A1(pmp_addr_i[128]), .A2(pmp_addr_i[129]), .ZN(n11910) );
  INV_X1 U1886 ( .A(pmp_addr_i[130]), .ZN(n1226) );
  OR2_X1 U1887 ( .A1(n11910), .A2(n1226), .ZN(n11897) );
  INV_X1 U1888 ( .A(pmp_addr_i[131]), .ZN(n1223) );
  NOR2_X1 U1889 ( .A1(n11897), .A2(n1223), .ZN(n11901) );
  NAND2_X1 U1890 ( .A1(n11901), .A2(pmp_addr_i[132]), .ZN(n11904) );
  INV_X1 U1891 ( .A(pmp_addr_i[133]), .ZN(n5267) );
  OR2_X1 U1892 ( .A1(n11904), .A2(n5267), .ZN(n11916) );
  INV_X1 U1893 ( .A(pmp_addr_i[134]), .ZN(n1148) );
  NOR2_X1 U1894 ( .A1(n11916), .A2(n1148), .ZN(n5591) );
  INV_X1 U1895 ( .A(pmp_cfg_i[36]), .ZN(n1216) );
  AOI21_X1 U1896 ( .B1(n5591), .B2(pmp_cfg_i[35]), .A(n1216), .ZN(n1219) );
  NAND2_X1 U1897 ( .A1(n1219), .A2(pmp_addr_i[135]), .ZN(n1149) );
  OAI21_X1 U1898 ( .B1(n1150), .B2(n4782), .A(n1149), .ZN(n9490) );
  INV_X1 U1899 ( .A(n9490), .ZN(n9649) );
  NOR2_X1 U1900 ( .A1(n4204), .A2(n9649), .ZN(n5537) );
  NAND2_X1 U1901 ( .A1(n5591), .A2(pmp_addr_i[135]), .ZN(n11921) );
  INV_X1 U1902 ( .A(pmp_addr_i[136]), .ZN(n5261) );
  OR2_X1 U1903 ( .A1(n11921), .A2(n5261), .ZN(n11929) );
  OAI21_X1 U1904 ( .B1(n11929), .B2(n1215), .A(pmp_cfg_i[36]), .ZN(n1211) );
  NAND2_X1 U1905 ( .A1(n9584), .A2(pmp_addr_i[104]), .ZN(n1151) );
  OAI21_X1 U1906 ( .B1(n1211), .B2(n5261), .A(n1151), .ZN(n9495) );
  INV_X1 U1907 ( .A(n9495), .ZN(n1152) );
  NOR2_X1 U1908 ( .A1(instr_addr_o_10_), .A2(n1152), .ZN(n5530) );
  NOR2_X1 U1909 ( .A1(n5537), .A2(n5530), .ZN(n1214) );
  NAND2_X1 U1910 ( .A1(n154), .A2(n9649), .ZN(n5603) );
  NAND2_X1 U1911 ( .A1(n12202), .A2(n1152), .ZN(n5614) );
  INV_X1 U1913 ( .A(pmp_addr_i[122]), .ZN(n1155) );
  INV_X1 U1914 ( .A(pmp_addr_i[137]), .ZN(n5249) );
  OR2_X1 U1915 ( .A1(n11929), .A2(n5249), .ZN(n5587) );
  AND2_X1 U1916 ( .A1(pmp_addr_i[140]), .A2(pmp_addr_i[139]), .ZN(n1198) );
  AND2_X1 U1917 ( .A1(n1198), .A2(pmp_addr_i[141]), .ZN(n5578) );
  NAND4_X1 U1918 ( .A1(n5578), .A2(pmp_addr_i[138]), .A3(pmp_addr_i[142]), 
        .A4(pmp_addr_i[143]), .ZN(n1153) );
  AND2_X1 U1919 ( .A1(pmp_cfg_i[35]), .A2(pmp_cfg_i[36]), .ZN(n11907) );
  OR2_X1 U1921 ( .A1(n1216), .A2(pmp_cfg_i[35]), .ZN(n9638) );
  NAND2_X1 U1922 ( .A1(n5567), .A2(n9638), .ZN(n5546) );
  NAND2_X1 U1923 ( .A1(n12224), .A2(pmp_addr_i[154]), .ZN(n1154) );
  OAI21_X1 U1924 ( .B1(n1150), .B2(n1155), .A(n1154), .ZN(n9619) );
  INV_X1 U1925 ( .A(n9619), .ZN(n1156) );
  OR2_X1 U1926 ( .A1(n5368), .A2(n1156), .ZN(n1252) );
  INV_X1 U1927 ( .A(pmp_addr_i[121]), .ZN(n1158) );
  NAND2_X1 U1928 ( .A1(n12225), .A2(pmp_addr_i[153]), .ZN(n1157) );
  OAI21_X1 U1929 ( .B1(n1150), .B2(n1158), .A(n1157), .ZN(n9586) );
  NAND2_X1 U1930 ( .A1(n4652), .A2(n9586), .ZN(n1159) );
  NAND2_X1 U1931 ( .A1(n12225), .A2(pmp_addr_i[157]), .ZN(n11943) );
  OAI21_X1 U1932 ( .B1(n1150), .B2(n4407), .A(n11943), .ZN(n9635) );
  NOR2_X1 U1933 ( .A1(pmp_addr_i[126]), .A2(pmp_addr_i[127]), .ZN(n4444) );
  AOI21_X1 U1934 ( .B1(n4005), .B2(n9635), .A(n197), .ZN(n1261) );
  INV_X1 U1935 ( .A(pmp_addr_i[124]), .ZN(n1161) );
  NAND2_X1 U1936 ( .A1(n5546), .A2(pmp_addr_i[156]), .ZN(n1160) );
  OAI21_X1 U1937 ( .B1(n1150), .B2(n1161), .A(n1160), .ZN(n9597) );
  INV_X1 U1938 ( .A(n9597), .ZN(n1162) );
  NOR2_X1 U1939 ( .A1(n12263), .A2(n1162), .ZN(n1258) );
  INV_X1 U1940 ( .A(pmp_addr_i[123]), .ZN(n1164) );
  NAND2_X1 U1941 ( .A1(n5546), .A2(pmp_addr_i[155]), .ZN(n1163) );
  OAI21_X1 U1942 ( .B1(n1150), .B2(n1164), .A(n1163), .ZN(n9632) );
  INV_X1 U1943 ( .A(n9632), .ZN(n1256) );
  NOR2_X1 U1944 ( .A1(n5149), .A2(n1256), .ZN(n1165) );
  INV_X1 U1945 ( .A(n1280), .ZN(n1191) );
  INV_X1 U1946 ( .A(pmp_addr_i[115]), .ZN(n1167) );
  NAND2_X1 U1947 ( .A1(n5546), .A2(pmp_addr_i[147]), .ZN(n1166) );
  OAI21_X1 U1948 ( .B1(n1150), .B2(n1167), .A(n1166), .ZN(n9625) );
  NOR2_X1 U1949 ( .A1(n5842), .A2(n9528), .ZN(n1171) );
  INV_X1 U1950 ( .A(pmp_addr_i[116]), .ZN(n1169) );
  NAND2_X1 U1951 ( .A1(n5546), .A2(pmp_addr_i[148]), .ZN(n1168) );
  OAI21_X1 U1952 ( .B1(n1150), .B2(n1169), .A(n1168), .ZN(n9624) );
  INV_X1 U1953 ( .A(n9624), .ZN(n1170) );
  NOR2_X1 U1954 ( .A1(n5181), .A2(n1170), .ZN(n1248) );
  INV_X1 U1955 ( .A(pmp_addr_i[113]), .ZN(n1173) );
  NAND2_X1 U1956 ( .A1(n12225), .A2(pmp_addr_i[145]), .ZN(n1172) );
  OAI21_X1 U1957 ( .B1(n1150), .B2(n1173), .A(n1172), .ZN(n9595) );
  INV_X1 U1958 ( .A(n9595), .ZN(n1244) );
  INV_X1 U1959 ( .A(pmp_addr_i[114]), .ZN(n1175) );
  NAND2_X1 U1960 ( .A1(n12224), .A2(pmp_addr_i[146]), .ZN(n1174) );
  OAI21_X1 U1961 ( .B1(n1150), .B2(n1175), .A(n1174), .ZN(n9588) );
  INV_X1 U1962 ( .A(n9588), .ZN(n1176) );
  NOR2_X1 U1963 ( .A1(n5187), .A2(n1176), .ZN(n1246) );
  INV_X1 U1964 ( .A(n1246), .ZN(n1177) );
  OAI21_X1 U1965 ( .B1(n5100), .B2(n1244), .A(n1177), .ZN(n1178) );
  NOR2_X1 U1966 ( .A1(n1243), .A2(n1178), .ZN(n1190) );
  INV_X1 U1967 ( .A(pmp_addr_i[117]), .ZN(n1180) );
  NAND2_X1 U1968 ( .A1(n12225), .A2(pmp_addr_i[149]), .ZN(n1179) );
  OAI21_X1 U1969 ( .B1(n1150), .B2(n1180), .A(n1179), .ZN(n9594) );
  INV_X1 U1970 ( .A(n9594), .ZN(n1268) );
  INV_X1 U1971 ( .A(pmp_addr_i[119]), .ZN(n1182) );
  NAND2_X1 U1972 ( .A1(n12224), .A2(pmp_addr_i[151]), .ZN(n1181) );
  OAI21_X1 U1973 ( .B1(n1150), .B2(n1182), .A(n1181), .ZN(n9618) );
  INV_X1 U1974 ( .A(n9618), .ZN(n1272) );
  NOR2_X1 U1975 ( .A1(n4644), .A2(n1272), .ZN(n1186) );
  INV_X1 U1976 ( .A(pmp_addr_i[120]), .ZN(n1184) );
  NAND2_X1 U1977 ( .A1(n12225), .A2(pmp_addr_i[152]), .ZN(n1183) );
  OAI21_X1 U1978 ( .B1(n1150), .B2(n1184), .A(n1183), .ZN(n9589) );
  INV_X1 U1979 ( .A(n9589), .ZN(n1185) );
  NOR2_X1 U1980 ( .A1(instr_addr_o_26_), .A2(n1185), .ZN(n1275) );
  INV_X1 U1981 ( .A(pmp_addr_i[118]), .ZN(n1188) );
  NAND2_X1 U1982 ( .A1(n12224), .A2(pmp_addr_i[150]), .ZN(n1187) );
  OAI21_X1 U1983 ( .B1(n1150), .B2(n1188), .A(n1187), .ZN(n9587) );
  OR2_X1 U1984 ( .A1(n6028), .A2(n9553), .ZN(n1267) );
  OAI211_X1 U1985 ( .C1(instr_addr_o_23_), .C2(n1268), .A(n1266), .B(n1267), 
        .ZN(n1242) );
  INV_X1 U1986 ( .A(n1242), .ZN(n1189) );
  INV_X1 U1987 ( .A(pmp_addr_i[112]), .ZN(n1193) );
  NAND2_X1 U1988 ( .A1(n12225), .A2(pmp_addr_i[144]), .ZN(n1192) );
  OAI21_X1 U1989 ( .B1(n1150), .B2(n1193), .A(n1192), .ZN(n9596) );
  INV_X1 U1990 ( .A(n9596), .ZN(n1194) );
  NOR2_X1 U1991 ( .A1(n6019), .A2(n1194), .ZN(n1295) );
  INV_X1 U1992 ( .A(pmp_addr_i[111]), .ZN(n1196) );
  NAND2_X1 U1993 ( .A1(n12224), .A2(pmp_addr_i[143]), .ZN(n1195) );
  OAI21_X1 U1994 ( .B1(n1150), .B2(n1196), .A(n1195), .ZN(n9519) );
  INV_X1 U1995 ( .A(n9519), .ZN(n1294) );
  NOR2_X1 U1996 ( .A1(n12265), .A2(n1294), .ZN(n5529) );
  NOR2_X1 U1997 ( .A1(n1295), .A2(n5529), .ZN(n1298) );
  INV_X1 U1998 ( .A(pmp_addr_i[109]), .ZN(n1200) );
  NAND2_X1 U1999 ( .A1(pmp_cfg_i[35]), .A2(pmp_addr_i[138]), .ZN(n1197) );
  OAI21_X1 U2000 ( .B1(n5587), .B2(n1197), .A(pmp_cfg_i[36]), .ZN(n1210) );
  OAI21_X1 U2001 ( .B1(n1198), .B2(n1216), .A(n1210), .ZN(n1206) );
  NAND2_X1 U2002 ( .A1(n1206), .A2(pmp_addr_i[141]), .ZN(n1199) );
  OAI21_X1 U2003 ( .B1(n1200), .B2(n1150), .A(n1199), .ZN(n9617) );
  INV_X1 U2004 ( .A(n9617), .ZN(n1292) );
  NOR2_X1 U2005 ( .A1(n5057), .A2(n1292), .ZN(n5549) );
  OR2_X1 U2006 ( .A1(n5578), .A2(n1216), .ZN(n1201) );
  INV_X1 U2007 ( .A(pmp_addr_i[142]), .ZN(n5225) );
  AOI21_X1 U2008 ( .B1(n1210), .B2(n1201), .A(n5225), .ZN(n1203) );
  INV_X1 U2009 ( .A(pmp_addr_i[110]), .ZN(n4767) );
  NOR2_X1 U2010 ( .A1(n1150), .A2(n4767), .ZN(n1202) );
  OR2_X1 U2011 ( .A1(n1203), .A2(n1202), .ZN(n11883) );
  INV_X1 U2012 ( .A(n11883), .ZN(n1293) );
  NOR2_X1 U2013 ( .A1(n3100), .A2(n1293), .ZN(n5525) );
  NOR2_X1 U2014 ( .A1(n5549), .A2(n5525), .ZN(n1204) );
  NAND2_X1 U2015 ( .A1(n1298), .A2(n1204), .ZN(n1300) );
  INV_X1 U2016 ( .A(pmp_addr_i[139]), .ZN(n5569) );
  NAND2_X1 U2017 ( .A1(n9584), .A2(pmp_addr_i[107]), .ZN(n1205) );
  OAI21_X1 U2018 ( .B1(n1210), .B2(n5569), .A(n1205), .ZN(n9604) );
  INV_X1 U2019 ( .A(n9604), .ZN(n1287) );
  NOR2_X1 U2020 ( .A1(n150), .A2(n1287), .ZN(n5536) );
  INV_X1 U2021 ( .A(pmp_addr_i[108]), .ZN(n1208) );
  NAND2_X1 U2022 ( .A1(n1206), .A2(pmp_addr_i[140]), .ZN(n1207) );
  OAI21_X1 U2023 ( .B1(n1150), .B2(n1208), .A(n1207), .ZN(n9616) );
  INV_X1 U2024 ( .A(n9616), .ZN(n1288) );
  NOR2_X1 U2025 ( .A1(n206), .A2(n1288), .ZN(n5519) );
  NOR2_X1 U2026 ( .A1(n5536), .A2(n5519), .ZN(n1291) );
  NAND2_X1 U2027 ( .A1(n9584), .A2(pmp_addr_i[106]), .ZN(n1209) );
  OAI21_X1 U2028 ( .B1(n1210), .B2(n1325), .A(n1209), .ZN(n9605) );
  INV_X1 U2029 ( .A(n9605), .ZN(n1285) );
  INV_X1 U2030 ( .A(pmp_addr_i[105]), .ZN(n4771) );
  OAI22_X1 U2031 ( .A1(n1211), .A2(n5249), .B1(n4771), .B2(n1150), .ZN(n9507)
         );
  INV_X1 U2032 ( .A(n9507), .ZN(n1284) );
  OR2_X1 U2033 ( .A1(n3934), .A2(n1284), .ZN(n5524) );
  NAND3_X1 U2034 ( .A1(n1291), .A2(n5527), .A3(n5524), .ZN(n1212) );
  NOR2_X1 U2035 ( .A1(n1300), .A2(n1212), .ZN(n1213) );
  OAI211_X1 U2036 ( .C1(n1214), .C2(n1238), .A(n1303), .B(n1213), .ZN(n1307)
         );
  INV_X1 U2037 ( .A(pmp_addr_i[101]), .ZN(n4776) );
  AND2_X1 U2038 ( .A1(pmp_addr_i[131]), .A2(pmp_addr_i[132]), .ZN(n1217) );
  OAI21_X1 U2039 ( .B1(n11897), .B2(n1215), .A(pmp_cfg_i[36]), .ZN(n1227) );
  OAI21_X1 U2040 ( .B1(n1217), .B2(n1216), .A(n1227), .ZN(n1221) );
  NAND2_X1 U2041 ( .A1(n1221), .A2(pmp_addr_i[133]), .ZN(n1218) );
  OAI21_X1 U2042 ( .B1(n1150), .B2(n4776), .A(n1218), .ZN(n9488) );
  INV_X1 U2043 ( .A(n9488), .ZN(n9636) );
  NOR2_X1 U2044 ( .A1(n4605), .A2(n9636), .ZN(n5518) );
  INV_X1 U2045 ( .A(pmp_addr_i[102]), .ZN(n4780) );
  NAND2_X1 U2046 ( .A1(n1219), .A2(pmp_addr_i[134]), .ZN(n1220) );
  OAI21_X1 U2047 ( .B1(n1150), .B2(n4780), .A(n1220), .ZN(n9487) );
  INV_X1 U2048 ( .A(n9487), .ZN(n9606) );
  NOR2_X1 U2049 ( .A1(n5342), .A2(n9606), .ZN(n5520) );
  NOR2_X1 U2050 ( .A1(n5518), .A2(n5520), .ZN(n1241) );
  INV_X1 U2051 ( .A(pmp_addr_i[100]), .ZN(n4763) );
  NAND2_X1 U2052 ( .A1(n1221), .A2(pmp_addr_i[132]), .ZN(n1222) );
  OAI21_X1 U2053 ( .B1(n1150), .B2(n4763), .A(n1222), .ZN(n9479) );
  INV_X1 U2054 ( .A(n9479), .ZN(n9642) );
  NOR2_X1 U2055 ( .A1(instr_addr_o_6_), .A2(n9642), .ZN(n1235) );
  INV_X1 U2056 ( .A(pmp_addr_i[99]), .ZN(n4762) );
  OAI22_X1 U2057 ( .A1(n1227), .A2(n1223), .B1(n4762), .B2(n1150), .ZN(n9478)
         );
  INV_X1 U2058 ( .A(n9478), .ZN(n9647) );
  NOR2_X1 U2059 ( .A1(n4596), .A2(n9647), .ZN(n1224) );
  OR2_X1 U2060 ( .A1(n1235), .A2(n1224), .ZN(n5557) );
  NAND2_X1 U2061 ( .A1(n9584), .A2(pmp_addr_i[98]), .ZN(n1225) );
  OAI21_X1 U2062 ( .B1(n1227), .B2(n1226), .A(n1225), .ZN(n9475) );
  INV_X1 U2063 ( .A(pmp_addr_i[96]), .ZN(n1229) );
  INV_X1 U2064 ( .A(pmp_addr_i[128]), .ZN(n1228) );
  OAI22_X1 U2065 ( .A1(n1229), .A2(n1150), .B1(n9638), .B2(n1228), .ZN(n9637)
         );
  INV_X1 U2066 ( .A(pmp_addr_i[97]), .ZN(n1232) );
  NAND2_X1 U2067 ( .A1(pmp_cfg_i[35]), .A2(pmp_addr_i[128]), .ZN(n1230) );
  NAND3_X1 U2068 ( .A1(n1230), .A2(pmp_cfg_i[36]), .A3(pmp_addr_i[129]), .ZN(
        n1231) );
  OAI21_X1 U2069 ( .B1(n1150), .B2(n1232), .A(n1231), .ZN(n9643) );
  OR2_X1 U2070 ( .A1(n9637), .A2(n9643), .ZN(n1233) );
  NAND2_X1 U2071 ( .A1(n9475), .A2(n1233), .ZN(n1234) );
  INV_X1 U2072 ( .A(n9475), .ZN(n9639) );
  INV_X1 U2073 ( .A(n1233), .ZN(n5547) );
  AOI22_X1 U2074 ( .A1(n3836), .A2(n1234), .B1(n9639), .B2(n5547), .ZN(n1237)
         );
  NAND2_X1 U2075 ( .A1(instr_addr_o_6_), .A2(n9642), .ZN(n5601) );
  NAND2_X1 U2076 ( .A1(n5293), .A2(n9647), .ZN(n5613) );
  OR2_X1 U2077 ( .A1(n5613), .A2(n1235), .ZN(n1236) );
  OAI211_X1 U2078 ( .C1(n5557), .C2(n1237), .A(n5601), .B(n1236), .ZN(n1240)
         );
  NAND2_X1 U2079 ( .A1(n5268), .A2(n9636), .ZN(n5600) );
  NAND2_X1 U2080 ( .A1(n205), .A2(n9606), .ZN(n5605) );
  OAI21_X1 U2081 ( .B1(n5520), .B2(n5600), .A(n5605), .ZN(n1239) );
  OR2_X1 U2082 ( .A1(n1280), .A2(n1242), .ZN(n1265) );
  INV_X1 U2083 ( .A(n1243), .ZN(n1251) );
  NAND2_X1 U2084 ( .A1(n3793), .A2(n1244), .ZN(n1245) );
  OAI22_X1 U2085 ( .A1(n1246), .A2(n1245), .B1(n4631), .B2(n9588), .ZN(n1250)
         );
  NAND2_X1 U2086 ( .A1(n3152), .A2(n9528), .ZN(n1247) );
  OAI22_X1 U2087 ( .A1(n1248), .A2(n1247), .B1(n5192), .B2(n9624), .ZN(n1249)
         );
  AOI21_X1 U2088 ( .B1(n1251), .B2(n1250), .A(n1249), .ZN(n1264) );
  INV_X1 U2089 ( .A(n1252), .ZN(n1255) );
  INV_X1 U2090 ( .A(n9586), .ZN(n1253) );
  NAND2_X1 U2091 ( .A1(n12195), .A2(n1253), .ZN(n1254) );
  OAI22_X1 U2092 ( .A1(n1255), .A2(n1254), .B1(n4438), .B2(n9619), .ZN(n1260)
         );
  NAND2_X1 U2093 ( .A1(n4900), .A2(n1256), .ZN(n1257) );
  OAI22_X1 U2094 ( .A1(n1258), .A2(n1257), .B1(n5115), .B2(n9597), .ZN(n1259)
         );
  INV_X1 U2095 ( .A(n1261), .ZN(n1262) );
  OAI22_X1 U2096 ( .A1(n1265), .A2(n1264), .B1(n1263), .B2(n1262), .ZN(n1283)
         );
  INV_X1 U2097 ( .A(n1267), .ZN(n1271) );
  NAND2_X1 U2098 ( .A1(n5208), .A2(n1268), .ZN(n1270) );
  OAI22_X1 U2099 ( .A1(n1271), .A2(n1270), .B1(n1269), .B2(n9587), .ZN(n1277)
         );
  NAND2_X1 U2100 ( .A1(n5202), .A2(n1272), .ZN(n1274) );
  OAI22_X1 U2101 ( .A1(n1275), .A2(n1274), .B1(n1273), .B2(n9589), .ZN(n1276)
         );
  AOI21_X1 U2102 ( .B1(n1266), .B2(n1277), .A(n1276), .ZN(n1281) );
  INV_X1 U2103 ( .A(n9635), .ZN(n1278) );
  NAND3_X1 U2104 ( .A1(n147), .A2(n1278), .A3(n4444), .ZN(n1279) );
  OAI21_X1 U2105 ( .B1(n1281), .B2(n1280), .A(n1279), .ZN(n1282) );
  NOR2_X1 U2106 ( .A1(n1283), .A2(n1282), .ZN(n1305) );
  INV_X1 U2107 ( .A(n5527), .ZN(n1286) );
  NAND2_X1 U2108 ( .A1(instr_addr_o_12_), .A2(n1285), .ZN(n5616) );
  OAI21_X1 U2109 ( .B1(n1286), .B2(n5607), .A(n5616), .ZN(n1290) );
  NAND2_X1 U2110 ( .A1(n5997), .A2(n1287), .ZN(n5602) );
  NAND2_X1 U2111 ( .A1(n206), .A2(n1288), .ZN(n5606) );
  OAI21_X1 U2112 ( .B1(n5519), .B2(n5602), .A(n5606), .ZN(n1289) );
  NAND2_X1 U2113 ( .A1(n208), .A2(n1292), .ZN(n5612) );
  NAND2_X1 U2114 ( .A1(n5226), .A2(n1293), .ZN(n5604) );
  OAI21_X1 U2115 ( .B1(n5525), .B2(n5612), .A(n5604), .ZN(n1297) );
  NAND2_X1 U2116 ( .A1(n5974), .A2(n1294), .ZN(n5615) );
  OAI22_X1 U2117 ( .A1(n1295), .A2(n5615), .B1(n1922), .B2(n9596), .ZN(n1296)
         );
  AOI21_X1 U2118 ( .B1(n1298), .B2(n1297), .A(n1296), .ZN(n1299) );
  OAI21_X1 U2119 ( .B1(n1301), .B2(n1300), .A(n1299), .ZN(n1302) );
  INV_X1 U2120 ( .A(pmp_addr_i[132]), .ZN(n1308) );
  NAND2_X1 U2121 ( .A1(instr_addr_o_6_), .A2(n1308), .ZN(n1313) );
  NOR2_X1 U2122 ( .A1(n4596), .A2(n1223), .ZN(n1309) );
  AOI22_X1 U2123 ( .A1(n1313), .A2(n1309), .B1(n2611), .B2(pmp_addr_i[132]), 
        .ZN(n1316) );
  NOR2_X1 U2124 ( .A1(pmp_addr_i[129]), .A2(pmp_addr_i[128]), .ZN(n1310) );
  AND2_X1 U2125 ( .A1(n1310), .A2(n1226), .ZN(n1311) );
  OAI22_X1 U2126 ( .A1(n3836), .A2(n1311), .B1(n1310), .B2(n1226), .ZN(n1312)
         );
  OAI211_X1 U2127 ( .C1(pmp_addr_i[131]), .C2(n3839), .A(n1313), .B(n1312), 
        .ZN(n1315) );
  NAND2_X1 U2128 ( .A1(instr_addr_o_8_), .A2(n1148), .ZN(n1318) );
  OAI21_X1 U2129 ( .B1(n4200), .B2(pmp_addr_i[133]), .A(n1318), .ZN(n1314) );
  NAND3_X1 U2132 ( .A1(n1318), .A2(n2424), .A3(pmp_addr_i[133]), .ZN(n1321) );
  NAND2_X1 U2133 ( .A1(n4606), .A2(pmp_addr_i[134]), .ZN(n1320) );
  NAND2_X1 U2134 ( .A1(n3846), .A2(pmp_addr_i[135]), .ZN(n1319) );
  INV_X1 U2135 ( .A(pmp_addr_i[135]), .ZN(n1322) );
  INV_X1 U2136 ( .A(pmp_addr_i[140]), .ZN(n1323) );
  NAND2_X1 U2137 ( .A1(n4788), .A2(n1323), .ZN(n1333) );
  NAND2_X1 U2138 ( .A1(n4061), .A2(n5569), .ZN(n1324) );
  NAND2_X1 U2139 ( .A1(n1333), .A2(n1324), .ZN(n1335) );
  INV_X1 U2140 ( .A(pmp_addr_i[138]), .ZN(n1325) );
  NAND2_X1 U2141 ( .A1(n5250), .A2(n1325), .ZN(n1331) );
  OAI21_X1 U2142 ( .B1(n5052), .B2(pmp_addr_i[137]), .A(n1331), .ZN(n1326) );
  NAND2_X1 U2143 ( .A1(n3100), .A2(n5225), .ZN(n1344) );
  OAI21_X1 U2144 ( .B1(n4578), .B2(pmp_addr_i[141]), .A(n1344), .ZN(n1328) );
  INV_X1 U2145 ( .A(pmp_addr_i[144]), .ZN(n1327) );
  NAND2_X1 U2146 ( .A1(n5047), .A2(n1327), .ZN(n1341) );
  OAI21_X1 U2147 ( .B1(n5048), .B2(pmp_addr_i[143]), .A(n1341), .ZN(n1345) );
  NOR2_X1 U2148 ( .A1(n1328), .A2(n1345), .ZN(n1337) );
  INV_X1 U2149 ( .A(n1431), .ZN(n4493) );
  NOR2_X1 U2150 ( .A1(n4493), .A2(n5249), .ZN(n1330) );
  AOI22_X1 U2151 ( .A1(n1331), .A2(n1330), .B1(n5070), .B2(pmp_addr_i[138]), 
        .ZN(n1336) );
  NOR2_X1 U2152 ( .A1(n5997), .A2(n5569), .ZN(n1332) );
  AOI22_X1 U2153 ( .A1(n1333), .A2(n1332), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[140]), .ZN(n1334) );
  OAI21_X1 U2154 ( .B1(n1336), .B2(n1335), .A(n1334), .ZN(n1338) );
  INV_X1 U2155 ( .A(pmp_addr_i[143]), .ZN(n1339) );
  NOR2_X1 U2156 ( .A1(n4069), .A2(n1339), .ZN(n1340) );
  AOI22_X1 U2157 ( .A1(n1341), .A2(n1340), .B1(n2750), .B2(pmp_addr_i[144]), 
        .ZN(n1348) );
  INV_X1 U2158 ( .A(pmp_addr_i[141]), .ZN(n1342) );
  NOR2_X1 U2159 ( .A1(n208), .A2(n1342), .ZN(n1343) );
  AOI22_X1 U2160 ( .A1(n1344), .A2(n1343), .B1(n5058), .B2(pmp_addr_i[142]), 
        .ZN(n1346) );
  INV_X1 U2161 ( .A(pmp_addr_i[156]), .ZN(n1349) );
  NAND2_X1 U2162 ( .A1(n12161), .A2(n1349), .ZN(n1393) );
  OAI21_X1 U2163 ( .B1(n4656), .B2(pmp_addr_i[155]), .A(n1393), .ZN(n1395) );
  INV_X1 U2164 ( .A(pmp_addr_i[154]), .ZN(n1350) );
  INV_X1 U2165 ( .A(pmp_addr_i[157]), .ZN(n1373) );
  NAND2_X1 U2166 ( .A1(n6018), .A2(n1373), .ZN(n1398) );
  INV_X1 U2167 ( .A(pmp_addr_i[152]), .ZN(n1351) );
  NAND2_X1 U2168 ( .A1(n12158), .A2(n1351), .ZN(n1369) );
  INV_X1 U2169 ( .A(pmp_addr_i[151]), .ZN(n1367) );
  NAND2_X1 U2170 ( .A1(n5202), .A2(n1367), .ZN(n1352) );
  NAND2_X1 U2171 ( .A1(n1369), .A2(n1352), .ZN(n1372) );
  INV_X1 U2172 ( .A(pmp_addr_i[150]), .ZN(n1353) );
  NAND2_X1 U2173 ( .A1(n4835), .A2(n1353), .ZN(n1366) );
  OAI21_X1 U2174 ( .B1(n5086), .B2(pmp_addr_i[149]), .A(n1366), .ZN(n1354) );
  NOR2_X1 U2175 ( .A1(n1372), .A2(n1354), .ZN(n1376) );
  INV_X1 U2176 ( .A(pmp_addr_i[148]), .ZN(n1355) );
  NAND2_X1 U2177 ( .A1(n12157), .A2(n1355), .ZN(n1384) );
  INV_X1 U2178 ( .A(pmp_addr_i[147]), .ZN(n1383) );
  NAND2_X1 U2179 ( .A1(n3152), .A2(n1383), .ZN(n1356) );
  NAND2_X1 U2180 ( .A1(n1384), .A2(n1356), .ZN(n1387) );
  INV_X1 U2181 ( .A(pmp_addr_i[146]), .ZN(n1357) );
  NAND2_X1 U2182 ( .A1(n6027), .A2(n1357), .ZN(n1381) );
  INV_X1 U2183 ( .A(pmp_addr_i[145]), .ZN(n1380) );
  NAND2_X1 U2184 ( .A1(n3793), .A2(n1380), .ZN(n1358) );
  NAND2_X1 U2185 ( .A1(n1381), .A2(n1358), .ZN(n1359) );
  NOR2_X1 U2186 ( .A1(n1387), .A2(n1359), .ZN(n1360) );
  INV_X1 U2187 ( .A(pmp_addr_i[149]), .ZN(n1364) );
  NOR2_X1 U2188 ( .A1(n5208), .A2(n1364), .ZN(n1365) );
  AOI22_X1 U2189 ( .A1(n1366), .A2(n1365), .B1(n1269), .B2(pmp_addr_i[150]), 
        .ZN(n1371) );
  NOR2_X1 U2190 ( .A1(n5365), .A2(n1367), .ZN(n1368) );
  AOI22_X1 U2191 ( .A1(n1369), .A2(n1368), .B1(n3806), .B2(pmp_addr_i[152]), 
        .ZN(n1370) );
  OAI21_X1 U2192 ( .B1(n1372), .B2(n1371), .A(n1370), .ZN(n1375) );
  NOR2_X1 U2193 ( .A1(pmp_addr_i[159]), .A2(pmp_addr_i[158]), .ZN(n9451) );
  OAI21_X1 U2194 ( .B1(n6018), .B2(n1373), .A(n9451), .ZN(n1374) );
  AOI21_X1 U2195 ( .B1(n1377), .B2(n1375), .A(n1374), .ZN(n1402) );
  INV_X1 U2196 ( .A(n1376), .ZN(n1379) );
  NOR2_X1 U2197 ( .A1(n1379), .A2(n1378), .ZN(n1400) );
  NOR2_X1 U2198 ( .A1(n5100), .A2(n1380), .ZN(n1382) );
  AOI22_X1 U2199 ( .A1(n1382), .A2(n1381), .B1(n2569), .B2(pmp_addr_i[146]), 
        .ZN(n1388) );
  NOR2_X1 U2200 ( .A1(instr_addr_o_21_), .A2(n1383), .ZN(n1385) );
  AOI22_X1 U2201 ( .A1(n1385), .A2(n1384), .B1(n999), .B2(pmp_addr_i[148]), 
        .ZN(n1386) );
  OAI21_X1 U2202 ( .B1(n1388), .B2(n1387), .A(n1386), .ZN(n1399) );
  INV_X1 U2203 ( .A(pmp_addr_i[153]), .ZN(n1389) );
  NOR2_X1 U2204 ( .A1(n5162), .A2(n1389), .ZN(n1390) );
  AOI22_X1 U2205 ( .A1(n1391), .A2(n1390), .B1(n5111), .B2(pmp_addr_i[154]), 
        .ZN(n1396) );
  NOR2_X1 U2206 ( .A1(instr_addr_o_29_), .A2(n5148), .ZN(n1392) );
  AOI22_X1 U2207 ( .A1(n1393), .A2(n1392), .B1(n5115), .B2(pmp_addr_i[156]), 
        .ZN(n1394) );
  OAI21_X1 U2208 ( .B1(n1396), .B2(n1395), .A(n1394), .ZN(n1397) );
  AOI22_X1 U2209 ( .A1(n1400), .A2(n1399), .B1(n1398), .B2(n1397), .ZN(n1401)
         );
  INV_X1 U2210 ( .A(pmp_cfg_i[99]), .ZN(n1452) );
  OR2_X1 U2211 ( .A1(n1452), .A2(pmp_cfg_i[100]), .ZN(n3475) );
  NAND2_X1 U2212 ( .A1(pmp_addr_i[384]), .A2(pmp_addr_i[385]), .ZN(n3474) );
  INV_X1 U2213 ( .A(pmp_addr_i[386]), .ZN(n3526) );
  OR2_X1 U2214 ( .A1(n3474), .A2(n3526), .ZN(n3461) );
  INV_X1 U2215 ( .A(pmp_addr_i[387]), .ZN(n3513) );
  NOR2_X1 U2216 ( .A1(n3461), .A2(n3513), .ZN(n11420) );
  NAND2_X1 U2217 ( .A1(n11420), .A2(pmp_cfg_i[99]), .ZN(n1441) );
  AND2_X1 U2218 ( .A1(pmp_addr_i[388]), .A2(pmp_addr_i[389]), .ZN(n1442) );
  AND2_X1 U2219 ( .A1(pmp_addr_i[390]), .A2(pmp_addr_i[391]), .ZN(n1414) );
  NAND2_X1 U2220 ( .A1(n1442), .A2(n1414), .ZN(n1408) );
  OR2_X1 U2221 ( .A1(n1441), .A2(n1408), .ZN(n1433) );
  NAND3_X1 U2222 ( .A1(n1433), .A2(pmp_addr_i[392]), .A3(pmp_cfg_i[100]), .ZN(
        n1409) );
  OAI21_X1 U2223 ( .B1(n3475), .B2(n3127), .A(n1409), .ZN(n8544) );
  INV_X1 U2224 ( .A(n8544), .ZN(n8670) );
  OR2_X1 U2225 ( .A1(n5262), .A2(n8670), .ZN(n1411) );
  INV_X1 U2226 ( .A(n1411), .ZN(n3450) );
  INV_X1 U2227 ( .A(pmp_addr_i[359]), .ZN(n2959) );
  NAND3_X1 U2228 ( .A1(n1433), .A2(pmp_addr_i[391]), .A3(pmp_cfg_i[100]), .ZN(
        n1410) );
  OAI21_X1 U2229 ( .B1(n3475), .B2(n2959), .A(n1410), .ZN(n8543) );
  INV_X1 U2230 ( .A(n8543), .ZN(n8673) );
  NOR2_X1 U2231 ( .A1(n4204), .A2(n8673), .ZN(n3411) );
  AND2_X1 U2232 ( .A1(n153), .A2(n8673), .ZN(n3419) );
  AOI22_X1 U2233 ( .A1(n3419), .A2(n1411), .B1(n12202), .B2(n8670), .ZN(n1440)
         );
  OAI21_X1 U2234 ( .B1(n3450), .B2(n3411), .A(n1440), .ZN(n1439) );
  NAND2_X1 U2235 ( .A1(pmp_addr_i[392]), .A2(pmp_addr_i[393]), .ZN(n1432) );
  NAND2_X1 U2236 ( .A1(pmp_addr_i[395]), .A2(pmp_addr_i[394]), .ZN(n1412) );
  OR2_X1 U2237 ( .A1(n1432), .A2(n1412), .ZN(n3463) );
  NAND2_X1 U2238 ( .A1(pmp_addr_i[396]), .A2(pmp_addr_i[397]), .ZN(n1413) );
  NOR2_X1 U2239 ( .A1(n3463), .A2(n1413), .ZN(n1419) );
  AND4_X1 U2240 ( .A1(n1442), .A2(n1414), .A3(pmp_addr_i[399]), .A4(
        pmp_addr_i[398]), .ZN(n1415) );
  INV_X1 U2241 ( .A(pmp_addr_i[400]), .ZN(n3589) );
  NAND2_X1 U2242 ( .A1(n1644), .A2(pmp_addr_i[368]), .ZN(n1416) );
  OAI21_X1 U2243 ( .B1(n3476), .B2(n3589), .A(n1416), .ZN(n8652) );
  INV_X1 U2244 ( .A(n8652), .ZN(n1417) );
  NOR2_X1 U2245 ( .A1(n6019), .A2(n1417), .ZN(n1472) );
  INV_X1 U2246 ( .A(pmp_addr_i[399]), .ZN(n3541) );
  NAND2_X1 U2247 ( .A1(n1644), .A2(pmp_addr_i[367]), .ZN(n1418) );
  OAI21_X1 U2248 ( .B1(n3476), .B2(n3541), .A(n1418), .ZN(n8514) );
  INV_X1 U2249 ( .A(n8514), .ZN(n8691) );
  NOR2_X1 U2250 ( .A1(n5974), .A2(n8691), .ZN(n3451) );
  OR2_X1 U2251 ( .A1(n1472), .A2(n3451), .ZN(n1470) );
  INV_X1 U2252 ( .A(n1419), .ZN(n1420) );
  OAI21_X1 U2253 ( .B1(n1433), .B2(n1420), .A(pmp_cfg_i[100]), .ZN(n1424) );
  INV_X1 U2254 ( .A(pmp_addr_i[397]), .ZN(n3455) );
  NAND2_X1 U2255 ( .A1(n1644), .A2(pmp_addr_i[365]), .ZN(n1421) );
  OAI21_X1 U2256 ( .B1(n1424), .B2(n3455), .A(n1421), .ZN(n8512) );
  INV_X1 U2257 ( .A(n8512), .ZN(n8678) );
  NOR2_X1 U2258 ( .A1(n208), .A2(n8678), .ZN(n3410) );
  INV_X1 U2259 ( .A(pmp_addr_i[398]), .ZN(n1423) );
  NAND2_X1 U2260 ( .A1(n1644), .A2(pmp_addr_i[366]), .ZN(n1422) );
  OAI21_X1 U2261 ( .B1(n1424), .B2(n1423), .A(n1422), .ZN(n8690) );
  INV_X1 U2262 ( .A(n8690), .ZN(n11409) );
  NOR2_X1 U2263 ( .A1(n3100), .A2(n11409), .ZN(n3426) );
  OR2_X1 U2264 ( .A1(n3410), .A2(n3426), .ZN(n1425) );
  NOR2_X1 U2265 ( .A1(n1470), .A2(n1425), .ZN(n1469) );
  OAI21_X1 U2266 ( .B1(n1433), .B2(n3463), .A(pmp_cfg_i[100]), .ZN(n1430) );
  INV_X1 U2267 ( .A(pmp_addr_i[395]), .ZN(n1427) );
  NAND2_X1 U2268 ( .A1(n1644), .A2(pmp_addr_i[363]), .ZN(n1426) );
  OAI21_X1 U2269 ( .B1(n1430), .B2(n1427), .A(n1426), .ZN(n8692) );
  INV_X1 U2270 ( .A(n8692), .ZN(n8676) );
  NOR2_X1 U2271 ( .A1(n149), .A2(n8676), .ZN(n3412) );
  INV_X1 U2272 ( .A(pmp_addr_i[396]), .ZN(n1429) );
  NAND2_X1 U2273 ( .A1(n1644), .A2(pmp_addr_i[364]), .ZN(n1428) );
  OAI21_X1 U2274 ( .B1(n1430), .B2(n1429), .A(n1428), .ZN(n8520) );
  INV_X1 U2275 ( .A(n8520), .ZN(n8679) );
  NOR2_X1 U2276 ( .A1(n206), .A2(n8679), .ZN(n3438) );
  NOR2_X1 U2277 ( .A1(n3412), .A2(n3438), .ZN(n1468) );
  OAI21_X1 U2278 ( .B1(n1433), .B2(n1432), .A(pmp_cfg_i[100]), .ZN(n1437) );
  INV_X1 U2279 ( .A(pmp_addr_i[393]), .ZN(n3420) );
  NAND2_X1 U2280 ( .A1(n1644), .A2(pmp_addr_i[361]), .ZN(n1434) );
  OAI21_X1 U2281 ( .B1(n1437), .B2(n3420), .A(n1434), .ZN(n8517) );
  INV_X1 U2282 ( .A(n8517), .ZN(n8671) );
  INV_X1 U2283 ( .A(pmp_addr_i[394]), .ZN(n1436) );
  NAND2_X1 U2284 ( .A1(n1644), .A2(pmp_addr_i[362]), .ZN(n1435) );
  OAI21_X1 U2285 ( .B1(n1437), .B2(n1436), .A(n1435), .ZN(n8518) );
  INV_X1 U2286 ( .A(n8518), .ZN(n8677) );
  NOR2_X1 U2287 ( .A1(instr_addr_o_12_), .A2(n8677), .ZN(n3427) );
  NOR2_X1 U2288 ( .A1(n3442), .A2(n3427), .ZN(n1438) );
  INV_X1 U2289 ( .A(n1440), .ZN(n1448) );
  NAND2_X1 U2290 ( .A1(n1441), .A2(pmp_cfg_i[100]), .ZN(n1451) );
  OAI21_X1 U2291 ( .B1(n1442), .B2(n220), .A(n1451), .ZN(n1444) );
  NAND2_X1 U2292 ( .A1(n1444), .A2(pmp_addr_i[390]), .ZN(n1443) );
  OAI21_X1 U2293 ( .B1(n3475), .B2(n3123), .A(n1443), .ZN(n8540) );
  INV_X1 U2294 ( .A(n8540), .ZN(n8672) );
  OR2_X1 U2295 ( .A1(n5342), .A2(n8672), .ZN(n3439) );
  INV_X1 U2296 ( .A(n3439), .ZN(n1446) );
  NAND2_X1 U2297 ( .A1(n1444), .A2(pmp_addr_i[389]), .ZN(n1445) );
  OAI21_X1 U2298 ( .B1(n3475), .B2(n3129), .A(n1445), .ZN(n8541) );
  INV_X1 U2299 ( .A(n8541), .ZN(n8665) );
  NAND2_X1 U2300 ( .A1(n5268), .A2(n8665), .ZN(n3445) );
  NAND2_X1 U2301 ( .A1(n205), .A2(n8672), .ZN(n3431) );
  OAI21_X1 U2302 ( .B1(n1446), .B2(n3445), .A(n3431), .ZN(n1447) );
  NOR2_X1 U2303 ( .A1(n1448), .A2(n1447), .ZN(n1463) );
  INV_X1 U2304 ( .A(pmp_addr_i[388]), .ZN(n3553) );
  NAND2_X1 U2305 ( .A1(n1644), .A2(pmp_addr_i[356]), .ZN(n1449) );
  OAI21_X1 U2306 ( .B1(n1451), .B2(n3553), .A(n1449), .ZN(n8533) );
  INV_X1 U2307 ( .A(n8533), .ZN(n8524) );
  NOR2_X1 U2308 ( .A1(n12152), .A2(n8524), .ZN(n3409) );
  NAND2_X1 U2309 ( .A1(n1644), .A2(pmp_addr_i[355]), .ZN(n1450) );
  OAI21_X1 U2310 ( .B1(n1451), .B2(n3513), .A(n1450), .ZN(n8534) );
  INV_X1 U2311 ( .A(n8534), .ZN(n8694) );
  NOR2_X1 U2312 ( .A1(n4596), .A2(n8694), .ZN(n3467) );
  OAI21_X1 U2313 ( .B1(n3474), .B2(n1452), .A(pmp_cfg_i[100]), .ZN(n1456) );
  INV_X1 U2314 ( .A(pmp_addr_i[385]), .ZN(n1453) );
  INV_X1 U2315 ( .A(pmp_addr_i[353]), .ZN(n5950) );
  OAI22_X1 U2316 ( .A1(n1456), .A2(n1453), .B1(n3475), .B2(n5950), .ZN(n8660)
         );
  INV_X1 U2317 ( .A(pmp_addr_i[352]), .ZN(n5949) );
  NAND2_X1 U2318 ( .A1(n1454), .A2(pmp_addr_i[384]), .ZN(n1455) );
  OAI21_X1 U2319 ( .B1(n3475), .B2(n5949), .A(n1455), .ZN(n8696) );
  OR2_X1 U2320 ( .A1(n8660), .A2(n8696), .ZN(n1457) );
  INV_X1 U2321 ( .A(pmp_addr_i[354]), .ZN(n2937) );
  OAI22_X1 U2322 ( .A1(n1456), .A2(n3526), .B1(n3475), .B2(n2937), .ZN(n8530)
         );
  NAND2_X1 U2323 ( .A1(n1457), .A2(n8530), .ZN(n1458) );
  INV_X1 U2324 ( .A(n8530), .ZN(n8661) );
  INV_X1 U2325 ( .A(n1457), .ZN(n3477) );
  AOI22_X1 U2326 ( .A1(n3836), .A2(n1458), .B1(n8661), .B2(n3477), .ZN(n1459)
         );
  NOR3_X1 U2327 ( .A1(n3409), .A2(n3467), .A3(n1459), .ZN(n1461) );
  NAND2_X1 U2328 ( .A1(n5293), .A2(n8694), .ZN(n3466) );
  NAND2_X1 U2329 ( .A1(instr_addr_o_6_), .A2(n8524), .ZN(n3418) );
  OAI21_X1 U2330 ( .B1(n3409), .B2(n3466), .A(n3418), .ZN(n1460) );
  OR2_X1 U2331 ( .A1(n12267), .A2(n8665), .ZN(n3444) );
  OAI211_X1 U2332 ( .C1(n1461), .C2(n1460), .A(n3439), .B(n3444), .ZN(n1462)
         );
  AND2_X1 U2333 ( .A1(n1463), .A2(n1462), .ZN(n1464) );
  NOR2_X1 U2334 ( .A1(n1465), .A2(n1464), .ZN(n1507) );
  NAND2_X1 U2335 ( .A1(instr_addr_o_11_), .A2(n8671), .ZN(n3441) );
  NAND2_X1 U2336 ( .A1(n5250), .A2(n8677), .ZN(n3428) );
  OAI21_X1 U2337 ( .B1(n3427), .B2(n3441), .A(n3428), .ZN(n1467) );
  NAND2_X1 U2338 ( .A1(n149), .A2(n8676), .ZN(n3421) );
  OAI22_X1 U2339 ( .A1(n3438), .A2(n3421), .B1(instr_addr_o_14__BAR), .B2(
        n8520), .ZN(n1466) );
  AOI21_X1 U2340 ( .B1(n1468), .B2(n1467), .A(n1466), .ZN(n1478) );
  INV_X1 U2341 ( .A(n1469), .ZN(n1477) );
  INV_X1 U2342 ( .A(n1470), .ZN(n1475) );
  NAND2_X1 U2343 ( .A1(n12179), .A2(n8678), .ZN(n1471) );
  OAI22_X1 U2344 ( .A1(n3426), .A2(n1471), .B1(n5058), .B2(n8690), .ZN(n1474)
         );
  NAND2_X1 U2345 ( .A1(n5974), .A2(n8691), .ZN(n3452) );
  OAI22_X1 U2346 ( .A1(n1472), .A2(n3452), .B1(n2082), .B2(n8652), .ZN(n1473)
         );
  AOI21_X1 U2347 ( .B1(n1475), .B2(n1474), .A(n1473), .ZN(n1476) );
  OAI21_X1 U2348 ( .B1(n1478), .B2(n1477), .A(n1476), .ZN(n1506) );
  INV_X1 U2349 ( .A(pmp_addr_i[408]), .ZN(n3591) );
  NAND2_X1 U2350 ( .A1(n1644), .A2(pmp_addr_i[376]), .ZN(n1479) );
  OAI21_X1 U2351 ( .B1(n3476), .B2(n3591), .A(n1479), .ZN(n8636) );
  INV_X1 U2352 ( .A(n8636), .ZN(n1480) );
  NOR2_X1 U2353 ( .A1(n12158), .A2(n1480), .ZN(n1544) );
  INV_X1 U2354 ( .A(pmp_addr_i[407]), .ZN(n3628) );
  NAND2_X1 U2355 ( .A1(n1644), .A2(pmp_addr_i[375]), .ZN(n1481) );
  OAI21_X1 U2356 ( .B1(n3476), .B2(n3628), .A(n1481), .ZN(n8653) );
  INV_X1 U2357 ( .A(n8653), .ZN(n1542) );
  INV_X1 U2359 ( .A(pmp_addr_i[405]), .ZN(n3601) );
  NAND2_X1 U2360 ( .A1(n1644), .A2(pmp_addr_i[373]), .ZN(n1483) );
  OAI21_X1 U2361 ( .B1(n3476), .B2(n3601), .A(n1483), .ZN(n8643) );
  INV_X1 U2362 ( .A(n8643), .ZN(n1539) );
  INV_X1 U2363 ( .A(pmp_addr_i[406]), .ZN(n3605) );
  NAND2_X1 U2364 ( .A1(n1644), .A2(pmp_addr_i[374]), .ZN(n1484) );
  OAI21_X1 U2365 ( .B1(n3476), .B2(n3605), .A(n1484), .ZN(n8635) );
  INV_X1 U2366 ( .A(n8635), .ZN(n1485) );
  OR2_X1 U2367 ( .A1(n5330), .A2(n1485), .ZN(n1538) );
  OAI21_X1 U2368 ( .B1(n5208), .B2(n1539), .A(n1538), .ZN(n1486) );
  INV_X1 U2369 ( .A(pmp_addr_i[403]), .ZN(n3581) );
  NAND2_X1 U2370 ( .A1(n1644), .A2(pmp_addr_i[371]), .ZN(n1487) );
  OAI21_X1 U2371 ( .B1(n3476), .B2(n3581), .A(n1487), .ZN(n8642) );
  INV_X1 U2372 ( .A(n8642), .ZN(n1516) );
  INV_X1 U2373 ( .A(pmp_addr_i[404]), .ZN(n3603) );
  NAND2_X1 U2374 ( .A1(n1644), .A2(pmp_addr_i[372]), .ZN(n1488) );
  INV_X1 U2375 ( .A(n8634), .ZN(n1489) );
  OR2_X1 U2376 ( .A1(n12157), .A2(n1489), .ZN(n1515) );
  OAI21_X1 U2377 ( .B1(n3152), .B2(n1516), .A(n1515), .ZN(n1510) );
  INV_X1 U2378 ( .A(pmp_addr_i[401]), .ZN(n3583) );
  NAND2_X1 U2379 ( .A1(n1644), .A2(pmp_addr_i[369]), .ZN(n1490) );
  OAI21_X1 U2380 ( .B1(n3476), .B2(n3583), .A(n1490), .ZN(n8633) );
  INV_X1 U2381 ( .A(n8633), .ZN(n1512) );
  INV_X1 U2382 ( .A(pmp_addr_i[402]), .ZN(n3607) );
  NAND2_X1 U2383 ( .A1(n1644), .A2(pmp_addr_i[370]), .ZN(n1491) );
  OAI21_X1 U2384 ( .B1(n3476), .B2(n3607), .A(n1491), .ZN(n8641) );
  INV_X1 U2385 ( .A(n8641), .ZN(n1492) );
  OR2_X1 U2386 ( .A1(n4802), .A2(n1492), .ZN(n1511) );
  OAI21_X1 U2387 ( .B1(n5100), .B2(n1512), .A(n1511), .ZN(n1493) );
  NOR2_X1 U2388 ( .A1(n1510), .A2(n1493), .ZN(n1494) );
  NAND2_X1 U2389 ( .A1(n1508), .A2(n1494), .ZN(n1504) );
  NAND2_X1 U2390 ( .A1(n1644), .A2(pmp_addr_i[380]), .ZN(n1495) );
  OAI21_X1 U2391 ( .B1(n3476), .B2(n1598), .A(n1495), .ZN(n8651) );
  INV_X1 U2392 ( .A(n8651), .ZN(n1496) );
  NOR2_X1 U2393 ( .A1(n4753), .A2(n1496), .ZN(n1528) );
  NAND2_X1 U2394 ( .A1(n1644), .A2(pmp_addr_i[379]), .ZN(n1497) );
  OAI21_X1 U2395 ( .B1(n3476), .B2(n1631), .A(n1497), .ZN(n8659) );
  INV_X1 U2396 ( .A(n8659), .ZN(n1526) );
  NOR2_X1 U2397 ( .A1(n5149), .A2(n1526), .ZN(n1498) );
  NOR2_X1 U2398 ( .A1(n1528), .A2(n1498), .ZN(n1531) );
  INV_X1 U2399 ( .A(pmp_addr_i[381]), .ZN(n1499) );
  INV_X1 U2400 ( .A(pmp_addr_i[413]), .ZN(n12085) );
  OR2_X1 U2401 ( .A1(n3476), .A2(n12085), .ZN(n11459) );
  OAI21_X1 U2402 ( .B1(n1499), .B2(n3475), .A(n11459), .ZN(n8584) );
  NOR2_X1 U2403 ( .A1(pmp_addr_i[382]), .A2(pmp_addr_i[383]), .ZN(n10111) );
  INV_X1 U2404 ( .A(n10111), .ZN(n1548) );
  AOI21_X1 U2405 ( .B1(n4660), .B2(n8584), .A(n1548), .ZN(n1532) );
  INV_X1 U2406 ( .A(pmp_addr_i[410]), .ZN(n3623) );
  NAND2_X1 U2407 ( .A1(n1644), .A2(pmp_addr_i[378]), .ZN(n1500) );
  OAI21_X1 U2408 ( .B1(n3476), .B2(n3623), .A(n1500), .ZN(n8654) );
  INV_X1 U2409 ( .A(n8654), .ZN(n1501) );
  OR2_X1 U2410 ( .A1(n5368), .A2(n1501), .ZN(n1522) );
  INV_X1 U2411 ( .A(pmp_addr_i[409]), .ZN(n3625) );
  NAND2_X1 U2412 ( .A1(n1644), .A2(pmp_addr_i[377]), .ZN(n1502) );
  OAI21_X1 U2413 ( .B1(n3476), .B2(n3625), .A(n1502), .ZN(n8644) );
  NAND2_X1 U2414 ( .A1(n4147), .A2(n8644), .ZN(n1503) );
  NAND4_X1 U2415 ( .A1(n1531), .A2(n1532), .A3(n1522), .A4(n1503), .ZN(n1550)
         );
  NOR2_X1 U2416 ( .A1(n1504), .A2(n1550), .ZN(n1505) );
  OAI21_X1 U2417 ( .B1(n1507), .B2(n1506), .A(n1505), .ZN(n1554) );
  OR2_X1 U2418 ( .A1(n1550), .A2(n1509), .ZN(n1536) );
  INV_X1 U2419 ( .A(n1510), .ZN(n1521) );
  INV_X1 U2420 ( .A(n1511), .ZN(n1514) );
  NAND2_X1 U2421 ( .A1(instr_addr_o_19_), .A2(n1512), .ZN(n1513) );
  OAI22_X1 U2422 ( .A1(n1514), .A2(n1513), .B1(n4631), .B2(n8641), .ZN(n1520)
         );
  INV_X1 U2423 ( .A(n1515), .ZN(n1518) );
  NAND2_X1 U2424 ( .A1(n3152), .A2(n1516), .ZN(n1517) );
  OAI22_X1 U2425 ( .A1(n1518), .A2(n1517), .B1(n999), .B2(n8634), .ZN(n1519)
         );
  AOI21_X1 U2426 ( .B1(n1521), .B2(n1520), .A(n1519), .ZN(n1535) );
  INV_X1 U2427 ( .A(n1522), .ZN(n1525) );
  INV_X1 U2428 ( .A(n8644), .ZN(n1523) );
  NAND2_X1 U2429 ( .A1(n12195), .A2(n1523), .ZN(n1524) );
  OAI22_X1 U2430 ( .A1(n1525), .A2(n1524), .B1(n5111), .B2(n8654), .ZN(n1530)
         );
  NAND2_X1 U2431 ( .A1(n5550), .A2(n1526), .ZN(n1527) );
  OAI22_X1 U2432 ( .A1(n1528), .A2(n1527), .B1(n5115), .B2(n8651), .ZN(n1529)
         );
  AOI21_X1 U2433 ( .B1(n1531), .B2(n1530), .A(n1529), .ZN(n1534) );
  INV_X1 U2434 ( .A(n1532), .ZN(n1533) );
  INV_X1 U2436 ( .A(n1537), .ZN(n1547) );
  INV_X1 U2437 ( .A(n1538), .ZN(n1541) );
  NAND2_X1 U2438 ( .A1(n5208), .A2(n1539), .ZN(n1540) );
  OAI22_X1 U2439 ( .A1(n1541), .A2(n1540), .B1(n1269), .B2(n8635), .ZN(n1546)
         );
  NAND2_X1 U2440 ( .A1(n5202), .A2(n1542), .ZN(n1543) );
  OAI22_X1 U2441 ( .A1(n1544), .A2(n1543), .B1(n3806), .B2(n8636), .ZN(n1545)
         );
  AOI21_X1 U2442 ( .B1(n1547), .B2(n1546), .A(n1545), .ZN(n1551) );
  INV_X1 U2443 ( .A(n8584), .ZN(n8693) );
  NAND3_X1 U2444 ( .A1(instr_addr_o_31_), .A2(n8693), .A3(n10111), .ZN(n1549)
         );
  OAI21_X1 U2445 ( .B1(n1551), .B2(n1550), .A(n1549), .ZN(n1552) );
  NAND2_X1 U2446 ( .A1(n5047), .A2(n3589), .ZN(n1565) );
  OAI21_X1 U2447 ( .B1(n5048), .B2(pmp_addr_i[399]), .A(n1565), .ZN(n1567) );
  NAND2_X1 U2448 ( .A1(n3100), .A2(n1423), .ZN(n1563) );
  OAI21_X1 U2449 ( .B1(n6017), .B2(pmp_addr_i[397]), .A(n1563), .ZN(n1555) );
  NOR2_X1 U2450 ( .A1(n1567), .A2(n1555), .ZN(n1594) );
  NAND2_X1 U2451 ( .A1(n5250), .A2(n1436), .ZN(n1590) );
  NOR2_X1 U2452 ( .A1(n5069), .A2(n3420), .ZN(n1556) );
  AOI22_X1 U2453 ( .A1(n1590), .A2(n1556), .B1(n5070), .B2(pmp_addr_i[394]), 
        .ZN(n1561) );
  NAND2_X1 U2454 ( .A1(n5251), .A2(n1429), .ZN(n1559) );
  NAND2_X1 U2455 ( .A1(n4061), .A2(n1427), .ZN(n1557) );
  NAND2_X1 U2456 ( .A1(n1559), .A2(n1557), .ZN(n1592) );
  NOR2_X1 U2457 ( .A1(n150), .A2(n1427), .ZN(n1558) );
  AOI22_X1 U2458 ( .A1(n1559), .A2(n1558), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[396]), .ZN(n1560) );
  OAI21_X1 U2459 ( .B1(n1561), .B2(n1592), .A(n1560), .ZN(n1570) );
  NOR2_X1 U2460 ( .A1(n12178), .A2(n3455), .ZN(n1562) );
  AOI22_X1 U2461 ( .A1(n1563), .A2(n1562), .B1(n5058), .B2(pmp_addr_i[398]), 
        .ZN(n1568) );
  NOR2_X1 U2462 ( .A1(n4069), .A2(n3541), .ZN(n1564) );
  NAND2_X1 U2464 ( .A1(instr_addr_o_6_), .A2(n3553), .ZN(n1576) );
  NOR2_X1 U2465 ( .A1(n4596), .A2(n3513), .ZN(n1571) );
  AOI22_X1 U2466 ( .A1(n1576), .A2(n1571), .B1(n2611), .B2(pmp_addr_i[388]), 
        .ZN(n1580) );
  OR2_X1 U2467 ( .A1(pmp_addr_i[385]), .A2(pmp_addr_i[384]), .ZN(n1572) );
  NOR2_X1 U2468 ( .A1(n1572), .A2(pmp_addr_i[386]), .ZN(n1574) );
  INV_X1 U2469 ( .A(n1572), .ZN(n1573) );
  OAI22_X1 U2470 ( .A1(n5899), .A2(n1574), .B1(n1573), .B2(n3526), .ZN(n1575)
         );
  OAI211_X1 U2471 ( .C1(pmp_addr_i[387]), .C2(n3839), .A(n1576), .B(n1575), 
        .ZN(n1579) );
  INV_X1 U2472 ( .A(pmp_addr_i[390]), .ZN(n1577) );
  NAND2_X1 U2473 ( .A1(n205), .A2(n1577), .ZN(n1581) );
  OAI21_X1 U2474 ( .B1(n3844), .B2(pmp_addr_i[389]), .A(n1581), .ZN(n1578) );
  AOI21_X1 U2475 ( .B1(n1580), .B2(n1579), .A(n1578), .ZN(n1597) );
  NAND3_X1 U2476 ( .A1(n1581), .A2(n3844), .A3(pmp_addr_i[389]), .ZN(n1585) );
  INV_X1 U2477 ( .A(pmp_addr_i[392]), .ZN(n1586) );
  NOR2_X1 U2478 ( .A1(n5270), .A2(n1586), .ZN(n1588) );
  INV_X1 U2479 ( .A(n1588), .ZN(n1584) );
  NAND2_X1 U2480 ( .A1(n3894), .A2(pmp_addr_i[390]), .ZN(n1583) );
  NAND2_X1 U2481 ( .A1(n3846), .A2(pmp_addr_i[391]), .ZN(n1582) );
  NAND4_X1 U2482 ( .A1(n1585), .A2(n1584), .A3(n1583), .A4(n1582), .ZN(n1596)
         );
  INV_X1 U2483 ( .A(pmp_addr_i[391]), .ZN(n1587) );
  AOI22_X1 U2484 ( .A1(n155), .A2(n1587), .B1(instr_addr_o_10_), .B2(n1586), 
        .ZN(n1589) );
  NOR2_X1 U2485 ( .A1(n1589), .A2(n1588), .ZN(n1593) );
  OAI21_X1 U2486 ( .B1(n5052), .B2(pmp_addr_i[393]), .A(n1590), .ZN(n1591) );
  NOR3_X1 U2487 ( .A1(n1593), .A2(n1592), .A3(n1591), .ZN(n1595) );
  OAI211_X1 U2488 ( .C1(n1597), .C2(n1596), .A(n1595), .B(n1594), .ZN(n1605)
         );
  INV_X1 U2489 ( .A(pmp_addr_i[412]), .ZN(n1598) );
  NAND2_X1 U2490 ( .A1(n12161), .A2(n1598), .ZN(n1634) );
  OAI21_X1 U2491 ( .B1(n4623), .B2(pmp_addr_i[411]), .A(n1634), .ZN(n1636) );
  NAND2_X1 U2492 ( .A1(n5368), .A2(n3623), .ZN(n1630) );
  NAND2_X1 U2493 ( .A1(n4866), .A2(n12085), .ZN(n1638) );
  OAI211_X1 U2494 ( .C1(n5094), .C2(pmp_addr_i[409]), .A(n1630), .B(n1638), 
        .ZN(n1599) );
  NOR2_X1 U2495 ( .A1(n1636), .A2(n1599), .ZN(n1627) );
  NAND2_X1 U2496 ( .A1(n4836), .A2(n3603), .ZN(n1621) );
  NAND2_X1 U2497 ( .A1(n3152), .A2(n3581), .ZN(n1600) );
  AND2_X1 U2498 ( .A1(n1621), .A2(n1600), .ZN(n1618) );
  NAND2_X1 U2499 ( .A1(n12158), .A2(n3591), .ZN(n1610) );
  NAND2_X1 U2500 ( .A1(n5202), .A2(n3628), .ZN(n1601) );
  NAND2_X1 U2501 ( .A1(n1610), .A2(n1601), .ZN(n1613) );
  NAND2_X1 U2502 ( .A1(n5330), .A2(n3605), .ZN(n1608) );
  OAI21_X1 U2503 ( .B1(n5086), .B2(pmp_addr_i[405]), .A(n1608), .ZN(n1602) );
  NOR2_X1 U2504 ( .A1(n1613), .A2(n1602), .ZN(n1626) );
  NAND2_X1 U2505 ( .A1(n6027), .A2(n3607), .ZN(n1619) );
  NAND2_X1 U2506 ( .A1(instr_addr_o_19_), .A2(n3583), .ZN(n1603) );
  AND2_X1 U2507 ( .A1(n1619), .A2(n1603), .ZN(n1604) );
  NOR2_X1 U2508 ( .A1(instr_addr_o_23_), .A2(n3601), .ZN(n1607) );
  AOI22_X1 U2509 ( .A1(n1608), .A2(n1607), .B1(n2580), .B2(pmp_addr_i[406]), 
        .ZN(n1612) );
  NOR2_X1 U2510 ( .A1(n5365), .A2(n3628), .ZN(n1609) );
  AOI22_X1 U2511 ( .A1(n1610), .A2(n1609), .B1(n1273), .B2(pmp_addr_i[408]), 
        .ZN(n1611) );
  OAI21_X1 U2512 ( .B1(n1613), .B2(n1612), .A(n1611), .ZN(n1614) );
  NAND2_X1 U2513 ( .A1(n1627), .A2(n1614), .ZN(n1617) );
  NOR2_X1 U2514 ( .A1(pmp_addr_i[415]), .A2(pmp_addr_i[414]), .ZN(n1616) );
  BUF_X1 U2515 ( .A(n3295), .Z(n4660) );
  NAND2_X1 U2516 ( .A1(n4660), .A2(pmp_addr_i[413]), .ZN(n1615) );
  INV_X1 U2517 ( .A(n1618), .ZN(n1625) );
  NOR2_X1 U2518 ( .A1(n5100), .A2(n3583), .ZN(n1620) );
  AOI22_X1 U2519 ( .A1(n1620), .A2(n1619), .B1(n4631), .B2(pmp_addr_i[402]), 
        .ZN(n1624) );
  NOR2_X1 U2520 ( .A1(n5183), .A2(n3581), .ZN(n1622) );
  AOI22_X1 U2521 ( .A1(n1622), .A2(n1621), .B1(n999), .B2(pmp_addr_i[404]), 
        .ZN(n1623) );
  OAI21_X1 U2522 ( .B1(n1625), .B2(n1624), .A(n1623), .ZN(n1628) );
  NAND3_X1 U2523 ( .A1(n1628), .A2(n1627), .A3(n1626), .ZN(n1641) );
  NOR2_X1 U2524 ( .A1(n5162), .A2(n3625), .ZN(n1629) );
  AOI22_X1 U2525 ( .A1(n1630), .A2(n1629), .B1(n5111), .B2(pmp_addr_i[410]), 
        .ZN(n1637) );
  INV_X1 U2526 ( .A(pmp_addr_i[411]), .ZN(n1631) );
  NOR2_X1 U2527 ( .A1(instr_addr_o_29_), .A2(n1631), .ZN(n1633) );
  AOI22_X1 U2528 ( .A1(n1634), .A2(n1633), .B1(n4658), .B2(pmp_addr_i[412]), 
        .ZN(n1635) );
  OAI21_X1 U2529 ( .B1(n1637), .B2(n1636), .A(n1635), .ZN(n1639) );
  NAND2_X1 U2530 ( .A1(n1639), .A2(n1638), .ZN(n1640) );
  INV_X1 U2532 ( .A(pmp_cfg_i[67]), .ZN(n1742) );
  NAND2_X1 U2533 ( .A1(pmp_addr_i[259]), .A2(pmp_addr_i[260]), .ZN(n1748) );
  NAND2_X1 U2534 ( .A1(pmp_addr_i[262]), .A2(pmp_addr_i[261]), .ZN(n1645) );
  AND3_X1 U2535 ( .A1(pmp_addr_i[266]), .A2(pmp_addr_i[263]), .A3(
        pmp_addr_i[258]), .ZN(n1647) );
  AND2_X1 U2536 ( .A1(pmp_addr_i[256]), .A2(pmp_addr_i[257]), .ZN(n5732) );
  AND2_X1 U2537 ( .A1(pmp_addr_i[264]), .A2(pmp_addr_i[265]), .ZN(n1646) );
  NAND4_X1 U2538 ( .A1(n5734), .A2(n1647), .A3(n5732), .A4(n1646), .ZN(n11603)
         );
  OR2_X1 U2539 ( .A1(n11603), .A2(n1823), .ZN(n11587) );
  INV_X1 U2540 ( .A(pmp_addr_i[268]), .ZN(n1648) );
  NAND2_X1 U2541 ( .A1(n11583), .A2(pmp_addr_i[269]), .ZN(n11605) );
  INV_X1 U2542 ( .A(pmp_addr_i[270]), .ZN(n2223) );
  OR2_X1 U2543 ( .A1(n11605), .A2(n2223), .ZN(n5749) );
  INV_X1 U2544 ( .A(pmp_addr_i[271]), .ZN(n2218) );
  AND2_X1 U2545 ( .A1(pmp_cfg_i[68]), .A2(pmp_cfg_i[67]), .ZN(n5741) );
  OAI21_X1 U2546 ( .B1(n5749), .B2(n2218), .A(n5741), .ZN(n11595) );
  INV_X1 U2547 ( .A(pmp_cfg_i[68]), .ZN(n1738) );
  OR2_X1 U2548 ( .A1(n1738), .A2(pmp_cfg_i[67]), .ZN(n9009) );
  NAND2_X1 U2549 ( .A1(n5783), .A2(pmp_addr_i[284]), .ZN(n1649) );
  OAI21_X1 U2550 ( .B1(n509), .B2(n35), .A(n1649), .ZN(n8952) );
  INV_X1 U2551 ( .A(n8952), .ZN(n1650) );
  NOR2_X1 U2552 ( .A1(n4560), .A2(n1650), .ZN(n1684) );
  NAND2_X1 U2553 ( .A1(n5783), .A2(pmp_addr_i[283]), .ZN(n1651) );
  OAI21_X1 U2554 ( .B1(n584), .B2(n35), .A(n1651), .ZN(n9002) );
  INV_X1 U2555 ( .A(n9002), .ZN(n1682) );
  NOR2_X1 U2556 ( .A1(n5149), .A2(n1682), .ZN(n1652) );
  NOR2_X1 U2557 ( .A1(n1684), .A2(n1652), .ZN(n1687) );
  NAND2_X1 U2558 ( .A1(n5783), .A2(pmp_addr_i[285]), .ZN(n12111) );
  OAI21_X1 U2559 ( .B1(n603), .B2(n35), .A(n12111), .ZN(n9007) );
  INV_X1 U2560 ( .A(n7116), .ZN(n1703) );
  AOI21_X1 U2561 ( .B1(n4005), .B2(n9007), .A(n1703), .ZN(n1688) );
  NAND2_X1 U2562 ( .A1(n5783), .A2(pmp_addr_i[282]), .ZN(n1653) );
  OAI21_X1 U2563 ( .B1(n510), .B2(n35), .A(n1653), .ZN(n8951) );
  INV_X1 U2564 ( .A(n8951), .ZN(n1654) );
  OR2_X1 U2565 ( .A1(n5368), .A2(n1654), .ZN(n1678) );
  NAND2_X1 U2566 ( .A1(n5783), .A2(pmp_addr_i[281]), .ZN(n1655) );
  OAI21_X1 U2567 ( .B1(n581), .B2(n35), .A(n1655), .ZN(n8960) );
  NAND2_X1 U2568 ( .A1(n4147), .A2(n8960), .ZN(n1656) );
  NAND4_X1 U2569 ( .A1(n1687), .A2(n1688), .A3(n1678), .A4(n1656), .ZN(n1718)
         );
  NAND2_X1 U2570 ( .A1(n5783), .A2(pmp_addr_i[277]), .ZN(n1657) );
  OAI21_X1 U2571 ( .B1(n594), .B2(n35), .A(n1657), .ZN(n8958) );
  INV_X1 U2572 ( .A(n8958), .ZN(n1695) );
  INV_X2 U2573 ( .A(n1658), .ZN(n6025) );
  NAND2_X1 U2574 ( .A1(n5783), .A2(pmp_addr_i[280]), .ZN(n1659) );
  OAI21_X1 U2575 ( .B1(n513), .B2(n35), .A(n1659), .ZN(n8950) );
  INV_X1 U2576 ( .A(n8950), .ZN(n1660) );
  NOR2_X1 U2577 ( .A1(instr_addr_o_26_), .A2(n1660), .ZN(n1700) );
  NAND2_X1 U2578 ( .A1(n5783), .A2(pmp_addr_i[279]), .ZN(n1661) );
  OAI21_X1 U2579 ( .B1(n597), .B2(n35), .A(n1661), .ZN(n8996) );
  INV_X1 U2580 ( .A(n8996), .ZN(n1698) );
  NOR2_X1 U2581 ( .A1(n4644), .A2(n1698), .ZN(n1662) );
  NAND2_X1 U2582 ( .A1(n5783), .A2(pmp_addr_i[278]), .ZN(n1663) );
  OAI21_X1 U2583 ( .B1(n515), .B2(n35), .A(n1663), .ZN(n8995) );
  INV_X1 U2584 ( .A(n8995), .ZN(n1664) );
  OR2_X1 U2585 ( .A1(n5330), .A2(n1664), .ZN(n1694) );
  OAI211_X1 U2586 ( .C1(n1695), .C2(n6025), .A(n1693), .B(n1694), .ZN(n1709)
         );
  OR2_X1 U2587 ( .A1(n1718), .A2(n1709), .ZN(n1692) );
  NAND2_X1 U2588 ( .A1(n5783), .A2(pmp_addr_i[275]), .ZN(n1665) );
  OAI21_X1 U2589 ( .B1(n574), .B2(n35), .A(n1665), .ZN(n8985) );
  NOR2_X1 U2590 ( .A1(n5191), .A2(n8909), .ZN(n1668) );
  NAND2_X1 U2591 ( .A1(n5783), .A2(pmp_addr_i[276]), .ZN(n1666) );
  OAI21_X1 U2592 ( .B1(n517), .B2(n35), .A(n1666), .ZN(n8959) );
  INV_X1 U2593 ( .A(n8959), .ZN(n1667) );
  NOR2_X1 U2594 ( .A1(n4836), .A2(n1667), .ZN(n1674) );
  NAND2_X1 U2595 ( .A1(n5783), .A2(pmp_addr_i[274]), .ZN(n1669) );
  OAI21_X1 U2596 ( .B1(n519), .B2(n35), .A(n1669), .ZN(n9001) );
  INV_X1 U2597 ( .A(n9001), .ZN(n1670) );
  NOR2_X1 U2598 ( .A1(instr_addr_o_20_), .A2(n1670), .ZN(n1711) );
  NAND2_X1 U2599 ( .A1(n5783), .A2(pmp_addr_i[273]), .ZN(n1671) );
  OAI21_X1 U2600 ( .B1(n571), .B2(n35), .A(n1671), .ZN(n8953) );
  INV_X1 U2601 ( .A(n8953), .ZN(n1713) );
  NAND2_X1 U2602 ( .A1(n3793), .A2(n1713), .ZN(n1672) );
  OAI22_X1 U2603 ( .A1(n1711), .A2(n1672), .B1(n1996), .B2(n9001), .ZN(n1676)
         );
  NAND2_X1 U2604 ( .A1(n5191), .A2(n8909), .ZN(n1673) );
  OAI22_X1 U2605 ( .A1(n1674), .A2(n1673), .B1(n5192), .B2(n8959), .ZN(n1675)
         );
  AOI21_X1 U2606 ( .B1(n1677), .B2(n1676), .A(n1675), .ZN(n1691) );
  INV_X1 U2607 ( .A(n1678), .ZN(n1681) );
  INV_X1 U2608 ( .A(n8960), .ZN(n1679) );
  NAND2_X1 U2609 ( .A1(instr_addr_o_27_), .A2(n1679), .ZN(n1680) );
  OAI22_X1 U2610 ( .A1(n1681), .A2(n1680), .B1(n5111), .B2(n8951), .ZN(n1686)
         );
  NAND2_X1 U2611 ( .A1(n4900), .A2(n1682), .ZN(n1683) );
  OAI22_X1 U2612 ( .A1(n1684), .A2(n1683), .B1(n4658), .B2(n8952), .ZN(n1685)
         );
  AOI21_X1 U2613 ( .B1(n1687), .B2(n1686), .A(n1685), .ZN(n1690) );
  INV_X1 U2614 ( .A(n1688), .ZN(n1689) );
  OAI22_X1 U2615 ( .A1(n1692), .A2(n1691), .B1(n1690), .B2(n1689), .ZN(n1708)
         );
  INV_X1 U2616 ( .A(n1694), .ZN(n1697) );
  NAND2_X1 U2617 ( .A1(n5208), .A2(n1695), .ZN(n1696) );
  OAI22_X1 U2618 ( .A1(n1697), .A2(n1696), .B1(n2580), .B2(n8995), .ZN(n1702)
         );
  NAND2_X1 U2619 ( .A1(instr_addr_o_25_), .A2(n1698), .ZN(n1699) );
  OAI22_X1 U2620 ( .A1(n1700), .A2(n1699), .B1(n3806), .B2(n8950), .ZN(n1701)
         );
  AOI21_X1 U2621 ( .B1(n1693), .B2(n1702), .A(n1701), .ZN(n1706) );
  INV_X1 U2622 ( .A(n9007), .ZN(n1704) );
  NAND3_X1 U2623 ( .A1(n5136), .A2(n1704), .A3(n7116), .ZN(n1705) );
  OAI21_X1 U2624 ( .B1(n1706), .B2(n1718), .A(n1705), .ZN(n1707) );
  NOR2_X1 U2625 ( .A1(n1708), .A2(n1707), .ZN(n1788) );
  INV_X1 U2626 ( .A(n1709), .ZN(n1717) );
  INV_X2 U2627 ( .A(n2339), .ZN(n6020) );
  INV_X1 U2628 ( .A(n1711), .ZN(n1712) );
  OAI21_X1 U2629 ( .B1(n1713), .B2(n6020), .A(n1712), .ZN(n1714) );
  NOR2_X1 U2630 ( .A1(n1715), .A2(n1714), .ZN(n1716) );
  NAND2_X1 U2631 ( .A1(n1717), .A2(n1716), .ZN(n1719) );
  NOR2_X1 U2632 ( .A1(n1719), .A2(n1718), .ZN(n1785) );
  INV_X1 U2633 ( .A(pmp_addr_i[240]), .ZN(n1721) );
  NAND2_X1 U2634 ( .A1(n5783), .A2(pmp_addr_i[272]), .ZN(n1720) );
  OAI21_X1 U2635 ( .B1(n1721), .B2(n35), .A(n1720), .ZN(n8961) );
  INV_X1 U2636 ( .A(n8961), .ZN(n1722) );
  NOR2_X1 U2637 ( .A1(n6019), .A2(n1722), .ZN(n1777) );
  NAND2_X1 U2638 ( .A1(n5783), .A2(pmp_addr_i[271]), .ZN(n1723) );
  OAI21_X1 U2639 ( .B1(n501), .B2(n35), .A(n1723), .ZN(n8879) );
  INV_X1 U2640 ( .A(n8879), .ZN(n1776) );
  NOR2_X1 U2641 ( .A1(n5974), .A2(n1776), .ZN(n5810) );
  NOR2_X1 U2642 ( .A1(n1777), .A2(n5810), .ZN(n1780) );
  NAND2_X1 U2643 ( .A1(n11583), .A2(pmp_cfg_i[67]), .ZN(n1730) );
  NAND3_X1 U2644 ( .A1(n1730), .A2(pmp_addr_i[269]), .A3(pmp_cfg_i[68]), .ZN(
        n1724) );
  OAI21_X1 U2645 ( .B1(n35), .B2(n497), .A(n1724), .ZN(n8830) );
  INV_X1 U2646 ( .A(n8830), .ZN(n9008) );
  NOR2_X1 U2647 ( .A1(instr_addr_o_15_), .A2(n9008), .ZN(n5788) );
  INV_X1 U2648 ( .A(pmp_addr_i[269]), .ZN(n1725) );
  OAI211_X1 U2649 ( .C1(n1730), .C2(n1725), .A(pmp_addr_i[270]), .B(
        pmp_cfg_i[68]), .ZN(n1726) );
  OAI21_X1 U2650 ( .B1(n35), .B2(n1727), .A(n1726), .ZN(n11607) );
  INV_X1 U2651 ( .A(n11607), .ZN(n11609) );
  NOR2_X1 U2652 ( .A1(n5226), .A2(n11609), .ZN(n5806) );
  NOR2_X1 U2653 ( .A1(n5788), .A2(n5806), .ZN(n1728) );
  NAND2_X1 U2654 ( .A1(n1780), .A2(n1728), .ZN(n1782) );
  OAI21_X1 U2655 ( .B1(n11603), .B2(n1742), .A(pmp_cfg_i[68]), .ZN(n1734) );
  NAND2_X1 U2656 ( .A1(n156), .A2(pmp_addr_i[235]), .ZN(n1729) );
  OAI21_X1 U2657 ( .B1(n1734), .B2(n1823), .A(n1729), .ZN(n8837) );
  INV_X1 U2658 ( .A(n8837), .ZN(n8986) );
  NOR2_X1 U2659 ( .A1(n150), .A2(n8986), .ZN(n5815) );
  NAND3_X1 U2660 ( .A1(n1730), .A2(pmp_addr_i[268]), .A3(pmp_cfg_i[68]), .ZN(
        n1731) );
  OAI21_X1 U2661 ( .B1(n35), .B2(n526), .A(n1731), .ZN(n8838) );
  INV_X1 U2662 ( .A(n8838), .ZN(n8988) );
  NOR2_X1 U2663 ( .A1(n206), .A2(n8988), .ZN(n5799) );
  INV_X1 U2664 ( .A(pmp_addr_i[266]), .ZN(n1733) );
  NAND2_X1 U2665 ( .A1(n156), .A2(pmp_addr_i[234]), .ZN(n1732) );
  OAI21_X1 U2666 ( .B1(n1734), .B2(n1733), .A(n1732), .ZN(n8835) );
  INV_X1 U2667 ( .A(n8835), .ZN(n8987) );
  OR2_X1 U2668 ( .A1(n5245), .A2(n8987), .ZN(n5808) );
  AND2_X1 U2669 ( .A1(pmp_addr_i[257]), .A2(pmp_addr_i[258]), .ZN(n1737) );
  NAND4_X1 U2670 ( .A1(n5734), .A2(pmp_addr_i[263]), .A3(pmp_addr_i[256]), 
        .A4(n1737), .ZN(n11618) );
  INV_X1 U2671 ( .A(pmp_addr_i[264]), .ZN(n2268) );
  OR2_X1 U2672 ( .A1(n11618), .A2(n2268), .ZN(n11586) );
  OAI211_X1 U2673 ( .C1(n11586), .C2(n1742), .A(pmp_addr_i[265]), .B(
        pmp_cfg_i[68]), .ZN(n1735) );
  OAI21_X1 U2674 ( .B1(n35), .B2(n523), .A(n1735), .ZN(n8834) );
  INV_X1 U2675 ( .A(n8834), .ZN(n8979) );
  OR2_X1 U2676 ( .A1(instr_addr_o_11_), .A2(n8979), .ZN(n5803) );
  NOR2_X1 U2677 ( .A1(n1782), .A2(n1736), .ZN(n1747) );
  AND2_X1 U2678 ( .A1(pmp_cfg_i[67]), .A2(pmp_addr_i[256]), .ZN(n1758) );
  NAND2_X1 U2679 ( .A1(n1758), .A2(n1737), .ZN(n1760) );
  INV_X1 U2680 ( .A(n1760), .ZN(n1739) );
  AOI21_X1 U2681 ( .B1(n1739), .B2(n5734), .A(n1738), .ZN(n1750) );
  NAND2_X1 U2682 ( .A1(n1750), .A2(pmp_addr_i[263]), .ZN(n1740) );
  OAI21_X1 U2683 ( .B1(n35), .B2(n1741), .A(n1740), .ZN(n8859) );
  INV_X1 U2684 ( .A(n8859), .ZN(n8981) );
  NAND2_X1 U2685 ( .A1(n154), .A2(n8981), .ZN(n5765) );
  OAI211_X1 U2686 ( .C1(n11618), .C2(n1742), .A(pmp_addr_i[264]), .B(
        pmp_cfg_i[68]), .ZN(n1743) );
  OAI21_X1 U2687 ( .B1(n35), .B2(n544), .A(n1743), .ZN(n8860) );
  INV_X1 U2688 ( .A(n8860), .ZN(n8978) );
  NOR2_X1 U2689 ( .A1(n5270), .A2(n8978), .ZN(n1744) );
  NAND2_X1 U2690 ( .A1(n5270), .A2(n8978), .ZN(n5774) );
  OAI21_X1 U2691 ( .B1(n5765), .B2(n1744), .A(n5774), .ZN(n1767) );
  NOR2_X1 U2692 ( .A1(n155), .A2(n8981), .ZN(n5814) );
  NAND2_X1 U2693 ( .A1(n1745), .A2(n316), .ZN(n1746) );
  AND2_X1 U2694 ( .A1(n1747), .A2(n1746), .ZN(n1771) );
  OAI21_X1 U2695 ( .B1(n1760), .B2(n1748), .A(pmp_cfg_i[68]), .ZN(n1754) );
  INV_X1 U2696 ( .A(pmp_addr_i[261]), .ZN(n5737) );
  NAND2_X1 U2697 ( .A1(n156), .A2(pmp_addr_i[229]), .ZN(n1749) );
  OAI21_X1 U2698 ( .B1(n1754), .B2(n5737), .A(n1749), .ZN(n8857) );
  INV_X1 U2699 ( .A(n8857), .ZN(n8969) );
  NOR2_X1 U2700 ( .A1(n5268), .A2(n8969), .ZN(n5800) );
  NAND2_X1 U2701 ( .A1(n1750), .A2(pmp_addr_i[262]), .ZN(n1751) );
  OAI21_X1 U2702 ( .B1(n35), .B2(n1752), .A(n1751), .ZN(n8856) );
  INV_X1 U2703 ( .A(n8856), .ZN(n8980) );
  NOR2_X1 U2704 ( .A1(n5342), .A2(n8980), .ZN(n5801) );
  NOR2_X1 U2705 ( .A1(n5800), .A2(n5801), .ZN(n1770) );
  INV_X1 U2706 ( .A(pmp_addr_i[260]), .ZN(n5735) );
  NAND2_X1 U2707 ( .A1(n156), .A2(pmp_addr_i[228]), .ZN(n1753) );
  OAI21_X1 U2708 ( .B1(n1754), .B2(n5735), .A(n1753), .ZN(n8842) );
  INV_X1 U2709 ( .A(n8842), .ZN(n8977) );
  NOR2_X1 U2710 ( .A1(n12152), .A2(n8977), .ZN(n1764) );
  INV_X1 U2711 ( .A(pmp_addr_i[227]), .ZN(n5353) );
  NAND3_X1 U2712 ( .A1(n1760), .A2(pmp_addr_i[259]), .A3(pmp_cfg_i[68]), .ZN(
        n1755) );
  OAI21_X1 U2713 ( .B1(n35), .B2(n5353), .A(n1755), .ZN(n9014) );
  INV_X1 U2714 ( .A(n9014), .ZN(n8968) );
  NOR2_X1 U2715 ( .A1(n5280), .A2(n8968), .ZN(n1756) );
  OR2_X1 U2716 ( .A1(n1764), .A2(n1756), .ZN(n5819) );
  INV_X1 U2717 ( .A(pmp_addr_i[256]), .ZN(n2258) );
  INV_X1 U2718 ( .A(pmp_addr_i[224]), .ZN(n11035) );
  OAI22_X1 U2719 ( .A1(n9009), .A2(n2258), .B1(n35), .B2(n11035), .ZN(n8972)
         );
  INV_X1 U2720 ( .A(pmp_addr_i[225]), .ZN(n1759) );
  NAND2_X1 U2721 ( .A1(pmp_cfg_i[68]), .A2(pmp_addr_i[257]), .ZN(n1757) );
  OAI22_X1 U2722 ( .A1(n35), .A2(n1759), .B1(n1758), .B2(n1757), .ZN(n8971) );
  OR2_X1 U2723 ( .A1(n8972), .A2(n8971), .ZN(n1762) );
  NAND3_X1 U2724 ( .A1(n1760), .A2(pmp_addr_i[258]), .A3(pmp_cfg_i[68]), .ZN(
        n1761) );
  OAI21_X1 U2725 ( .B1(n35), .B2(n550), .A(n1761), .ZN(n8974) );
  NAND2_X1 U2726 ( .A1(n1762), .A2(n8974), .ZN(n1763) );
  INV_X1 U2727 ( .A(n8974), .ZN(n5786) );
  INV_X1 U2728 ( .A(n1762), .ZN(n5784) );
  AOI22_X1 U2729 ( .A1(n3836), .A2(n1763), .B1(n5786), .B2(n5784), .ZN(n1766)
         );
  NAND2_X1 U2730 ( .A1(instr_addr_o_6_), .A2(n8977), .ZN(n5764) );
  NAND2_X1 U2731 ( .A1(n5293), .A2(n8968), .ZN(n5773) );
  OR2_X1 U2732 ( .A1(n5773), .A2(n1764), .ZN(n1765) );
  OAI211_X1 U2733 ( .C1(n5819), .C2(n1766), .A(n5764), .B(n1765), .ZN(n1769)
         );
  NAND2_X1 U2734 ( .A1(n5268), .A2(n8969), .ZN(n5769) );
  NAND2_X1 U2735 ( .A1(n5269), .A2(n8980), .ZN(n5767) );
  OAI21_X1 U2736 ( .B1(n5801), .B2(n5769), .A(n5767), .ZN(n1768) );
  INV_X1 U2737 ( .A(n5808), .ZN(n1772) );
  NAND2_X1 U2738 ( .A1(instr_addr_o_11_), .A2(n8979), .ZN(n5763) );
  NAND2_X1 U2739 ( .A1(n5250), .A2(n8987), .ZN(n5776) );
  OAI21_X1 U2740 ( .B1(n1772), .B2(n5763), .A(n5776), .ZN(n1774) );
  NAND2_X1 U2741 ( .A1(n149), .A2(n8986), .ZN(n5777) );
  NAND2_X1 U2742 ( .A1(n5251), .A2(n8988), .ZN(n5770) );
  OAI21_X1 U2743 ( .B1(n5799), .B2(n5777), .A(n5770), .ZN(n1773) );
  AOI21_X1 U2744 ( .B1(n1775), .B2(n1774), .A(n1773), .ZN(n1783) );
  NAND2_X1 U2745 ( .A1(n12178), .A2(n9008), .ZN(n5766) );
  NAND2_X1 U2746 ( .A1(n5226), .A2(n11609), .ZN(n5768) );
  OAI21_X1 U2747 ( .B1(n5766), .B2(n5806), .A(n5768), .ZN(n1779) );
  NAND2_X1 U2748 ( .A1(n5974), .A2(n1776), .ZN(n5775) );
  OAI22_X1 U2749 ( .A1(n1777), .A2(n5775), .B1(n2082), .B2(n8961), .ZN(n1778)
         );
  AOI21_X1 U2750 ( .B1(n1780), .B2(n1779), .A(n1778), .ZN(n1781) );
  OAI21_X1 U2751 ( .B1(n1783), .B2(n1782), .A(n1781), .ZN(n1784) );
  NAND2_X1 U2752 ( .A1(n1785), .A2(n1784), .ZN(n1786) );
  NAND2_X1 U2753 ( .A1(instr_addr_o_6_), .A2(n5735), .ZN(n1796) );
  INV_X1 U2754 ( .A(pmp_addr_i[259]), .ZN(n1789) );
  NOR2_X1 U2755 ( .A1(n4596), .A2(n1789), .ZN(n1790) );
  AOI22_X1 U2756 ( .A1(n1796), .A2(n1790), .B1(n2611), .B2(pmp_addr_i[260]), 
        .ZN(n1800) );
  OR2_X1 U2757 ( .A1(pmp_addr_i[257]), .A2(pmp_addr_i[256]), .ZN(n1791) );
  NOR2_X1 U2758 ( .A1(n1791), .A2(pmp_addr_i[258]), .ZN(n1794) );
  INV_X1 U2759 ( .A(n1791), .ZN(n1793) );
  INV_X1 U2760 ( .A(pmp_addr_i[258]), .ZN(n1792) );
  OAI22_X1 U2761 ( .A1(n5899), .A2(n1794), .B1(n1793), .B2(n1792), .ZN(n1795)
         );
  OAI211_X1 U2762 ( .C1(pmp_addr_i[259]), .C2(n5031), .A(n1796), .B(n1795), 
        .ZN(n1799) );
  INV_X1 U2763 ( .A(pmp_addr_i[262]), .ZN(n1797) );
  NAND2_X1 U2764 ( .A1(instr_addr_o_8_), .A2(n1797), .ZN(n1802) );
  OAI21_X1 U2765 ( .B1(n3844), .B2(pmp_addr_i[261]), .A(n1802), .ZN(n1798) );
  AOI21_X1 U2766 ( .B1(n1800), .B2(n1799), .A(n1798), .ZN(n1817) );
  INV_X1 U2767 ( .A(pmp_addr_i[263]), .ZN(n1809) );
  NOR2_X1 U2768 ( .A1(n5040), .A2(n1809), .ZN(n1801) );
  NAND2_X1 U2769 ( .A1(n5270), .A2(n2268), .ZN(n1811) );
  AOI22_X1 U2770 ( .A1(n1801), .A2(n1811), .B1(n4602), .B2(pmp_addr_i[264]), 
        .ZN(n1813) );
  NAND3_X1 U2771 ( .A1(n1802), .A2(n2424), .A3(pmp_addr_i[261]), .ZN(n1804) );
  NAND2_X1 U2772 ( .A1(n4606), .A2(pmp_addr_i[262]), .ZN(n1803) );
  NAND3_X1 U2773 ( .A1(n1813), .A2(n1804), .A3(n1803), .ZN(n1816) );
  INV_X1 U2774 ( .A(pmp_addr_i[272]), .ZN(n1805) );
  NAND2_X1 U2775 ( .A1(n5047), .A2(n1805), .ZN(n1833) );
  NAND2_X1 U2776 ( .A1(n5974), .A2(n2218), .ZN(n1806) );
  AND2_X1 U2777 ( .A1(n1833), .A2(n1806), .ZN(n1831) );
  NAND2_X1 U2778 ( .A1(n5226), .A2(n2223), .ZN(n1830) );
  OAI211_X1 U2779 ( .C1(pmp_addr_i[269]), .C2(n4578), .A(n1831), .B(n1830), 
        .ZN(n1818) );
  INV_X1 U2780 ( .A(pmp_addr_i[267]), .ZN(n1823) );
  NAND2_X1 U2781 ( .A1(n149), .A2(n1823), .ZN(n1807) );
  AND2_X1 U2782 ( .A1(n1825), .A2(n1807), .ZN(n1822) );
  NAND2_X1 U2783 ( .A1(n5250), .A2(n1733), .ZN(n1821) );
  OAI211_X1 U2784 ( .C1(pmp_addr_i[265]), .C2(n5052), .A(n1822), .B(n1821), 
        .ZN(n1808) );
  NOR2_X1 U2785 ( .A1(n1818), .A2(n1808), .ZN(n1815) );
  NAND2_X1 U2786 ( .A1(instr_addr_o_9_), .A2(n1809), .ZN(n1810) );
  NAND2_X1 U2787 ( .A1(n1811), .A2(n1810), .ZN(n1812) );
  NAND2_X1 U2788 ( .A1(n1813), .A2(n1812), .ZN(n1814) );
  OAI211_X1 U2789 ( .C1(n1817), .C2(n1816), .A(n1815), .B(n1814), .ZN(n1853)
         );
  INV_X1 U2790 ( .A(n1818), .ZN(n1839) );
  INV_X1 U2791 ( .A(pmp_addr_i[265]), .ZN(n1819) );
  NOR2_X1 U2792 ( .A1(n3934), .A2(n1819), .ZN(n1820) );
  AOI22_X1 U2793 ( .A1(n1821), .A2(n1820), .B1(n5070), .B2(pmp_addr_i[266]), 
        .ZN(n1828) );
  INV_X1 U2794 ( .A(n1822), .ZN(n1827) );
  NOR2_X1 U2795 ( .A1(n149), .A2(n1823), .ZN(n1824) );
  AOI22_X1 U2796 ( .A1(n1825), .A2(n1824), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[268]), .ZN(n1826) );
  OAI21_X1 U2797 ( .B1(n1828), .B2(n1827), .A(n1826), .ZN(n1838) );
  NOR2_X1 U2798 ( .A1(n208), .A2(n1725), .ZN(n1829) );
  AOI22_X1 U2799 ( .A1(n1830), .A2(n1829), .B1(n5058), .B2(pmp_addr_i[270]), 
        .ZN(n1836) );
  INV_X1 U2800 ( .A(n1831), .ZN(n1835) );
  NOR2_X1 U2801 ( .A1(n12265), .A2(n2218), .ZN(n1832) );
  AOI22_X1 U2802 ( .A1(n1833), .A2(n1832), .B1(n2082), .B2(pmp_addr_i[272]), 
        .ZN(n1834) );
  OAI21_X1 U2803 ( .B1(n1836), .B2(n1835), .A(n1834), .ZN(n1837) );
  AOI21_X1 U2804 ( .B1(n1839), .B2(n1838), .A(n1837), .ZN(n1852) );
  INV_X1 U2805 ( .A(pmp_addr_i[284]), .ZN(n1840) );
  NAND2_X1 U2806 ( .A1(n12161), .A2(n1840), .ZN(n1880) );
  OAI21_X1 U2807 ( .B1(n4623), .B2(pmp_addr_i[283]), .A(n1880), .ZN(n1882) );
  INV_X1 U2808 ( .A(pmp_addr_i[282]), .ZN(n1841) );
  NAND2_X1 U2809 ( .A1(n5368), .A2(n1841), .ZN(n1878) );
  NAND2_X1 U2810 ( .A1(n5154), .A2(n2147), .ZN(n1884) );
  OAI211_X1 U2811 ( .C1(n5094), .C2(pmp_addr_i[281]), .A(n1878), .B(n1884), 
        .ZN(n1842) );
  NOR2_X1 U2812 ( .A1(n1882), .A2(n1842), .ZN(n1875) );
  NAND2_X1 U2813 ( .A1(n12157), .A2(n2161), .ZN(n1858) );
  INV_X1 U2814 ( .A(pmp_addr_i[275]), .ZN(n1857) );
  NAND2_X1 U2815 ( .A1(n3152), .A2(n1857), .ZN(n1843) );
  INV_X1 U2816 ( .A(pmp_addr_i[280]), .ZN(n1844) );
  NAND2_X1 U2817 ( .A1(n210), .A2(n1844), .ZN(n1870) );
  INV_X1 U2818 ( .A(pmp_addr_i[279]), .ZN(n1868) );
  NAND2_X1 U2819 ( .A1(instr_addr_o_25_), .A2(n1868), .ZN(n1845) );
  NAND2_X1 U2820 ( .A1(n1870), .A2(n1845), .ZN(n1873) );
  INV_X1 U2821 ( .A(pmp_addr_i[278]), .ZN(n1846) );
  NAND2_X1 U2822 ( .A1(n5330), .A2(n1846), .ZN(n1867) );
  OAI21_X1 U2823 ( .B1(n5086), .B2(pmp_addr_i[277]), .A(n1867), .ZN(n1847) );
  NOR2_X1 U2824 ( .A1(n1873), .A2(n1847), .ZN(n1864) );
  INV_X1 U2825 ( .A(pmp_addr_i[274]), .ZN(n1848) );
  NAND2_X1 U2826 ( .A1(n4802), .A2(n1848), .ZN(n1854) );
  NAND2_X1 U2827 ( .A1(instr_addr_o_19_), .A2(n2168), .ZN(n1849) );
  AND2_X1 U2828 ( .A1(n1854), .A2(n1849), .ZN(n1850) );
  NAND4_X1 U2829 ( .A1(n1875), .A2(n1856), .A3(n1864), .A4(n1850), .ZN(n1851)
         );
  AOI21_X1 U2830 ( .B1(n1853), .B2(n1852), .A(n1851), .ZN(n1892) );
  NOR2_X1 U2831 ( .A1(n5100), .A2(n2168), .ZN(n1855) );
  AOI22_X1 U2832 ( .A1(n1855), .A2(n1854), .B1(n2569), .B2(pmp_addr_i[274]), 
        .ZN(n1862) );
  NOR2_X1 U2833 ( .A1(n5191), .A2(n1857), .ZN(n1859) );
  AOI22_X1 U2834 ( .A1(n1859), .A2(n1858), .B1(n5192), .B2(pmp_addr_i[276]), 
        .ZN(n1860) );
  OAI21_X1 U2835 ( .B1(n1862), .B2(n1861), .A(n1860), .ZN(n1863) );
  NAND3_X1 U2836 ( .A1(n1875), .A2(n1864), .A3(n1863), .ZN(n1890) );
  INV_X1 U2837 ( .A(pmp_addr_i[277]), .ZN(n1865) );
  NOR2_X1 U2838 ( .A1(n5208), .A2(n1865), .ZN(n1866) );
  AOI22_X1 U2839 ( .A1(n1867), .A2(n1866), .B1(n2580), .B2(pmp_addr_i[278]), 
        .ZN(n1872) );
  NOR2_X1 U2840 ( .A1(n137), .A2(n1868), .ZN(n1869) );
  AOI22_X1 U2841 ( .A1(n1870), .A2(n1869), .B1(n3806), .B2(pmp_addr_i[280]), 
        .ZN(n1871) );
  OAI21_X1 U2842 ( .B1(n1873), .B2(n1872), .A(n1871), .ZN(n1874) );
  NAND2_X1 U2843 ( .A1(n1875), .A2(n1874), .ZN(n1889) );
  INV_X1 U2844 ( .A(pmp_addr_i[281]), .ZN(n1876) );
  NOR2_X1 U2845 ( .A1(n5162), .A2(n1876), .ZN(n1877) );
  AOI22_X1 U2846 ( .A1(n1878), .A2(n1877), .B1(n4438), .B2(pmp_addr_i[282]), 
        .ZN(n1883) );
  NOR2_X1 U2847 ( .A1(n5149), .A2(n2145), .ZN(n1879) );
  AOI22_X1 U2848 ( .A1(n1880), .A2(n1879), .B1(n5115), .B2(pmp_addr_i[284]), 
        .ZN(n1881) );
  OAI21_X1 U2849 ( .B1(n1883), .B2(n1882), .A(n1881), .ZN(n1885) );
  NAND2_X1 U2850 ( .A1(n1885), .A2(n1884), .ZN(n1888) );
  NOR2_X1 U2851 ( .A1(pmp_addr_i[286]), .A2(pmp_addr_i[287]), .ZN(n8818) );
  OAI21_X1 U2852 ( .B1(n6018), .B2(n2147), .A(n8818), .ZN(n1886) );
  INV_X1 U2853 ( .A(n1886), .ZN(n1887) );
  NAND4_X1 U2854 ( .A1(n1890), .A2(n1889), .A3(n1888), .A4(n1887), .ZN(n1891)
         );
  OR2_X1 U2855 ( .A1(n1892), .A2(n1891), .ZN(n1893) );
  NAND2_X1 U2856 ( .A1(pmp_addr_i[66]), .A2(pmp_addr_i[65]), .ZN(n1947) );
  NAND2_X1 U2857 ( .A1(pmp_addr_i[68]), .A2(pmp_addr_i[67]), .ZN(n1895) );
  NOR2_X1 U2858 ( .A1(n1947), .A2(n1895), .ZN(n1896) );
  AND2_X1 U2859 ( .A1(pmp_cfg_i[19]), .A2(pmp_addr_i[64]), .ZN(n1953) );
  AND2_X1 U2860 ( .A1(n1896), .A2(n1953), .ZN(n1946) );
  NAND2_X1 U2861 ( .A1(pmp_addr_i[69]), .A2(pmp_addr_i[70]), .ZN(n1930) );
  NAND2_X1 U2862 ( .A1(pmp_addr_i[71]), .A2(pmp_addr_i[72]), .ZN(n1897) );
  NOR2_X1 U2863 ( .A1(n1930), .A2(n1897), .ZN(n5677) );
  NAND2_X1 U2864 ( .A1(n1946), .A2(n5677), .ZN(n1918) );
  NAND2_X1 U2865 ( .A1(pmp_addr_i[73]), .A2(pmp_addr_i[74]), .ZN(n5685) );
  OAI21_X1 U2866 ( .B1(n1918), .B2(n5685), .A(pmp_cfg_i[20]), .ZN(n1903) );
  INV_X1 U2867 ( .A(pmp_addr_i[75]), .ZN(n4219) );
  INV_X1 U2868 ( .A(pmp_cfg_i[19]), .ZN(n1898) );
  OR2_X1 U2869 ( .A1(n1898), .A2(pmp_cfg_i[20]), .ZN(n5662) );
  NAND2_X1 U2870 ( .A1(n6376), .A2(pmp_addr_i[43]), .ZN(n1899) );
  OAI21_X1 U2871 ( .B1(n1903), .B2(n4219), .A(n1899), .ZN(n6243) );
  INV_X1 U2872 ( .A(n6243), .ZN(n6102) );
  NOR2_X1 U2873 ( .A1(n150), .A2(n6102), .ZN(n5657) );
  AND2_X1 U2874 ( .A1(pmp_addr_i[76]), .A2(pmp_addr_i[75]), .ZN(n1900) );
  INV_X1 U2875 ( .A(pmp_cfg_i[20]), .ZN(n1948) );
  OAI21_X1 U2876 ( .B1(n1900), .B2(n1948), .A(n1903), .ZN(n1915) );
  NAND2_X1 U2877 ( .A1(n1915), .A2(pmp_addr_i[76]), .ZN(n1901) );
  OAI21_X1 U2878 ( .B1(n5662), .B2(n2889), .A(n1901), .ZN(n6244) );
  INV_X1 U2879 ( .A(n6244), .ZN(n11184) );
  NOR2_X1 U2880 ( .A1(n206), .A2(n11184), .ZN(n5626) );
  NOR2_X1 U2881 ( .A1(n5657), .A2(n5626), .ZN(n1937) );
  INV_X1 U2882 ( .A(pmp_addr_i[74]), .ZN(n4225) );
  NAND2_X1 U2883 ( .A1(n6376), .A2(pmp_addr_i[42]), .ZN(n1902) );
  OAI21_X1 U2884 ( .B1(n1903), .B2(n4225), .A(n1902), .ZN(n6241) );
  INV_X1 U2885 ( .A(n6241), .ZN(n6090) );
  NOR2_X1 U2886 ( .A1(instr_addr_o_12_), .A2(n6090), .ZN(n5643) );
  INV_X1 U2887 ( .A(pmp_addr_i[41]), .ZN(n4981) );
  NAND3_X1 U2888 ( .A1(n1918), .A2(pmp_addr_i[73]), .A3(pmp_cfg_i[20]), .ZN(
        n1904) );
  OAI21_X1 U2889 ( .B1(n5662), .B2(n4981), .A(n1904), .ZN(n6240) );
  INV_X1 U2890 ( .A(n6240), .ZN(n6068) );
  NAND2_X1 U2891 ( .A1(instr_addr_o_11_), .A2(n6068), .ZN(n5675) );
  NAND2_X1 U2892 ( .A1(n5250), .A2(n6090), .ZN(n5699) );
  OAI21_X1 U2893 ( .B1(n5643), .B2(n5675), .A(n5699), .ZN(n1906) );
  NAND2_X1 U2894 ( .A1(n5997), .A2(n6102), .ZN(n5721) );
  NAND2_X1 U2895 ( .A1(instr_addr_o_14_), .A2(n11184), .ZN(n5716) );
  OAI21_X1 U2896 ( .B1(n5626), .B2(n5721), .A(n5716), .ZN(n1905) );
  AOI21_X1 U2897 ( .B1(n1937), .B2(n1906), .A(n1905), .ZN(n1929) );
  NAND3_X1 U2898 ( .A1(pmp_addr_i[76]), .A2(pmp_addr_i[75]), .A3(
        pmp_addr_i[77]), .ZN(n1907) );
  NOR2_X1 U2899 ( .A1(n5685), .A2(n1907), .ZN(n5695) );
  AND3_X1 U2900 ( .A1(pmp_addr_i[79]), .A2(pmp_addr_i[68]), .A3(pmp_addr_i[66]), .ZN(n1910) );
  NAND2_X1 U2901 ( .A1(pmp_addr_i[64]), .A2(pmp_addr_i[65]), .ZN(n11151) );
  NAND2_X1 U2902 ( .A1(pmp_addr_i[78]), .A2(pmp_addr_i[67]), .ZN(n1908) );
  NOR2_X1 U2903 ( .A1(n11151), .A2(n1908), .ZN(n1909) );
  NAND4_X1 U2904 ( .A1(n5695), .A2(n5677), .A3(n1910), .A4(n1909), .ZN(n1911)
         );
  AND2_X1 U2905 ( .A1(pmp_cfg_i[19]), .A2(pmp_cfg_i[20]), .ZN(n11155) );
  NAND2_X1 U2906 ( .A1(n6376), .A2(pmp_addr_i[48]), .ZN(n1912) );
  OAI21_X1 U2907 ( .B1(n5663), .B2(n2053), .A(n1912), .ZN(n6236) );
  INV_X1 U2908 ( .A(n6236), .ZN(n1913) );
  NOR2_X1 U2909 ( .A1(n6019), .A2(n1913), .ZN(n1923) );
  NAND2_X1 U2910 ( .A1(n6376), .A2(pmp_addr_i[47]), .ZN(n1914) );
  OAI21_X1 U2911 ( .B1(n5663), .B2(n2081), .A(n1914), .ZN(n6237) );
  INV_X1 U2912 ( .A(n6237), .ZN(n6101) );
  NOR2_X1 U2913 ( .A1(n5974), .A2(n6101), .ZN(n5647) );
  INV_X1 U2915 ( .A(pmp_addr_i[45]), .ZN(n2724) );
  NAND2_X1 U2916 ( .A1(n1915), .A2(pmp_addr_i[77]), .ZN(n1916) );
  OAI21_X1 U2917 ( .B1(n5662), .B2(n2724), .A(n1916), .ZN(n6234) );
  INV_X1 U2918 ( .A(n6234), .ZN(n11187) );
  NOR2_X1 U2919 ( .A1(n5057), .A2(n11187), .ZN(n5667) );
  INV_X1 U2920 ( .A(n5695), .ZN(n1917) );
  OAI211_X1 U2921 ( .C1(n1918), .C2(n1917), .A(pmp_cfg_i[20]), .B(
        pmp_addr_i[78]), .ZN(n1919) );
  OAI21_X1 U2922 ( .B1(n5662), .B2(n2891), .A(n1919), .ZN(n11196) );
  INV_X1 U2923 ( .A(n11196), .ZN(n11194) );
  INV_X1 U2925 ( .A(n1938), .ZN(n1928) );
  INV_X1 U2926 ( .A(n1921), .ZN(n1926) );
  NAND2_X1 U2927 ( .A1(n5057), .A2(n11187), .ZN(n5720) );
  NAND2_X1 U2928 ( .A1(n12265), .A2(n6101), .ZN(n5714) );
  OAI22_X1 U2929 ( .A1(n1923), .A2(n5714), .B1(n1922), .B2(n6236), .ZN(n1924)
         );
  AOI21_X1 U2930 ( .B1(n1926), .B2(n1925), .A(n1924), .ZN(n1927) );
  OAI21_X1 U2931 ( .B1(n1929), .B2(n1928), .A(n1927), .ZN(n1991) );
  NOR2_X1 U2932 ( .A1(n6002), .A2(n6068), .ZN(n5625) );
  NOR2_X1 U2933 ( .A1(n5625), .A2(n5643), .ZN(n1936) );
  INV_X1 U2934 ( .A(pmp_addr_i[39]), .ZN(n2697) );
  INV_X1 U2935 ( .A(n1930), .ZN(n1931) );
  AOI21_X1 U2936 ( .B1(n1946), .B2(n1931), .A(n1948), .ZN(n1941) );
  NAND2_X1 U2937 ( .A1(n1941), .A2(pmp_addr_i[71]), .ZN(n1932) );
  OAI21_X1 U2938 ( .B1(n5662), .B2(n2697), .A(n1932), .ZN(n6266) );
  INV_X1 U2939 ( .A(n6266), .ZN(n6104) );
  INV_X1 U2940 ( .A(pmp_addr_i[40]), .ZN(n4937) );
  NOR2_X1 U2941 ( .A1(n1948), .A2(pmp_addr_i[71]), .ZN(n1933) );
  OAI21_X1 U2942 ( .B1(n1941), .B2(n1933), .A(pmp_addr_i[72]), .ZN(n1934) );
  OAI21_X1 U2943 ( .B1(n5662), .B2(n4937), .A(n1934), .ZN(n6267) );
  INV_X1 U2944 ( .A(n6267), .ZN(n6105) );
  OAI22_X1 U2945 ( .A1(n155), .A2(n6104), .B1(n214), .B2(n6105), .ZN(n5634) );
  NAND2_X1 U2946 ( .A1(n5270), .A2(n6105), .ZN(n5703) );
  NAND2_X1 U2947 ( .A1(n5634), .A2(n5703), .ZN(n1935) );
  NAND2_X1 U2948 ( .A1(pmp_cfg_i[20]), .A2(pmp_addr_i[69]), .ZN(n1940) );
  NAND2_X1 U2949 ( .A1(n6376), .A2(pmp_addr_i[37]), .ZN(n1939) );
  OAI21_X1 U2950 ( .B1(n1946), .B2(n1940), .A(n1939), .ZN(n6270) );
  INV_X1 U2951 ( .A(n6270), .ZN(n6093) );
  NOR2_X1 U2952 ( .A1(n5268), .A2(n6093), .ZN(n5624) );
  INV_X1 U2953 ( .A(pmp_addr_i[38]), .ZN(n1943) );
  NAND2_X1 U2954 ( .A1(n1941), .A2(pmp_addr_i[70]), .ZN(n1942) );
  OAI21_X1 U2955 ( .B1(n5662), .B2(n1943), .A(n1942), .ZN(n6269) );
  INV_X1 U2956 ( .A(n6269), .ZN(n6106) );
  NOR2_X1 U2957 ( .A1(n5342), .A2(n6106), .ZN(n5627) );
  NOR2_X1 U2958 ( .A1(n5624), .A2(n5627), .ZN(n1964) );
  NAND2_X1 U2959 ( .A1(pmp_cfg_i[20]), .A2(pmp_addr_i[68]), .ZN(n1945) );
  NAND2_X1 U2960 ( .A1(n6376), .A2(pmp_addr_i[36]), .ZN(n1944) );
  OAI21_X1 U2961 ( .B1(n1946), .B2(n1945), .A(n1944), .ZN(n6249) );
  INV_X1 U2962 ( .A(n6249), .ZN(n6094) );
  OR2_X1 U2963 ( .A1(n12152), .A2(n6094), .ZN(n1960) );
  INV_X1 U2964 ( .A(n1960), .ZN(n5656) );
  INV_X1 U2965 ( .A(pmp_addr_i[35]), .ZN(n2693) );
  INV_X1 U2966 ( .A(n1947), .ZN(n1949) );
  AOI21_X1 U2967 ( .B1(n1949), .B2(n1953), .A(n1948), .ZN(n1955) );
  NAND2_X1 U2968 ( .A1(n1955), .A2(pmp_addr_i[67]), .ZN(n1950) );
  OAI21_X1 U2969 ( .B1(n5662), .B2(n2693), .A(n1950), .ZN(n6248) );
  INV_X1 U2970 ( .A(n6248), .ZN(n6095) );
  NAND2_X1 U2971 ( .A1(n5293), .A2(n6095), .ZN(n5710) );
  NAND2_X1 U2972 ( .A1(n12152), .A2(n6094), .ZN(n5719) );
  INV_X1 U2973 ( .A(pmp_addr_i[32]), .ZN(n11482) );
  NAND2_X1 U2974 ( .A1(n6096), .A2(pmp_addr_i[64]), .ZN(n1951) );
  OAI21_X1 U2975 ( .B1(n5662), .B2(n11482), .A(n1951), .ZN(n6251) );
  INV_X1 U2976 ( .A(pmp_addr_i[33]), .ZN(n1954) );
  NAND2_X1 U2977 ( .A1(pmp_cfg_i[20]), .A2(pmp_addr_i[65]), .ZN(n1952) );
  OAI22_X1 U2978 ( .A1(n5662), .A2(n1954), .B1(n1953), .B2(n1952), .ZN(n6252)
         );
  NOR2_X1 U2979 ( .A1(n6251), .A2(n6252), .ZN(n5664) );
  INV_X1 U2980 ( .A(n5664), .ZN(n1959) );
  INV_X1 U2981 ( .A(pmp_addr_i[34]), .ZN(n2683) );
  NAND2_X1 U2982 ( .A1(n1955), .A2(pmp_addr_i[66]), .ZN(n1956) );
  OAI21_X1 U2983 ( .B1(n5662), .B2(n2683), .A(n1956), .ZN(n6257) );
  OAI21_X1 U2985 ( .B1(n6258), .B2(n5664), .A(n5291), .ZN(n1958) );
  OR2_X1 U2986 ( .A1(n5293), .A2(n6095), .ZN(n5648) );
  OAI211_X1 U2987 ( .C1(n5656), .C2(n5710), .A(n5719), .B(n1961), .ZN(n1963)
         );
  NAND2_X1 U2988 ( .A1(n5268), .A2(n6093), .ZN(n5718) );
  NAND2_X1 U2989 ( .A1(n5269), .A2(n6106), .ZN(n5694) );
  AND2_X1 U2990 ( .A1(n5694), .A2(n5703), .ZN(n5723) );
  NAND2_X1 U2991 ( .A1(instr_addr_o_9_), .A2(n6104), .ZN(n5711) );
  OAI211_X1 U2992 ( .C1(n5627), .C2(n5718), .A(n5723), .B(n5711), .ZN(n1962)
         );
  AOI21_X1 U2993 ( .B1(n1964), .B2(n1963), .A(n1962), .ZN(n1965) );
  NOR2_X1 U2994 ( .A1(n1966), .A2(n1965), .ZN(n1990) );
  INV_X1 U2995 ( .A(pmp_addr_i[88]), .ZN(n4283) );
  NAND2_X1 U2996 ( .A1(n6376), .A2(pmp_addr_i[56]), .ZN(n1967) );
  OAI21_X1 U2997 ( .B1(n5663), .B2(n4283), .A(n1967), .ZN(n6307) );
  NOR2_X1 U2998 ( .A1(instr_addr_o_26_), .A2(n6344), .ZN(n2024) );
  INV_X1 U2999 ( .A(pmp_addr_i[87]), .ZN(n4285) );
  NAND2_X1 U3000 ( .A1(n6376), .A2(pmp_addr_i[55]), .ZN(n1968) );
  OAI21_X1 U3001 ( .B1(n5663), .B2(n4285), .A(n1968), .ZN(n6306) );
  NOR2_X1 U3002 ( .A1(n4644), .A2(n6343), .ZN(n1969) );
  OR2_X1 U3003 ( .A1(n2024), .A2(n1969), .ZN(n2019) );
  INV_X1 U3004 ( .A(pmp_addr_i[85]), .ZN(n4280) );
  NAND2_X1 U3005 ( .A1(n6376), .A2(pmp_addr_i[53]), .ZN(n1970) );
  OAI21_X1 U3006 ( .B1(n5663), .B2(n4280), .A(n1970), .ZN(n6303) );
  INV_X1 U3007 ( .A(n6303), .ZN(n6082) );
  INV_X1 U3008 ( .A(pmp_addr_i[86]), .ZN(n4278) );
  NAND2_X1 U3009 ( .A1(n6376), .A2(pmp_addr_i[54]), .ZN(n1971) );
  OAI21_X1 U3010 ( .B1(n5663), .B2(n4278), .A(n1971), .ZN(n6304) );
  INV_X1 U3011 ( .A(n6304), .ZN(n6083) );
  OR2_X1 U3012 ( .A1(n5330), .A2(n6083), .ZN(n2020) );
  OAI21_X1 U3013 ( .B1(n5208), .B2(n6082), .A(n2020), .ZN(n1972) );
  INV_X1 U3014 ( .A(pmp_addr_i[83]), .ZN(n4273) );
  NAND2_X1 U3015 ( .A1(n6376), .A2(pmp_addr_i[51]), .ZN(n1973) );
  OAI21_X1 U3016 ( .B1(n5663), .B2(n4273), .A(n1973), .ZN(n6310) );
  INV_X1 U3017 ( .A(n6310), .ZN(n6078) );
  INV_X1 U3018 ( .A(pmp_addr_i[84]), .ZN(n4271) );
  NAND2_X1 U3019 ( .A1(n6376), .A2(pmp_addr_i[52]), .ZN(n1974) );
  OAI21_X1 U3020 ( .B1(n5663), .B2(n4271), .A(n1974), .ZN(n6311) );
  INV_X1 U3021 ( .A(n6311), .ZN(n6079) );
  OR2_X1 U3022 ( .A1(n5181), .A2(n6079), .ZN(n1999) );
  OAI21_X1 U3023 ( .B1(n5183), .B2(n6078), .A(n1999), .ZN(n1994) );
  INV_X1 U3024 ( .A(pmp_addr_i[81]), .ZN(n4268) );
  NAND2_X1 U3025 ( .A1(n6376), .A2(pmp_addr_i[49]), .ZN(n1975) );
  OAI21_X1 U3026 ( .B1(n5663), .B2(n4268), .A(n1975), .ZN(n6313) );
  INV_X1 U3027 ( .A(pmp_addr_i[82]), .ZN(n4266) );
  NAND2_X1 U3028 ( .A1(n6376), .A2(pmp_addr_i[50]), .ZN(n1976) );
  INV_X1 U3029 ( .A(n6314), .ZN(n1977) );
  OR2_X1 U3030 ( .A1(n5187), .A2(n1977), .ZN(n1995) );
  OAI21_X1 U3031 ( .B1(n5100), .B2(n6330), .A(n1995), .ZN(n1978) );
  NOR2_X1 U3032 ( .A1(n1994), .A2(n1978), .ZN(n1979) );
  NAND2_X1 U3033 ( .A1(n1992), .A2(n1979), .ZN(n1988) );
  INV_X1 U3034 ( .A(pmp_addr_i[92]), .ZN(n4290) );
  NAND2_X1 U3035 ( .A1(n6376), .A2(pmp_addr_i[60]), .ZN(n1980) );
  OAI21_X1 U3036 ( .B1(n5663), .B2(n4290), .A(n1980), .ZN(n6322) );
  INV_X1 U3037 ( .A(n6322), .ZN(n1981) );
  NOR2_X1 U3038 ( .A1(n4560), .A2(n1981), .ZN(n2010) );
  INV_X1 U3039 ( .A(pmp_addr_i[91]), .ZN(n4292) );
  NAND2_X1 U3040 ( .A1(n6376), .A2(pmp_addr_i[59]), .ZN(n1982) );
  OAI21_X1 U3041 ( .B1(n5663), .B2(n4292), .A(n1982), .ZN(n6321) );
  INV_X1 U3042 ( .A(n6321), .ZN(n6075) );
  NOR2_X1 U3043 ( .A1(n5149), .A2(n6075), .ZN(n1983) );
  NOR2_X1 U3044 ( .A1(n2010), .A2(n1983), .ZN(n2013) );
  INV_X1 U3045 ( .A(pmp_addr_i[61]), .ZN(n2758) );
  INV_X1 U3046 ( .A(pmp_addr_i[93]), .ZN(n12071) );
  OR2_X1 U3047 ( .A1(n5663), .A2(n12071), .ZN(n11204) );
  OAI21_X1 U3048 ( .B1(n5662), .B2(n2758), .A(n11204), .ZN(n6325) );
  OR2_X1 U3049 ( .A1(pmp_addr_i[62]), .A2(pmp_addr_i[63]), .ZN(n2028) );
  AOI21_X1 U3050 ( .B1(n4005), .B2(n6325), .A(n2028), .ZN(n2014) );
  INV_X1 U3051 ( .A(pmp_addr_i[90]), .ZN(n4297) );
  NAND2_X1 U3052 ( .A1(n6376), .A2(pmp_addr_i[58]), .ZN(n1984) );
  OAI21_X1 U3053 ( .B1(n5663), .B2(n4297), .A(n1984), .ZN(n6319) );
  INV_X1 U3054 ( .A(n6319), .ZN(n1985) );
  OR2_X1 U3055 ( .A1(n5368), .A2(n1985), .ZN(n2005) );
  INV_X1 U3056 ( .A(pmp_addr_i[89]), .ZN(n4295) );
  NAND2_X1 U3057 ( .A1(n6376), .A2(pmp_addr_i[57]), .ZN(n1986) );
  OAI21_X1 U3058 ( .B1(n5663), .B2(n4295), .A(n1986), .ZN(n6318) );
  NAND2_X1 U3059 ( .A1(n4147), .A2(n6318), .ZN(n1987) );
  NOR2_X1 U3060 ( .A1(n1988), .A2(n2030), .ZN(n1989) );
  OAI21_X1 U3061 ( .B1(n1991), .B2(n1990), .A(n1989), .ZN(n2035) );
  OR2_X1 U3062 ( .A1(n2030), .A2(n1993), .ZN(n2018) );
  INV_X1 U3063 ( .A(n1994), .ZN(n2004) );
  INV_X1 U3064 ( .A(n1995), .ZN(n1998) );
  NAND2_X1 U3065 ( .A1(n3793), .A2(n6330), .ZN(n1997) );
  OAI22_X1 U3066 ( .A1(n1998), .A2(n1997), .B1(n1996), .B2(n6314), .ZN(n2003)
         );
  INV_X1 U3067 ( .A(n1999), .ZN(n2001) );
  NAND2_X1 U3068 ( .A1(n5183), .A2(n6078), .ZN(n2000) );
  OAI22_X1 U3069 ( .A1(n2001), .A2(n2000), .B1(n999), .B2(n6311), .ZN(n2002)
         );
  AOI21_X1 U3070 ( .B1(n2004), .B2(n2003), .A(n2002), .ZN(n2017) );
  INV_X1 U3071 ( .A(n2005), .ZN(n2008) );
  INV_X1 U3072 ( .A(n6318), .ZN(n2006) );
  NAND2_X1 U3073 ( .A1(instr_addr_o_27_), .A2(n2006), .ZN(n2007) );
  OAI22_X1 U3074 ( .A1(n2008), .A2(n2007), .B1(n5111), .B2(n6319), .ZN(n2012)
         );
  NAND2_X1 U3075 ( .A1(n5550), .A2(n6075), .ZN(n2009) );
  OAI22_X1 U3076 ( .A1(n2010), .A2(n2009), .B1(n4658), .B2(n6322), .ZN(n2011)
         );
  AOI21_X1 U3077 ( .B1(n2013), .B2(n2012), .A(n2011), .ZN(n2016) );
  INV_X1 U3078 ( .A(n2014), .ZN(n2015) );
  OAI22_X1 U3079 ( .A1(n2018), .A2(n2017), .B1(n2016), .B2(n2015), .ZN(n2033)
         );
  INV_X1 U3080 ( .A(n2019), .ZN(n2027) );
  INV_X1 U3081 ( .A(n2020), .ZN(n2022) );
  NAND2_X1 U3082 ( .A1(instr_addr_o_23_), .A2(n6082), .ZN(n2021) );
  OAI22_X1 U3083 ( .A1(n2022), .A2(n2021), .B1(n2580), .B2(n6304), .ZN(n2026)
         );
  NAND2_X1 U3084 ( .A1(n5202), .A2(n6343), .ZN(n2023) );
  OAI22_X1 U3085 ( .A1(n2024), .A2(n2023), .B1(n1273), .B2(n6307), .ZN(n2025)
         );
  AOI21_X1 U3086 ( .B1(n2027), .B2(n2026), .A(n2025), .ZN(n2031) );
  INV_X1 U3087 ( .A(n6325), .ZN(n5632) );
  NAND3_X1 U3088 ( .A1(n147), .A2(n5632), .A3(n8193), .ZN(n2029) );
  OAI21_X1 U3089 ( .B1(n2031), .B2(n2030), .A(n2029), .ZN(n2032) );
  NAND2_X1 U3090 ( .A1(instr_addr_o_6_), .A2(n5676), .ZN(n2043) );
  INV_X1 U3091 ( .A(pmp_addr_i[67]), .ZN(n2036) );
  NOR2_X1 U3092 ( .A1(n4596), .A2(n2036), .ZN(n2037) );
  AOI22_X1 U3093 ( .A1(n2043), .A2(n2037), .B1(n16), .B2(pmp_addr_i[68]), .ZN(
        n2047) );
  OR2_X1 U3094 ( .A1(pmp_addr_i[65]), .A2(pmp_addr_i[64]), .ZN(n2038) );
  NOR2_X1 U3095 ( .A1(n2038), .A2(pmp_addr_i[66]), .ZN(n2041) );
  INV_X1 U3096 ( .A(n2038), .ZN(n2040) );
  INV_X1 U3097 ( .A(pmp_addr_i[66]), .ZN(n2039) );
  OAI22_X1 U3098 ( .A1(n5899), .A2(n2041), .B1(n2040), .B2(n2039), .ZN(n2042)
         );
  OAI211_X1 U3099 ( .C1(pmp_addr_i[67]), .C2(n5031), .A(n2043), .B(n2042), 
        .ZN(n2046) );
  INV_X1 U3100 ( .A(pmp_addr_i[70]), .ZN(n2044) );
  NAND2_X1 U3101 ( .A1(n5269), .A2(n2044), .ZN(n2050) );
  OAI21_X1 U3102 ( .B1(n3844), .B2(pmp_addr_i[69]), .A(n2050), .ZN(n2045) );
  AOI21_X1 U3103 ( .B1(n2047), .B2(n2046), .A(n2045), .ZN(n2066) );
  INV_X1 U3104 ( .A(pmp_addr_i[71]), .ZN(n2058) );
  NOR2_X1 U3105 ( .A1(n5040), .A2(n2058), .ZN(n2049) );
  INV_X1 U3106 ( .A(pmp_addr_i[72]), .ZN(n2048) );
  NAND2_X1 U3107 ( .A1(n5262), .A2(n2048), .ZN(n2060) );
  AOI22_X1 U3108 ( .A1(n2049), .A2(n2060), .B1(n4602), .B2(pmp_addr_i[72]), 
        .ZN(n2062) );
  NAND3_X1 U3109 ( .A1(n2050), .A2(n3844), .A3(pmp_addr_i[69]), .ZN(n2052) );
  NAND2_X1 U3110 ( .A1(n4606), .A2(pmp_addr_i[70]), .ZN(n2051) );
  NAND3_X1 U3111 ( .A1(n2062), .A2(n2052), .A3(n2051), .ZN(n2065) );
  INV_X1 U3112 ( .A(pmp_addr_i[80]), .ZN(n2053) );
  NAND2_X1 U3113 ( .A1(n5047), .A2(n2053), .ZN(n2084) );
  INV_X1 U3114 ( .A(pmp_addr_i[79]), .ZN(n2081) );
  NAND2_X1 U3115 ( .A1(n5974), .A2(n2081), .ZN(n2054) );
  AND2_X1 U3116 ( .A1(n2084), .A2(n2054), .ZN(n2080) );
  INV_X1 U3117 ( .A(pmp_addr_i[78]), .ZN(n2055) );
  NAND2_X1 U3118 ( .A1(n3100), .A2(n2055), .ZN(n2079) );
  OAI211_X1 U3119 ( .C1(pmp_addr_i[77]), .C2(n4578), .A(n2080), .B(n2079), 
        .ZN(n2067) );
  INV_X1 U3120 ( .A(pmp_addr_i[76]), .ZN(n2056) );
  NAND2_X1 U3121 ( .A1(n5251), .A2(n2056), .ZN(n2073) );
  NAND2_X1 U3122 ( .A1(n149), .A2(n4219), .ZN(n2057) );
  AND2_X1 U3123 ( .A1(n2073), .A2(n2057), .ZN(n2071) );
  NAND2_X1 U3124 ( .A1(n5250), .A2(n4225), .ZN(n2070) );
  NAND2_X1 U3125 ( .A1(instr_addr_o_9_), .A2(n2058), .ZN(n2059) );
  NAND2_X1 U3126 ( .A1(n2060), .A2(n2059), .ZN(n2061) );
  NAND2_X1 U3127 ( .A1(n2062), .A2(n2061), .ZN(n2063) );
  OAI211_X1 U3128 ( .C1(n2066), .C2(n2065), .A(n2064), .B(n2063), .ZN(n2099)
         );
  INV_X1 U3129 ( .A(n2067), .ZN(n2090) );
  INV_X1 U3130 ( .A(pmp_addr_i[73]), .ZN(n2068) );
  NOR2_X1 U3131 ( .A1(n3934), .A2(n2068), .ZN(n2069) );
  NOR2_X1 U3132 ( .A1(n149), .A2(n4219), .ZN(n2072) );
  AOI22_X1 U3133 ( .A1(n2073), .A2(n2072), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[76]), .ZN(n2074) );
  OAI21_X1 U3134 ( .B1(n2076), .B2(n2075), .A(n2074), .ZN(n2089) );
  INV_X1 U3135 ( .A(pmp_addr_i[77]), .ZN(n2077) );
  NOR2_X1 U3136 ( .A1(instr_addr_o_15_), .A2(n2077), .ZN(n2078) );
  AOI22_X1 U3137 ( .A1(n2079), .A2(n2078), .B1(n5058), .B2(pmp_addr_i[78]), 
        .ZN(n2087) );
  INV_X1 U3138 ( .A(n2080), .ZN(n2086) );
  NOR2_X1 U3139 ( .A1(n12156), .A2(n2081), .ZN(n2083) );
  AOI22_X1 U3140 ( .A1(n2084), .A2(n2083), .B1(n2082), .B2(pmp_addr_i[80]), 
        .ZN(n2085) );
  OAI21_X1 U3141 ( .B1(n2087), .B2(n2086), .A(n2085), .ZN(n2088) );
  AOI21_X1 U3142 ( .B1(n2089), .B2(n2090), .A(n2088), .ZN(n2098) );
  NAND2_X1 U3143 ( .A1(n12161), .A2(n4290), .ZN(n2122) );
  OAI21_X1 U3144 ( .B1(n4656), .B2(pmp_addr_i[91]), .A(n2122), .ZN(n2124) );
  NAND2_X1 U3145 ( .A1(n5368), .A2(n4297), .ZN(n2120) );
  NAND2_X1 U3146 ( .A1(n5154), .A2(n12071), .ZN(n2126) );
  OAI211_X1 U3147 ( .C1(n5094), .C2(pmp_addr_i[89]), .A(n2120), .B(n2126), 
        .ZN(n2091) );
  NOR2_X1 U3148 ( .A1(n2124), .A2(n2091), .ZN(n2118) );
  NAND2_X1 U3149 ( .A1(n12157), .A2(n4271), .ZN(n2104) );
  NAND2_X1 U3150 ( .A1(n3152), .A2(n4273), .ZN(n2092) );
  NAND2_X1 U3151 ( .A1(n12158), .A2(n4283), .ZN(n2114) );
  NAND2_X1 U3152 ( .A1(n5202), .A2(n4285), .ZN(n2093) );
  NAND2_X1 U3153 ( .A1(n2114), .A2(n2093), .ZN(n2116) );
  NAND2_X1 U3154 ( .A1(n5330), .A2(n4278), .ZN(n2112) );
  OAI21_X1 U3155 ( .B1(n5086), .B2(pmp_addr_i[85]), .A(n2112), .ZN(n2094) );
  NOR2_X1 U3156 ( .A1(n2116), .A2(n2094), .ZN(n2110) );
  NAND2_X1 U3157 ( .A1(n4802), .A2(n4266), .ZN(n2100) );
  NAND2_X1 U3158 ( .A1(instr_addr_o_19_), .A2(n4268), .ZN(n2095) );
  AND2_X1 U3159 ( .A1(n2100), .A2(n2095), .ZN(n2096) );
  NAND4_X1 U3160 ( .A1(n2118), .A2(n2102), .A3(n2110), .A4(n2096), .ZN(n2097)
         );
  AOI21_X1 U3161 ( .B1(n2098), .B2(n2099), .A(n2097), .ZN(n2135) );
  NOR2_X1 U3162 ( .A1(n5100), .A2(n4268), .ZN(n2101) );
  AOI22_X1 U3163 ( .A1(n2101), .A2(n2100), .B1(n1996), .B2(pmp_addr_i[82]), 
        .ZN(n2108) );
  NOR2_X1 U3164 ( .A1(n5183), .A2(n4273), .ZN(n2105) );
  AOI22_X1 U3165 ( .A1(n2105), .A2(n2104), .B1(n5192), .B2(pmp_addr_i[84]), 
        .ZN(n2106) );
  NOR2_X1 U3166 ( .A1(n5208), .A2(n4280), .ZN(n2111) );
  NOR2_X1 U3167 ( .A1(n137), .A2(n4285), .ZN(n2113) );
  AOI22_X1 U3168 ( .A1(n2114), .A2(n2113), .B1(n3806), .B2(pmp_addr_i[88]), 
        .ZN(n2115) );
  NAND2_X1 U3169 ( .A1(n2118), .A2(n2117), .ZN(n2132) );
  NOR2_X1 U3170 ( .A1(n5162), .A2(n4295), .ZN(n2119) );
  AOI22_X1 U3171 ( .A1(n2120), .A2(n2119), .B1(n5111), .B2(pmp_addr_i[90]), 
        .ZN(n2125) );
  NOR2_X1 U3172 ( .A1(n5149), .A2(n4292), .ZN(n2121) );
  AOI22_X1 U3173 ( .A1(n2122), .A2(n2121), .B1(n5115), .B2(pmp_addr_i[92]), 
        .ZN(n2123) );
  OAI21_X1 U3174 ( .B1(n2125), .B2(n2124), .A(n2123), .ZN(n2127) );
  NAND2_X1 U3175 ( .A1(n2127), .A2(n2126), .ZN(n2131) );
  NOR2_X1 U3176 ( .A1(pmp_addr_i[94]), .A2(pmp_addr_i[95]), .ZN(n2128) );
  OAI21_X1 U3177 ( .B1(n4866), .B2(n12071), .A(n2128), .ZN(n2129) );
  INV_X1 U3178 ( .A(n2129), .ZN(n2130) );
  NAND4_X1 U3179 ( .A1(n2133), .A2(n2132), .A3(n2131), .A4(n2130), .ZN(n2134)
         );
  OR2_X1 U3180 ( .A1(n2135), .A2(n2134), .ZN(n2136) );
  INV_X1 U3181 ( .A(pmp_cfg_i[75]), .ZN(n2227) );
  NAND2_X1 U3182 ( .A1(pmp_addr_i[288]), .A2(pmp_addr_i[289]), .ZN(n11835) );
  INV_X1 U3183 ( .A(pmp_addr_i[290]), .ZN(n2251) );
  OR2_X1 U3184 ( .A1(n11835), .A2(n2251), .ZN(n5425) );
  NAND2_X1 U3185 ( .A1(pmp_addr_i[292]), .A2(pmp_addr_i[291]), .ZN(n2236) );
  NOR2_X1 U3186 ( .A1(n5425), .A2(n2236), .ZN(n11842) );
  NAND2_X1 U3187 ( .A1(n11842), .A2(pmp_addr_i[293]), .ZN(n11849) );
  INV_X1 U3188 ( .A(pmp_addr_i[294]), .ZN(n2137) );
  OR2_X1 U3189 ( .A1(n11849), .A2(n2137), .ZN(n11850) );
  INV_X1 U3190 ( .A(pmp_addr_i[295]), .ZN(n2138) );
  NOR2_X1 U3191 ( .A1(n11850), .A2(n2138), .ZN(n11838) );
  NAND2_X1 U3192 ( .A1(n11838), .A2(pmp_addr_i[296]), .ZN(n11852) );
  OR2_X1 U3193 ( .A1(n11852), .A2(n2139), .ZN(n11862) );
  AND2_X1 U3194 ( .A1(pmp_addr_i[298]), .A2(pmp_addr_i[300]), .ZN(n2140) );
  NAND4_X1 U3195 ( .A1(n2140), .A2(pmp_addr_i[299]), .A3(pmp_addr_i[302]), 
        .A4(pmp_addr_i[301]), .ZN(n2141) );
  NOR2_X1 U3196 ( .A1(n11862), .A2(n2141), .ZN(n5417) );
  NAND2_X1 U3197 ( .A1(pmp_cfg_i[75]), .A2(pmp_cfg_i[76]), .ZN(n11831) );
  AOI21_X1 U3198 ( .B1(n5417), .B2(pmp_addr_i[303]), .A(n11831), .ZN(n5427) );
  INV_X1 U3199 ( .A(pmp_cfg_i[76]), .ZN(n2253) );
  NOR2_X1 U3200 ( .A1(n2253), .A2(pmp_cfg_i[75]), .ZN(n6985) );
  OR2_X1 U3201 ( .A1(n5427), .A2(n6985), .ZN(n5469) );
  NAND2_X1 U3202 ( .A1(n5469), .A2(pmp_addr_i[316]), .ZN(n2142) );
  OAI21_X1 U3203 ( .B1(n2219), .B2(n1840), .A(n2142), .ZN(n6972) );
  INV_X1 U3204 ( .A(n6972), .ZN(n2143) );
  NOR2_X1 U3205 ( .A1(n12263), .A2(n2143), .ZN(n2180) );
  INV_X1 U3206 ( .A(pmp_addr_i[283]), .ZN(n2145) );
  NAND2_X1 U3207 ( .A1(n5469), .A2(pmp_addr_i[315]), .ZN(n2144) );
  OAI21_X1 U3208 ( .B1(n2219), .B2(n2145), .A(n2144), .ZN(n6971) );
  NOR2_X1 U3209 ( .A1(n5149), .A2(n6916), .ZN(n2146) );
  NOR2_X1 U3210 ( .A1(n2180), .A2(n2146), .ZN(n2183) );
  INV_X1 U3211 ( .A(pmp_addr_i[285]), .ZN(n2147) );
  NAND2_X1 U3212 ( .A1(n5469), .A2(pmp_addr_i[317]), .ZN(n11944) );
  OAI21_X1 U3213 ( .B1(n2147), .B2(n2219), .A(n11944), .ZN(n7004) );
  OR2_X1 U3214 ( .A1(pmp_addr_i[287]), .A2(pmp_addr_i[286]), .ZN(n2199) );
  AOI21_X1 U3215 ( .B1(n4660), .B2(n7004), .A(n2199), .ZN(n2184) );
  NAND2_X1 U3216 ( .A1(n5469), .A2(pmp_addr_i[314]), .ZN(n2148) );
  OAI21_X1 U3217 ( .B1(n2219), .B2(n1841), .A(n2148), .ZN(n6970) );
  INV_X1 U3218 ( .A(n6970), .ZN(n2149) );
  OR2_X1 U3219 ( .A1(n5368), .A2(n2149), .ZN(n2175) );
  NAND2_X1 U3220 ( .A1(n5469), .A2(pmp_addr_i[313]), .ZN(n2150) );
  OAI21_X1 U3221 ( .B1(n2219), .B2(n1876), .A(n2150), .ZN(n6969) );
  NAND2_X1 U3222 ( .A1(n4652), .A2(n6969), .ZN(n2151) );
  NAND2_X1 U3223 ( .A1(n5469), .A2(pmp_addr_i[309]), .ZN(n2152) );
  OAI21_X1 U3224 ( .B1(n2219), .B2(n1865), .A(n2152), .ZN(n6961) );
  INV_X1 U3225 ( .A(n6961), .ZN(n2190) );
  NAND2_X1 U3226 ( .A1(n5469), .A2(pmp_addr_i[312]), .ZN(n2153) );
  OAI21_X1 U3227 ( .B1(n2219), .B2(n1844), .A(n2153), .ZN(n6964) );
  INV_X1 U3228 ( .A(n6964), .ZN(n2154) );
  NOR2_X1 U3229 ( .A1(n12158), .A2(n2154), .ZN(n2195) );
  NAND2_X1 U3230 ( .A1(n5469), .A2(pmp_addr_i[311]), .ZN(n2155) );
  OAI21_X1 U3231 ( .B1(n2219), .B2(n1868), .A(n2155), .ZN(n6963) );
  INV_X1 U3232 ( .A(n6963), .ZN(n2193) );
  NOR2_X1 U3233 ( .A1(n136), .A2(n2193), .ZN(n2157) );
  NOR2_X1 U3234 ( .A1(n2195), .A2(n2157), .ZN(n2198) );
  NAND2_X1 U3235 ( .A1(n5469), .A2(pmp_addr_i[310]), .ZN(n2158) );
  OAI21_X1 U3236 ( .B1(n2219), .B2(n1846), .A(n2158), .ZN(n6962) );
  INV_X1 U3237 ( .A(n6962), .ZN(n2159) );
  OR2_X1 U3238 ( .A1(n5330), .A2(n2159), .ZN(n2189) );
  OAI211_X1 U3239 ( .C1(n5208), .C2(n2190), .A(n2198), .B(n2189), .ZN(n2211)
         );
  OR2_X1 U3240 ( .A1(n2211), .A2(n2214), .ZN(n2188) );
  INV_X1 U3241 ( .A(pmp_addr_i[276]), .ZN(n2161) );
  NAND2_X1 U3242 ( .A1(n5469), .A2(pmp_addr_i[308]), .ZN(n2160) );
  OAI21_X1 U3243 ( .B1(n2219), .B2(n2161), .A(n2160), .ZN(n6956) );
  INV_X1 U3244 ( .A(n6956), .ZN(n2162) );
  NOR2_X1 U3245 ( .A1(n12157), .A2(n2162), .ZN(n2172) );
  NAND2_X1 U3246 ( .A1(n5469), .A2(pmp_addr_i[307]), .ZN(n2163) );
  OAI21_X1 U3247 ( .B1(n2219), .B2(n1857), .A(n2163), .ZN(n6955) );
  INV_X1 U3248 ( .A(n6955), .ZN(n2170) );
  NOR2_X1 U3249 ( .A1(n5842), .A2(n2170), .ZN(n2164) );
  NOR2_X1 U3250 ( .A1(n2172), .A2(n2164), .ZN(n2205) );
  NAND2_X1 U3251 ( .A1(n5469), .A2(pmp_addr_i[306]), .ZN(n2165) );
  OAI21_X1 U3252 ( .B1(n2219), .B2(n1848), .A(n2165), .ZN(n6954) );
  INV_X1 U3253 ( .A(n6954), .ZN(n2166) );
  NOR2_X1 U3254 ( .A1(instr_addr_o_20_), .A2(n2166), .ZN(n2206) );
  INV_X1 U3255 ( .A(pmp_addr_i[273]), .ZN(n2168) );
  NAND2_X1 U3256 ( .A1(n5469), .A2(pmp_addr_i[305]), .ZN(n2167) );
  OAI21_X1 U3257 ( .B1(n2219), .B2(n2168), .A(n2167), .ZN(n6953) );
  INV_X1 U3258 ( .A(n6953), .ZN(n2208) );
  NAND2_X1 U3259 ( .A1(n3793), .A2(n2208), .ZN(n2169) );
  OAI22_X1 U3260 ( .A1(n2206), .A2(n2169), .B1(n2569), .B2(n6954), .ZN(n2174)
         );
  NAND2_X1 U3261 ( .A1(n5183), .A2(n2170), .ZN(n2171) );
  OAI22_X1 U3262 ( .A1(n2172), .A2(n2171), .B1(n999), .B2(n6956), .ZN(n2173)
         );
  AOI21_X1 U3263 ( .B1(n2205), .B2(n2174), .A(n2173), .ZN(n2187) );
  INV_X1 U3264 ( .A(n2175), .ZN(n2178) );
  INV_X1 U3265 ( .A(n6969), .ZN(n2176) );
  NAND2_X1 U3266 ( .A1(instr_addr_o_27_), .A2(n2176), .ZN(n2177) );
  OAI22_X1 U3267 ( .A1(n2178), .A2(n2177), .B1(n5111), .B2(n6970), .ZN(n2182)
         );
  NAND2_X1 U3268 ( .A1(n5550), .A2(n6916), .ZN(n2179) );
  OAI22_X1 U3269 ( .A1(n2180), .A2(n2179), .B1(n5115), .B2(n6972), .ZN(n2181)
         );
  AOI21_X1 U3270 ( .B1(n2183), .B2(n2182), .A(n2181), .ZN(n2186) );
  INV_X1 U3271 ( .A(n2184), .ZN(n2185) );
  OAI22_X1 U3272 ( .A1(n2188), .A2(n2187), .B1(n2186), .B2(n2185), .ZN(n2204)
         );
  INV_X1 U3273 ( .A(n2189), .ZN(n2192) );
  NAND2_X1 U3274 ( .A1(n5208), .A2(n2190), .ZN(n2191) );
  OAI22_X1 U3275 ( .A1(n2192), .A2(n2191), .B1(n1269), .B2(n6962), .ZN(n2197)
         );
  NAND2_X1 U3276 ( .A1(n5202), .A2(n2193), .ZN(n2194) );
  OAI22_X1 U3277 ( .A1(n2195), .A2(n2194), .B1(n1273), .B2(n6964), .ZN(n2196)
         );
  AOI21_X1 U3278 ( .B1(n2198), .B2(n2197), .A(n2196), .ZN(n2202) );
  INV_X1 U3279 ( .A(n7004), .ZN(n2200) );
  NAND3_X1 U3280 ( .A1(n4866), .A2(n2200), .A3(n6929), .ZN(n2201) );
  OAI21_X1 U3281 ( .B1(n2202), .B2(n2214), .A(n2201), .ZN(n2203) );
  NOR2_X1 U3282 ( .A1(n2204), .A2(n2203), .ZN(n2295) );
  INV_X1 U3283 ( .A(n2205), .ZN(n2210) );
  INV_X1 U3284 ( .A(n2206), .ZN(n2207) );
  OAI21_X1 U3285 ( .B1(instr_addr_o_19_), .B2(n2208), .A(n2207), .ZN(n2209) );
  NOR2_X1 U3286 ( .A1(n2210), .A2(n2209), .ZN(n2213) );
  INV_X1 U3287 ( .A(n2211), .ZN(n2212) );
  NAND2_X1 U3288 ( .A1(n5469), .A2(pmp_addr_i[304]), .ZN(n2215) );
  OAI21_X1 U3289 ( .B1(n2219), .B2(n1805), .A(n2215), .ZN(n6948) );
  INV_X1 U3290 ( .A(n6948), .ZN(n2216) );
  NOR2_X1 U3291 ( .A1(n6019), .A2(n2216), .ZN(n2284) );
  NAND2_X1 U3292 ( .A1(n5469), .A2(pmp_addr_i[303]), .ZN(n2217) );
  OAI21_X1 U3293 ( .B1(n2219), .B2(n2218), .A(n2217), .ZN(n6947) );
  INV_X1 U3294 ( .A(n6947), .ZN(n2283) );
  NOR2_X1 U3295 ( .A1(n5062), .A2(n2283), .ZN(n5505) );
  NOR2_X1 U3296 ( .A1(n2284), .A2(n5505), .ZN(n2287) );
  INV_X1 U3297 ( .A(pmp_addr_i[298]), .ZN(n2234) );
  OR2_X1 U3298 ( .A1(n11862), .A2(n2234), .ZN(n11828) );
  NOR2_X1 U3299 ( .A1(n11828), .A2(n2229), .ZN(n5414) );
  NAND2_X1 U3300 ( .A1(n5414), .A2(pmp_addr_i[300]), .ZN(n11870) );
  OAI21_X1 U3301 ( .B1(n11870), .B2(n2227), .A(pmp_cfg_i[76]), .ZN(n2232) );
  NAND2_X1 U3302 ( .A1(n6935), .A2(pmp_addr_i[269]), .ZN(n2220) );
  OAI21_X1 U3303 ( .B1(n2232), .B2(n5434), .A(n2220), .ZN(n6866) );
  INV_X1 U3304 ( .A(n6866), .ZN(n5421) );
  NOR2_X1 U3305 ( .A1(n208), .A2(n5421), .ZN(n5473) );
  NAND2_X1 U3306 ( .A1(n5434), .A2(pmp_cfg_i[76]), .ZN(n2222) );
  INV_X1 U3307 ( .A(pmp_addr_i[302]), .ZN(n2221) );
  AOI21_X1 U3308 ( .B1(n2232), .B2(n2222), .A(n2221), .ZN(n2225) );
  NOR2_X1 U3309 ( .A1(n2219), .A2(n2223), .ZN(n2224) );
  OR2_X1 U3310 ( .A1(n2225), .A2(n2224), .ZN(n11821) );
  NOR2_X1 U3311 ( .A1(n5226), .A2(n6875), .ZN(n5502) );
  NOR2_X1 U3312 ( .A1(n5473), .A2(n5502), .ZN(n2226) );
  NAND2_X1 U3313 ( .A1(n2287), .A2(n2226), .ZN(n2289) );
  OAI21_X1 U3314 ( .B1(n11828), .B2(n2227), .A(pmp_cfg_i[76]), .ZN(n2235) );
  NAND2_X1 U3315 ( .A1(n6935), .A2(pmp_addr_i[267]), .ZN(n2228) );
  OAI21_X1 U3316 ( .B1(n2235), .B2(n2229), .A(n2228), .ZN(n6862) );
  INV_X1 U3317 ( .A(n6862), .ZN(n5420) );
  NOR2_X1 U3318 ( .A1(n149), .A2(n5420), .ZN(n5492) );
  INV_X1 U3319 ( .A(pmp_addr_i[300]), .ZN(n2231) );
  NAND2_X1 U3320 ( .A1(n6935), .A2(pmp_addr_i[268]), .ZN(n2230) );
  OAI21_X1 U3321 ( .B1(n2232), .B2(n2231), .A(n2230), .ZN(n6865) );
  INV_X1 U3322 ( .A(n6865), .ZN(n2279) );
  NOR2_X1 U3323 ( .A1(n206), .A2(n2279), .ZN(n5494) );
  NOR2_X1 U3324 ( .A1(n5492), .A2(n5494), .ZN(n2282) );
  NAND2_X1 U3325 ( .A1(n6935), .A2(pmp_addr_i[266]), .ZN(n2233) );
  OAI21_X1 U3326 ( .B1(n2235), .B2(n2234), .A(n2233), .ZN(n6859) );
  INV_X1 U3327 ( .A(n6859), .ZN(n5433) );
  OR2_X1 U3328 ( .A1(n5245), .A2(n5433), .ZN(n2278) );
  INV_X1 U3329 ( .A(n2236), .ZN(n2237) );
  AOI21_X1 U3330 ( .B1(pmp_cfg_i[76]), .B2(n5425), .A(n6985), .ZN(n2252) );
  OAI21_X1 U3331 ( .B1(n2237), .B2(n2253), .A(n2252), .ZN(n2246) );
  NAND2_X1 U3332 ( .A1(pmp_addr_i[294]), .A2(pmp_addr_i[293]), .ZN(n2238) );
  AND2_X1 U3333 ( .A1(n2238), .A2(pmp_cfg_i[76]), .ZN(n2239) );
  OR2_X1 U3334 ( .A1(n2246), .A2(n2239), .ZN(n2264) );
  NOR2_X1 U3335 ( .A1(n2253), .A2(pmp_addr_i[295]), .ZN(n2240) );
  OR2_X1 U3336 ( .A1(n2264), .A2(n2240), .ZN(n2266) );
  NOR2_X1 U3337 ( .A1(n11831), .A2(pmp_addr_i[296]), .ZN(n2241) );
  OAI21_X1 U3338 ( .B1(n2266), .B2(n2241), .A(pmp_addr_i[297]), .ZN(n2242) );
  OAI21_X1 U3339 ( .B1(n2219), .B2(n1819), .A(n2242), .ZN(n6822) );
  INV_X1 U3340 ( .A(n6822), .ZN(n6982) );
  OR2_X1 U3341 ( .A1(instr_addr_o_11_), .A2(n6982), .ZN(n5495) );
  NAND3_X1 U3342 ( .A1(n2282), .A2(n2278), .A3(n5495), .ZN(n2243) );
  NOR2_X1 U3343 ( .A1(n2289), .A2(n2243), .ZN(n2277) );
  NAND2_X1 U3344 ( .A1(n2246), .A2(pmp_addr_i[293]), .ZN(n2244) );
  OAI21_X1 U3345 ( .B1(n2219), .B2(n5737), .A(n2244), .ZN(n6842) );
  INV_X1 U3346 ( .A(n6842), .ZN(n6995) );
  NOR2_X1 U3347 ( .A1(n4605), .A2(n6995), .ZN(n5493) );
  NAND2_X1 U3348 ( .A1(n2264), .A2(pmp_addr_i[294]), .ZN(n2245) );
  OAI21_X1 U3349 ( .B1(n2219), .B2(n1797), .A(n2245), .ZN(n6841) );
  INV_X1 U3350 ( .A(n6841), .ZN(n6999) );
  NOR2_X1 U3351 ( .A1(n5342), .A2(n6999), .ZN(n5496) );
  NOR2_X1 U3352 ( .A1(n5493), .A2(n5496), .ZN(n2271) );
  NAND2_X1 U3353 ( .A1(n2246), .A2(pmp_addr_i[292]), .ZN(n2247) );
  OAI21_X1 U3354 ( .B1(n2219), .B2(n5735), .A(n2247), .ZN(n6834) );
  INV_X1 U3355 ( .A(n6834), .ZN(n6937) );
  NOR2_X1 U3356 ( .A1(n12152), .A2(n6937), .ZN(n2261) );
  NAND2_X1 U3357 ( .A1(n6935), .A2(pmp_addr_i[259]), .ZN(n2248) );
  OAI21_X1 U3358 ( .B1(n2252), .B2(n89), .A(n2248), .ZN(n6833) );
  INV_X1 U3359 ( .A(n6833), .ZN(n6996) );
  OR2_X1 U3360 ( .A1(n2261), .A2(n2249), .ZN(n5484) );
  NAND2_X1 U3361 ( .A1(n6935), .A2(pmp_addr_i[258]), .ZN(n2250) );
  OAI21_X1 U3362 ( .B1(n2252), .B2(n2251), .A(n2250), .ZN(n6830) );
  INV_X1 U3363 ( .A(pmp_addr_i[257]), .ZN(n2256) );
  NOR2_X1 U3364 ( .A1(n2253), .A2(pmp_addr_i[288]), .ZN(n2254) );
  OAI21_X1 U3365 ( .B1(n6985), .B2(n2254), .A(pmp_addr_i[289]), .ZN(n2255) );
  OAI21_X1 U3366 ( .B1(n2219), .B2(n2256), .A(n2255), .ZN(n6989) );
  NAND2_X1 U3367 ( .A1(n6985), .A2(pmp_addr_i[288]), .ZN(n2257) );
  OAI21_X1 U3368 ( .B1(n2219), .B2(n2258), .A(n2257), .ZN(n6984) );
  OR2_X1 U3369 ( .A1(n6989), .A2(n6984), .ZN(n2259) );
  NAND2_X1 U3370 ( .A1(n6830), .A2(n2259), .ZN(n2260) );
  INV_X1 U3371 ( .A(n6830), .ZN(n6983) );
  INV_X1 U3372 ( .A(n2259), .ZN(n5470) );
  AOI22_X1 U3373 ( .A1(n3836), .A2(n2260), .B1(n6983), .B2(n5470), .ZN(n2263)
         );
  NAND2_X1 U3374 ( .A1(instr_addr_o_6_), .A2(n6937), .ZN(n5447) );
  NAND2_X1 U3375 ( .A1(n5293), .A2(n6996), .ZN(n5458) );
  OR2_X1 U3376 ( .A1(n5458), .A2(n2261), .ZN(n2262) );
  OAI211_X1 U3377 ( .C1(n5484), .C2(n2263), .A(n5447), .B(n2262), .ZN(n2270)
         );
  NAND2_X1 U3378 ( .A1(n5740), .A2(n6995), .ZN(n5446) );
  NAND2_X1 U3379 ( .A1(n5269), .A2(n6999), .ZN(n5452) );
  OAI21_X1 U3380 ( .B1(n5496), .B2(n5446), .A(n5452), .ZN(n2269) );
  NAND2_X1 U3381 ( .A1(n2264), .A2(pmp_addr_i[295]), .ZN(n2265) );
  OAI21_X1 U3382 ( .B1(n2219), .B2(n1809), .A(n2265), .ZN(n6844) );
  INV_X1 U3383 ( .A(n6844), .ZN(n6998) );
  NAND2_X1 U3384 ( .A1(instr_addr_o_9_), .A2(n6998), .ZN(n5457) );
  NAND2_X1 U3385 ( .A1(n2266), .A2(pmp_addr_i[296]), .ZN(n2267) );
  OAI21_X1 U3386 ( .B1(n2219), .B2(n2268), .A(n2267), .ZN(n6939) );
  INV_X1 U3387 ( .A(n6939), .ZN(n6981) );
  NOR2_X1 U3388 ( .A1(n213), .A2(n6981), .ZN(n5504) );
  NAND2_X1 U3389 ( .A1(n5270), .A2(n6981), .ZN(n5459) );
  OAI21_X1 U3390 ( .B1(n5457), .B2(n5504), .A(n5459), .ZN(n2273) );
  AOI211_X1 U3391 ( .C1(n2271), .C2(n2270), .A(n2269), .B(n2273), .ZN(n2275)
         );
  NOR2_X1 U3392 ( .A1(n4204), .A2(n6998), .ZN(n5491) );
  NOR2_X1 U3393 ( .A1(n5491), .A2(n5504), .ZN(n2272) );
  NOR2_X1 U3394 ( .A1(n2275), .A2(n2274), .ZN(n2276) );
  INV_X1 U3395 ( .A(n2278), .ZN(n5503) );
  NAND2_X1 U3396 ( .A1(instr_addr_o_11_), .A2(n6982), .ZN(n5449) );
  NAND2_X1 U3397 ( .A1(n5250), .A2(n5433), .ZN(n5451) );
  OAI21_X1 U3398 ( .B1(n5503), .B2(n5449), .A(n5451), .ZN(n2281) );
  NAND2_X1 U3399 ( .A1(n150), .A2(n5420), .ZN(n5448) );
  NAND2_X1 U3400 ( .A1(n5251), .A2(n2279), .ZN(n5453) );
  OAI21_X1 U3401 ( .B1(n5494), .B2(n5448), .A(n5453), .ZN(n2280) );
  AOI21_X1 U3402 ( .B1(n2282), .B2(n2281), .A(n2280), .ZN(n2290) );
  NAND2_X1 U3403 ( .A1(instr_addr_o_15_), .A2(n5421), .ZN(n5461) );
  OAI21_X1 U3404 ( .B1(n5502), .B2(n5461), .A(n5450), .ZN(n2286) );
  NAND2_X1 U3405 ( .A1(n12156), .A2(n2283), .ZN(n5460) );
  OAI22_X1 U3406 ( .A1(n2284), .A2(n5460), .B1(n1922), .B2(n6948), .ZN(n2285)
         );
  AOI21_X1 U3407 ( .B1(n2287), .B2(n2286), .A(n2285), .ZN(n2288) );
  OAI21_X1 U3408 ( .B1(n2290), .B2(n2289), .A(n2288), .ZN(n2291) );
  NAND2_X1 U3411 ( .A1(n5226), .A2(n2221), .ZN(n2334) );
  NOR2_X1 U3412 ( .A1(n12179), .A2(n5434), .ZN(n2296) );
  AOI22_X1 U3413 ( .A1(n2334), .A2(n2296), .B1(n5058), .B2(pmp_addr_i[302]), 
        .ZN(n2300) );
  NAND2_X1 U3414 ( .A1(n5047), .A2(n883), .ZN(n2298) );
  OAI21_X1 U3415 ( .B1(n5048), .B2(pmp_addr_i[303]), .A(n2298), .ZN(n2336) );
  NOR2_X1 U3416 ( .A1(n12156), .A2(n886), .ZN(n2297) );
  AOI22_X1 U3417 ( .A1(n2298), .A2(n2297), .B1(n2082), .B2(pmp_addr_i[304]), 
        .ZN(n2299) );
  NAND2_X1 U3419 ( .A1(n5250), .A2(n2234), .ZN(n2322) );
  NOR2_X1 U3420 ( .A1(n3934), .A2(n2139), .ZN(n2301) );
  AOI22_X1 U3421 ( .A1(n2322), .A2(n2301), .B1(n5070), .B2(pmp_addr_i[298]), 
        .ZN(n2306) );
  NAND2_X1 U3422 ( .A1(n5251), .A2(n2231), .ZN(n2304) );
  NAND2_X1 U3423 ( .A1(n4061), .A2(n2229), .ZN(n2302) );
  NAND2_X1 U3424 ( .A1(n2304), .A2(n2302), .ZN(n2324) );
  NOR2_X1 U3425 ( .A1(n149), .A2(n2229), .ZN(n2303) );
  AOI22_X1 U3426 ( .A1(n2304), .A2(n2303), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[300]), .ZN(n2305) );
  OAI21_X1 U3427 ( .B1(n2306), .B2(n2324), .A(n2305), .ZN(n2307) );
  NOR2_X1 U3428 ( .A1(n153), .A2(n2138), .ZN(n2308) );
  NAND2_X1 U3429 ( .A1(n5262), .A2(n894), .ZN(n2326) );
  AOI22_X1 U3430 ( .A1(n2308), .A2(n2326), .B1(n4602), .B2(pmp_addr_i[296]), 
        .ZN(n2328) );
  NAND2_X1 U3431 ( .A1(instr_addr_o_8_), .A2(n2137), .ZN(n2318) );
  NAND3_X1 U3432 ( .A1(n2318), .A2(n3844), .A3(pmp_addr_i[293]), .ZN(n2310) );
  NAND2_X1 U3433 ( .A1(n3894), .A2(pmp_addr_i[294]), .ZN(n2309) );
  NAND3_X1 U3434 ( .A1(n2328), .A2(n2310), .A3(n2309), .ZN(n2332) );
  INV_X1 U3435 ( .A(pmp_addr_i[292]), .ZN(n2311) );
  NAND2_X1 U3436 ( .A1(n12152), .A2(n2311), .ZN(n2317) );
  NOR2_X1 U3437 ( .A1(n20), .A2(n89), .ZN(n2312) );
  AOI22_X1 U3438 ( .A1(n2317), .A2(n2312), .B1(n2611), .B2(pmp_addr_i[292]), 
        .ZN(n2321) );
  OR2_X1 U3439 ( .A1(pmp_addr_i[289]), .A2(pmp_addr_i[288]), .ZN(n2313) );
  NOR2_X1 U3440 ( .A1(n2313), .A2(pmp_addr_i[290]), .ZN(n2315) );
  INV_X1 U3441 ( .A(n2313), .ZN(n2314) );
  OAI22_X1 U3442 ( .A1(n3836), .A2(n2315), .B1(n2314), .B2(n2251), .ZN(n2316)
         );
  OAI21_X1 U3443 ( .B1(n3844), .B2(pmp_addr_i[293]), .A(n2318), .ZN(n2319) );
  AOI21_X1 U3444 ( .B1(n2321), .B2(n2320), .A(n2319), .ZN(n2331) );
  OAI21_X1 U3445 ( .B1(n5052), .B2(pmp_addr_i[297]), .A(n2322), .ZN(n2323) );
  NOR2_X1 U3446 ( .A1(n2324), .A2(n2323), .ZN(n2330) );
  NAND2_X1 U3447 ( .A1(instr_addr_o_9_), .A2(n2138), .ZN(n2325) );
  NAND2_X1 U3448 ( .A1(n2326), .A2(n2325), .ZN(n2327) );
  NAND2_X1 U3449 ( .A1(n2328), .A2(n2327), .ZN(n2329) );
  OAI211_X1 U3450 ( .C1(n2332), .C2(n2331), .A(n2330), .B(n2329), .ZN(n2333)
         );
  OAI21_X1 U3451 ( .B1(n6017), .B2(pmp_addr_i[301]), .A(n2334), .ZN(n2335) );
  NOR2_X1 U3452 ( .A1(n2336), .A2(n2335), .ZN(n2337) );
  BUF_X2 U3453 ( .A(n3025), .Z(n5313) );
  NAND2_X1 U3454 ( .A1(n12157), .A2(n963), .ZN(n2353) );
  NAND2_X1 U3455 ( .A1(n3152), .A2(n961), .ZN(n2340) );
  AND2_X1 U3456 ( .A1(n2353), .A2(n2340), .ZN(n2352) );
  NAND2_X1 U3457 ( .A1(instr_addr_o_20_), .A2(n968), .ZN(n2350) );
  OAI211_X1 U3458 ( .C1(pmp_addr_i[305]), .C2(n12208), .A(n2352), .B(n2350), 
        .ZN(n2345) );
  INV_X1 U3459 ( .A(pmp_addr_i[312]), .ZN(n2341) );
  NAND2_X1 U3460 ( .A1(n210), .A2(n2341), .ZN(n2376) );
  INV_X1 U3461 ( .A(pmp_addr_i[311]), .ZN(n2374) );
  NAND2_X1 U3462 ( .A1(n5365), .A2(n2374), .ZN(n2342) );
  AND2_X1 U3463 ( .A1(n2376), .A2(n2342), .ZN(n2371) );
  NAND2_X1 U3464 ( .A1(n5330), .A2(n957), .ZN(n2373) );
  OAI211_X1 U3465 ( .C1(pmp_addr_i[309]), .C2(n5086), .A(n2371), .B(n2373), 
        .ZN(n2349) );
  NAND2_X1 U3466 ( .A1(n4753), .A2(n973), .ZN(n2362) );
  NAND2_X1 U3467 ( .A1(instr_addr_o_29_), .A2(n976), .ZN(n2343) );
  AND2_X1 U3468 ( .A1(n2362), .A2(n2343), .ZN(n2360) );
  NAND2_X1 U3469 ( .A1(instr_addr_o_27_), .A2(n982), .ZN(n2344) );
  NAND2_X1 U3470 ( .A1(n138), .A2(n979), .ZN(n2359) );
  NAND2_X1 U3471 ( .A1(n147), .A2(n983), .ZN(n2367) );
  NAND4_X1 U3472 ( .A1(n2360), .A2(n2344), .A3(n2359), .A4(n2367), .ZN(n2370)
         );
  NOR2_X1 U3473 ( .A1(n2349), .A2(n2370), .ZN(n2369) );
  NOR2_X1 U3474 ( .A1(n5100), .A2(n966), .ZN(n2351) );
  AOI22_X1 U3475 ( .A1(n2351), .A2(n2350), .B1(n2569), .B2(pmp_addr_i[306]), 
        .ZN(n2357) );
  INV_X1 U3476 ( .A(n2352), .ZN(n2356) );
  NOR2_X1 U3477 ( .A1(instr_addr_o_21_), .A2(n961), .ZN(n2354) );
  AOI22_X1 U3478 ( .A1(n2354), .A2(n2353), .B1(n5192), .B2(pmp_addr_i[308]), 
        .ZN(n2355) );
  OAI21_X1 U3479 ( .B1(n2357), .B2(n2356), .A(n2355), .ZN(n2368) );
  NOR2_X1 U3480 ( .A1(instr_addr_o_27_), .A2(n982), .ZN(n2358) );
  AOI22_X1 U3481 ( .A1(n2359), .A2(n2358), .B1(n5111), .B2(pmp_addr_i[314]), 
        .ZN(n2365) );
  INV_X1 U3482 ( .A(n2360), .ZN(n2364) );
  NOR2_X1 U3483 ( .A1(instr_addr_o_29_), .A2(n976), .ZN(n2361) );
  AOI22_X1 U3484 ( .A1(n2362), .A2(n2361), .B1(n5115), .B2(pmp_addr_i[316]), 
        .ZN(n2363) );
  OAI21_X1 U3485 ( .B1(n2365), .B2(n2364), .A(n2363), .ZN(n2366) );
  AOI22_X1 U3486 ( .A1(n2369), .A2(n2368), .B1(n2367), .B2(n2366), .ZN(n2384)
         );
  INV_X1 U3487 ( .A(n2370), .ZN(n2382) );
  INV_X1 U3488 ( .A(n2371), .ZN(n2379) );
  NOR2_X1 U3489 ( .A1(n6025), .A2(n955), .ZN(n2372) );
  AOI22_X1 U3490 ( .A1(n2373), .A2(n2372), .B1(n2580), .B2(pmp_addr_i[310]), 
        .ZN(n2378) );
  NOR2_X1 U3491 ( .A1(n137), .A2(n2374), .ZN(n2375) );
  AOI22_X1 U3492 ( .A1(n2376), .A2(n2375), .B1(n3806), .B2(pmp_addr_i[312]), 
        .ZN(n2377) );
  OAI21_X1 U3493 ( .B1(n2379), .B2(n2378), .A(n2377), .ZN(n2381) );
  NOR2_X1 U3494 ( .A1(pmp_addr_i[318]), .A2(pmp_addr_i[319]), .ZN(n6801) );
  OAI21_X1 U3495 ( .B1(n4866), .B2(n983), .A(n6801), .ZN(n2380) );
  NAND2_X1 U3497 ( .A1(pmp_addr_i[448]), .A2(pmp_addr_i[449]), .ZN(n3219) );
  INV_X1 U3498 ( .A(pmp_addr_i[450]), .ZN(n2391) );
  OR2_X1 U3499 ( .A1(n3219), .A2(n2391), .ZN(n3207) );
  NAND2_X1 U3500 ( .A1(pmp_addr_i[452]), .A2(pmp_addr_i[451]), .ZN(n2392) );
  NOR2_X1 U3501 ( .A1(n3207), .A2(n2392), .ZN(n11106) );
  NAND2_X1 U3502 ( .A1(n11106), .A2(pmp_addr_i[453]), .ZN(n11094) );
  NAND2_X1 U3503 ( .A1(pmp_cfg_i[115]), .A2(pmp_addr_i[454]), .ZN(n2393) );
  OAI21_X1 U3504 ( .B1(n11094), .B2(n2393), .A(pmp_cfg_i[116]), .ZN(n2401) );
  INV_X1 U3505 ( .A(pmp_addr_i[455]), .ZN(n3906) );
  INV_X1 U3506 ( .A(pmp_cfg_i[115]), .ZN(n2394) );
  NAND2_X1 U3507 ( .A1(n7923), .A2(pmp_addr_i[423]), .ZN(n2395) );
  OAI21_X1 U3508 ( .B1(n2401), .B2(n3906), .A(n2395), .ZN(n7819) );
  INV_X1 U3509 ( .A(n7819), .ZN(n7667) );
  INV_X1 U3510 ( .A(n3260), .ZN(n2398) );
  NAND2_X1 U3511 ( .A1(pmp_addr_i[454]), .A2(pmp_addr_i[455]), .ZN(n2396) );
  OR2_X1 U3512 ( .A1(n11094), .A2(n2396), .ZN(n3229) );
  NAND2_X1 U3513 ( .A1(pmp_cfg_i[115]), .A2(pmp_addr_i[456]), .ZN(n2397) );
  NOR2_X1 U3514 ( .A1(n3229), .A2(n2397), .ZN(n2452) );
  INV_X1 U3515 ( .A(pmp_cfg_i[116]), .ZN(n2450) );
  OR2_X1 U3516 ( .A1(n2452), .A2(n2450), .ZN(n2449) );
  INV_X1 U3517 ( .A(pmp_addr_i[456]), .ZN(n3903) );
  INV_X1 U3518 ( .A(pmp_addr_i[424]), .ZN(n3522) );
  OAI22_X1 U3519 ( .A1(n2449), .A2(n3903), .B1(n3522), .B2(n23), .ZN(n7821) );
  INV_X1 U3520 ( .A(n7821), .ZN(n7659) );
  INV_X1 U3521 ( .A(pmp_addr_i[454]), .ZN(n2400) );
  NAND2_X1 U3522 ( .A1(n7923), .A2(pmp_addr_i[422]), .ZN(n2399) );
  OAI21_X1 U3523 ( .B1(n2401), .B2(n2400), .A(n2399), .ZN(n7815) );
  INV_X1 U3524 ( .A(n7815), .ZN(n7632) );
  OR2_X1 U3525 ( .A1(n2623), .A2(n7632), .ZN(n3286) );
  INV_X1 U3526 ( .A(n3286), .ZN(n2425) );
  AOI21_X1 U3527 ( .B1(n11106), .B2(pmp_cfg_i[115]), .A(n2450), .ZN(n2406) );
  NAND2_X1 U3528 ( .A1(n2406), .A2(pmp_addr_i[453]), .ZN(n2402) );
  OAI21_X1 U3529 ( .B1(n23), .B2(n4604), .A(n2402), .ZN(n7817) );
  INV_X1 U3530 ( .A(n7817), .ZN(n7648) );
  NAND2_X1 U3531 ( .A1(n5740), .A2(n7648), .ZN(n3243) );
  NAND2_X1 U3532 ( .A1(n5269), .A2(n7632), .ZN(n3248) );
  OAI21_X1 U3533 ( .B1(n2425), .B2(n3243), .A(n3248), .ZN(n2405) );
  NAND2_X1 U3534 ( .A1(n155), .A2(n7667), .ZN(n3238) );
  INV_X1 U3535 ( .A(n3278), .ZN(n2403) );
  NAND2_X1 U3536 ( .A1(n5270), .A2(n7659), .ZN(n3252) );
  OAI21_X1 U3537 ( .B1(n3238), .B2(n2403), .A(n3252), .ZN(n2404) );
  INV_X1 U3539 ( .A(pmp_addr_i[420]), .ZN(n2408) );
  NAND2_X1 U3540 ( .A1(n2406), .A2(pmp_addr_i[452]), .ZN(n2407) );
  OAI21_X1 U3541 ( .B1(n23), .B2(n2408), .A(n2407), .ZN(n7798) );
  INV_X1 U3542 ( .A(n7798), .ZN(n7656) );
  INV_X1 U3543 ( .A(pmp_addr_i[419]), .ZN(n3514) );
  NAND2_X1 U3544 ( .A1(n3207), .A2(pmp_cfg_i[116]), .ZN(n2409) );
  OR2_X1 U3545 ( .A1(n2450), .A2(pmp_cfg_i[115]), .ZN(n3250) );
  NAND2_X1 U3546 ( .A1(n2409), .A2(n3250), .ZN(n2417) );
  NAND2_X1 U3547 ( .A1(n2417), .A2(pmp_addr_i[451]), .ZN(n2410) );
  OAI21_X1 U3548 ( .B1(n23), .B2(n3514), .A(n2410), .ZN(n7797) );
  INV_X1 U3549 ( .A(n7797), .ZN(n11122) );
  OR2_X1 U3550 ( .A1(instr_addr_o_5_), .A2(n11122), .ZN(n3277) );
  INV_X1 U3551 ( .A(n3277), .ZN(n2422) );
  INV_X1 U3552 ( .A(pmp_addr_i[416]), .ZN(n11977) );
  INV_X1 U3553 ( .A(pmp_addr_i[448]), .ZN(n2411) );
  OAI22_X1 U3554 ( .A1(n11977), .A2(n23), .B1(n3250), .B2(n2411), .ZN(n7800)
         );
  NAND2_X1 U3555 ( .A1(n2411), .A2(pmp_cfg_i[116]), .ZN(n2413) );
  INV_X1 U3556 ( .A(pmp_addr_i[449]), .ZN(n2412) );
  AOI21_X1 U3557 ( .B1(n3250), .B2(n2413), .A(n2412), .ZN(n2416) );
  INV_X1 U3558 ( .A(pmp_addr_i[417]), .ZN(n2414) );
  NOR2_X1 U3559 ( .A1(n23), .A2(n2414), .ZN(n2415) );
  OR2_X1 U3560 ( .A1(n2416), .A2(n2415), .ZN(n11097) );
  NOR2_X1 U3561 ( .A1(n7800), .A2(n11097), .ZN(n3266) );
  INV_X1 U3562 ( .A(n3266), .ZN(n2419) );
  INV_X1 U3563 ( .A(pmp_addr_i[418]), .ZN(n3497) );
  NAND2_X1 U3564 ( .A1(n2417), .A2(pmp_addr_i[450]), .ZN(n2418) );
  OAI21_X1 U3565 ( .B1(n3497), .B2(n23), .A(n2418), .ZN(n11101) );
  NAND2_X1 U3566 ( .A1(n2419), .A2(n11101), .ZN(n2420) );
  INV_X1 U3567 ( .A(n11101), .ZN(n11103) );
  AOI22_X1 U3568 ( .A1(n5291), .A2(n2420), .B1(n11103), .B2(n3266), .ZN(n2421)
         );
  NOR3_X1 U3569 ( .A1(n2423), .A2(n2422), .A3(n2421), .ZN(n2430) );
  AND2_X1 U3570 ( .A1(instr_addr_o_5_), .A2(n11122), .ZN(n3209) );
  NAND2_X1 U3572 ( .A1(instr_addr_o_6_), .A2(n7656), .ZN(n3241) );
  OAI21_X1 U3573 ( .B1(n2423), .B2(n3253), .A(n3241), .ZN(n2429) );
  OR2_X1 U3574 ( .A1(instr_addr_i[7]), .A2(n7648), .ZN(n3297) );
  INV_X1 U3575 ( .A(n3297), .ZN(n2426) );
  NOR2_X1 U3576 ( .A1(n2426), .A2(n2425), .ZN(n2427) );
  OAI211_X1 U3577 ( .C1(n2429), .C2(n2430), .A(n2428), .B(n2427), .ZN(n2431)
         );
  INV_X1 U3578 ( .A(pmp_addr_i[432]), .ZN(n2437) );
  NAND3_X1 U3579 ( .A1(pmp_addr_i[456]), .A2(pmp_addr_i[460]), .A3(
        pmp_addr_i[457]), .ZN(n2434) );
  NAND2_X1 U3580 ( .A1(pmp_addr_i[459]), .A2(pmp_addr_i[458]), .ZN(n2433) );
  NOR2_X1 U3581 ( .A1(n2434), .A2(n2433), .ZN(n2442) );
  NAND4_X1 U3582 ( .A1(n2442), .A2(pmp_addr_i[461]), .A3(pmp_addr_i[463]), 
        .A4(pmp_addr_i[462]), .ZN(n2435) );
  AND2_X1 U3583 ( .A1(pmp_cfg_i[115]), .A2(pmp_cfg_i[116]), .ZN(n3206) );
  OAI21_X1 U3584 ( .B1(n3229), .B2(n2435), .A(n3206), .ZN(n3208) );
  NAND2_X1 U3585 ( .A1(n3208), .A2(n3250), .ZN(n2632) );
  NAND2_X1 U3586 ( .A1(n2632), .A2(pmp_addr_i[464]), .ZN(n2436) );
  OAI21_X1 U3587 ( .B1(n23), .B2(n2437), .A(n2436), .ZN(n7786) );
  INV_X1 U3588 ( .A(n7786), .ZN(n2438) );
  NOR2_X1 U3589 ( .A1(n5047), .A2(n2438), .ZN(n2467) );
  INV_X1 U3590 ( .A(pmp_addr_i[431]), .ZN(n2440) );
  NAND2_X1 U3591 ( .A1(n2632), .A2(pmp_addr_i[463]), .ZN(n2439) );
  OAI21_X1 U3592 ( .B1(n23), .B2(n2440), .A(n2439), .ZN(n7787) );
  INV_X1 U3593 ( .A(n7787), .ZN(n7666) );
  NAND2_X1 U3594 ( .A1(n2442), .A2(pmp_cfg_i[115]), .ZN(n2443) );
  OAI21_X1 U3595 ( .B1(n3229), .B2(n2443), .A(pmp_cfg_i[116]), .ZN(n2461) );
  INV_X1 U3596 ( .A(pmp_addr_i[461]), .ZN(n3226) );
  NAND2_X1 U3597 ( .A1(n7923), .A2(pmp_addr_i[429]), .ZN(n2444) );
  OAI21_X1 U3598 ( .B1(n2461), .B2(n3226), .A(n2444), .ZN(n7784) );
  INV_X1 U3599 ( .A(n7784), .ZN(n7651) );
  INV_X1 U3600 ( .A(n3228), .ZN(n12266) );
  NAND2_X1 U3601 ( .A1(n3226), .A2(pmp_cfg_i[116]), .ZN(n2445) );
  INV_X1 U3602 ( .A(pmp_addr_i[462]), .ZN(n11133) );
  AOI21_X1 U3603 ( .B1(n2461), .B2(n2445), .A(n11133), .ZN(n2447) );
  INV_X1 U3604 ( .A(pmp_addr_i[430]), .ZN(n3507) );
  NOR2_X1 U3605 ( .A1(n23), .A2(n3507), .ZN(n2446) );
  OR2_X1 U3606 ( .A1(n2447), .A2(n2446), .ZN(n11139) );
  INV_X1 U3607 ( .A(n11139), .ZN(n7655) );
  OR2_X1 U3608 ( .A1(n12266), .A2(n7655), .ZN(n3285) );
  INV_X1 U3609 ( .A(n3285), .ZN(n2466) );
  INV_X1 U3610 ( .A(pmp_addr_i[457]), .ZN(n3933) );
  NAND2_X1 U3611 ( .A1(n7923), .A2(pmp_addr_i[425]), .ZN(n2448) );
  OAI21_X1 U3612 ( .B1(n2449), .B2(n3933), .A(n2448), .ZN(n7791) );
  INV_X1 U3613 ( .A(n7791), .ZN(n7660) );
  OR2_X1 U3614 ( .A1(instr_addr_o_11_), .A2(n7660), .ZN(n3301) );
  INV_X1 U3616 ( .A(pmp_addr_i[426]), .ZN(n3538) );
  AND2_X1 U3617 ( .A1(pmp_addr_i[458]), .A2(pmp_addr_i[457]), .ZN(n2451) );
  AOI21_X1 U3618 ( .B1(n2452), .B2(n2451), .A(n2450), .ZN(n2457) );
  NAND2_X1 U3619 ( .A1(n2457), .A2(pmp_addr_i[458]), .ZN(n2453) );
  OAI21_X1 U3620 ( .B1(n23), .B2(n3538), .A(n2453), .ZN(n2454) );
  INV_X1 U3621 ( .A(n2454), .ZN(n7646) );
  OR2_X1 U3622 ( .A1(n5250), .A2(n7646), .ZN(n3287) );
  INV_X1 U3623 ( .A(n3287), .ZN(n2455) );
  NAND2_X1 U3625 ( .A1(n2457), .A2(pmp_addr_i[459]), .ZN(n2458) );
  OAI21_X1 U3626 ( .B1(n23), .B2(n4582), .A(n2458), .ZN(n2459) );
  INV_X1 U3627 ( .A(n2459), .ZN(n7647) );
  NOR2_X1 U3628 ( .A1(n5997), .A2(n7647), .ZN(n3261) );
  INV_X1 U3629 ( .A(n3261), .ZN(n2462) );
  INV_X1 U3630 ( .A(pmp_addr_i[460]), .ZN(n3926) );
  NAND2_X1 U3631 ( .A1(n7923), .A2(pmp_addr_i[428]), .ZN(n2460) );
  OAI21_X1 U3632 ( .B1(n2461), .B2(n3926), .A(n2460), .ZN(n7793) );
  INV_X1 U3633 ( .A(n7793), .ZN(n7652) );
  OR2_X1 U3634 ( .A1(n5251), .A2(n7652), .ZN(n3300) );
  INV_X1 U3635 ( .A(n2465), .ZN(n2470) );
  NAND2_X1 U3636 ( .A1(n208), .A2(n7651), .ZN(n3239) );
  NAND2_X1 U3637 ( .A1(n12266), .A2(n7655), .ZN(n3246) );
  OAI21_X1 U3638 ( .B1(n2466), .B2(n3239), .A(n3246), .ZN(n2469) );
  NAND2_X1 U3639 ( .A1(n12156), .A2(n7666), .ZN(n3225) );
  OAI22_X1 U3640 ( .A1(n2467), .A2(n3225), .B1(instr_addr_o_18__BAR), .B2(
        n7786), .ZN(n2468) );
  NAND2_X1 U3641 ( .A1(instr_addr_o_11_), .A2(n7660), .ZN(n3240) );
  NAND2_X1 U3642 ( .A1(n5250), .A2(n7646), .ZN(n3247) );
  OAI21_X1 U3643 ( .B1(n3240), .B2(n2455), .A(n3247), .ZN(n2472) );
  INV_X1 U3644 ( .A(n3300), .ZN(n2473) );
  NAND2_X1 U3645 ( .A1(n4061), .A2(n7647), .ZN(n3242) );
  NAND2_X1 U3646 ( .A1(n206), .A2(n7652), .ZN(n3249) );
  OAI21_X1 U3647 ( .B1(n2473), .B2(n3242), .A(n3249), .ZN(n2475) );
  OAI21_X1 U3648 ( .B1(n2476), .B2(n2475), .A(n2474), .ZN(n2477) );
  INV_X1 U3649 ( .A(pmp_addr_i[440]), .ZN(n2481) );
  NAND2_X1 U3650 ( .A1(n2632), .A2(pmp_addr_i[472]), .ZN(n2480) );
  OAI21_X1 U3651 ( .B1(n23), .B2(n2481), .A(n2480), .ZN(n7856) );
  INV_X1 U3652 ( .A(n7856), .ZN(n2482) );
  NOR2_X1 U3653 ( .A1(n12158), .A2(n2482), .ZN(n2534) );
  INV_X1 U3654 ( .A(pmp_addr_i[439]), .ZN(n2484) );
  NAND2_X1 U3655 ( .A1(n2632), .A2(pmp_addr_i[471]), .ZN(n2483) );
  OAI21_X1 U3656 ( .B1(n23), .B2(n2484), .A(n2483), .ZN(n7855) );
  INV_X1 U3657 ( .A(n7855), .ZN(n2532) );
  OR2_X1 U3659 ( .A1(n2534), .A2(n2485), .ZN(n2527) );
  INV_X1 U3660 ( .A(pmp_addr_i[437]), .ZN(n2487) );
  NAND2_X1 U3661 ( .A1(n2632), .A2(pmp_addr_i[469]), .ZN(n2486) );
  OAI21_X1 U3662 ( .B1(n23), .B2(n2487), .A(n2486), .ZN(n7852) );
  INV_X1 U3663 ( .A(n7852), .ZN(n2529) );
  INV_X1 U3664 ( .A(pmp_addr_i[438]), .ZN(n2489) );
  NAND2_X1 U3665 ( .A1(n2632), .A2(pmp_addr_i[470]), .ZN(n2488) );
  OAI21_X1 U3666 ( .B1(n23), .B2(n2489), .A(n2488), .ZN(n7853) );
  INV_X1 U3667 ( .A(n7853), .ZN(n2490) );
  OR2_X1 U3668 ( .A1(n5330), .A2(n2490), .ZN(n2528) );
  OAI21_X1 U3669 ( .B1(n5208), .B2(n2529), .A(n2528), .ZN(n2491) );
  NOR2_X1 U3670 ( .A1(n2527), .A2(n2491), .ZN(n2526) );
  INV_X1 U3671 ( .A(pmp_addr_i[436]), .ZN(n2493) );
  NAND2_X1 U3672 ( .A1(n2632), .A2(pmp_addr_i[468]), .ZN(n2492) );
  OAI21_X1 U3673 ( .B1(n23), .B2(n2493), .A(n2492), .ZN(n7860) );
  INV_X1 U3674 ( .A(n7860), .ZN(n3289) );
  NOR2_X1 U3675 ( .A1(instr_addr_o_22_), .A2(n3289), .ZN(n2522) );
  INV_X1 U3676 ( .A(pmp_addr_i[435]), .ZN(n2495) );
  NAND2_X1 U3677 ( .A1(n2632), .A2(pmp_addr_i[467]), .ZN(n2494) );
  OAI21_X1 U3678 ( .B1(n23), .B2(n2495), .A(n2494), .ZN(n7859) );
  INV_X1 U3679 ( .A(n7859), .ZN(n2520) );
  NOR2_X1 U3680 ( .A1(n5183), .A2(n2520), .ZN(n2496) );
  NOR2_X1 U3681 ( .A1(n2522), .A2(n2496), .ZN(n2525) );
  INV_X1 U3682 ( .A(pmp_addr_i[434]), .ZN(n2498) );
  NAND2_X1 U3683 ( .A1(n2632), .A2(pmp_addr_i[466]), .ZN(n2497) );
  OAI21_X1 U3684 ( .B1(n23), .B2(n2498), .A(n2497), .ZN(n7863) );
  INV_X1 U3685 ( .A(n7863), .ZN(n3291) );
  OR2_X1 U3686 ( .A1(n4802), .A2(n3291), .ZN(n2516) );
  INV_X1 U3687 ( .A(pmp_addr_i[433]), .ZN(n2500) );
  NAND2_X1 U3688 ( .A1(n2632), .A2(pmp_addr_i[465]), .ZN(n2499) );
  OAI21_X1 U3689 ( .B1(n23), .B2(n2500), .A(n2499), .ZN(n7862) );
  NAND2_X1 U3690 ( .A1(n12208), .A2(n7862), .ZN(n2501) );
  NAND4_X1 U3691 ( .A1(n2526), .A2(n2525), .A3(n2516), .A4(n2501), .ZN(n2514)
         );
  INV_X1 U3692 ( .A(pmp_addr_i[444]), .ZN(n2503) );
  NAND2_X1 U3693 ( .A1(n2632), .A2(pmp_addr_i[476]), .ZN(n2502) );
  OAI21_X1 U3694 ( .B1(n23), .B2(n2503), .A(n2502), .ZN(n7871) );
  INV_X1 U3695 ( .A(n7871), .ZN(n2550) );
  NOR2_X1 U3696 ( .A1(n4753), .A2(n2550), .ZN(n2553) );
  INV_X1 U3697 ( .A(pmp_addr_i[443]), .ZN(n2505) );
  NAND2_X1 U3698 ( .A1(n2632), .A2(pmp_addr_i[475]), .ZN(n2504) );
  OAI21_X1 U3699 ( .B1(n23), .B2(n2505), .A(n2504), .ZN(n7870) );
  INV_X1 U3700 ( .A(n7870), .ZN(n2548) );
  NOR2_X1 U3701 ( .A1(n5149), .A2(n2548), .ZN(n2506) );
  NOR2_X1 U3702 ( .A1(n2553), .A2(n2506), .ZN(n2556) );
  INV_X1 U3703 ( .A(pmp_addr_i[445]), .ZN(n2507) );
  NAND2_X1 U3704 ( .A1(n2632), .A2(pmp_addr_i[477]), .ZN(n11145) );
  OAI21_X1 U3705 ( .B1(n23), .B2(n2507), .A(n11145), .ZN(n7874) );
  INV_X1 U3706 ( .A(n7874), .ZN(n2549) );
  NOR2_X1 U3707 ( .A1(pmp_addr_i[446]), .A2(pmp_addr_i[447]), .ZN(n9764) );
  OAI21_X1 U3708 ( .B1(n4866), .B2(n2549), .A(n9764), .ZN(n2557) );
  INV_X1 U3709 ( .A(n2557), .ZN(n2513) );
  INV_X1 U3710 ( .A(pmp_addr_i[441]), .ZN(n2509) );
  NAND2_X1 U3711 ( .A1(n2632), .A2(pmp_addr_i[473]), .ZN(n2508) );
  OAI21_X1 U3712 ( .B1(n23), .B2(n2509), .A(n2508), .ZN(n7867) );
  NAND2_X1 U3713 ( .A1(n5094), .A2(n7867), .ZN(n2512) );
  INV_X1 U3714 ( .A(pmp_addr_i[442]), .ZN(n2511) );
  NAND2_X1 U3715 ( .A1(n2632), .A2(pmp_addr_i[474]), .ZN(n2510) );
  OAI21_X1 U3716 ( .B1(n23), .B2(n2511), .A(n2510), .ZN(n7868) );
  OR2_X1 U3717 ( .A1(n138), .A2(n7901), .ZN(n2544) );
  NAND4_X1 U3718 ( .A1(n2556), .A2(n2513), .A3(n2512), .A4(n2544), .ZN(n2541)
         );
  NOR2_X1 U3719 ( .A1(n2514), .A2(n2541), .ZN(n2515) );
  INV_X1 U3720 ( .A(n2516), .ZN(n2519) );
  INV_X1 U3721 ( .A(n7862), .ZN(n2517) );
  NAND2_X1 U3722 ( .A1(instr_addr_o_19_), .A2(n2517), .ZN(n2518) );
  OAI22_X1 U3723 ( .A1(n2519), .A2(n2518), .B1(n2569), .B2(n7863), .ZN(n2524)
         );
  NAND2_X1 U3724 ( .A1(n5191), .A2(n2520), .ZN(n2521) );
  OAI22_X1 U3725 ( .A1(n2522), .A2(n2521), .B1(n999), .B2(n7860), .ZN(n2523)
         );
  AOI21_X1 U3726 ( .B1(n2525), .B2(n2524), .A(n2523), .ZN(n2540) );
  INV_X1 U3727 ( .A(n2526), .ZN(n2539) );
  INV_X1 U3728 ( .A(n2527), .ZN(n2537) );
  INV_X1 U3729 ( .A(n2528), .ZN(n2531) );
  NAND2_X1 U3730 ( .A1(instr_addr_o_23_), .A2(n2529), .ZN(n2530) );
  OAI22_X1 U3731 ( .A1(n2531), .A2(n2530), .B1(n2580), .B2(n7853), .ZN(n2536)
         );
  NAND2_X1 U3732 ( .A1(n5365), .A2(n2532), .ZN(n2533) );
  OAI22_X1 U3733 ( .A1(n2534), .A2(n2533), .B1(n1273), .B2(n7856), .ZN(n2535)
         );
  AOI21_X1 U3734 ( .B1(n2537), .B2(n2536), .A(n2535), .ZN(n2538) );
  OAI21_X1 U3735 ( .B1(n2540), .B2(n2539), .A(n2538), .ZN(n2543) );
  INV_X1 U3736 ( .A(n2541), .ZN(n2542) );
  NAND2_X1 U3737 ( .A1(n2543), .A2(n2542), .ZN(n2560) );
  INV_X1 U3738 ( .A(n2544), .ZN(n2547) );
  INV_X1 U3739 ( .A(n7867), .ZN(n2545) );
  NAND2_X1 U3740 ( .A1(instr_addr_o_27_), .A2(n2545), .ZN(n2546) );
  OAI22_X1 U3741 ( .A1(n2547), .A2(n2546), .B1(n4438), .B2(n7868), .ZN(n2555)
         );
  NAND2_X1 U3742 ( .A1(instr_addr_o_29_), .A2(n2548), .ZN(n2552) );
  AOI22_X1 U3743 ( .A1(n12199), .A2(n2550), .B1(n4866), .B2(n2549), .ZN(n2551)
         );
  OAI21_X1 U3744 ( .B1(n2553), .B2(n2552), .A(n2551), .ZN(n2554) );
  AOI21_X1 U3745 ( .B1(n2556), .B2(n2555), .A(n2554), .ZN(n2558) );
  INV_X1 U3746 ( .A(pmp_addr_i[476]), .ZN(n2562) );
  NAND2_X1 U3747 ( .A1(n12161), .A2(n2562), .ZN(n2599) );
  OAI21_X1 U3748 ( .B1(n4656), .B2(pmp_addr_i[475]), .A(n2599), .ZN(n2601) );
  INV_X1 U3749 ( .A(pmp_addr_i[474]), .ZN(n2563) );
  INV_X1 U3751 ( .A(pmp_addr_i[477]), .ZN(n2590) );
  NAND2_X1 U3752 ( .A1(n5136), .A2(n2590), .ZN(n2603) );
  NOR2_X1 U3754 ( .A1(n2601), .A2(n2564), .ZN(n2593) );
  INV_X1 U3755 ( .A(instr_addr_i[25]), .ZN(n3992) );
  INV_X1 U3756 ( .A(pmp_addr_i[472]), .ZN(n2565) );
  NAND2_X1 U3757 ( .A1(n12158), .A2(n2565), .ZN(n2585) );
  OAI21_X1 U3758 ( .B1(n135), .B2(pmp_addr_i[471]), .A(n2585), .ZN(n2588) );
  INV_X1 U3759 ( .A(n2588), .ZN(n2568) );
  INV_X1 U3760 ( .A(pmp_addr_i[470]), .ZN(n2566) );
  NAND2_X1 U3761 ( .A1(n5330), .A2(n2566), .ZN(n2582) );
  INV_X1 U3762 ( .A(pmp_addr_i[469]), .ZN(n2579) );
  NAND2_X1 U3763 ( .A1(n5208), .A2(n2579), .ZN(n2567) );
  NAND4_X1 U3764 ( .A1(n2593), .A2(n2568), .A3(n2582), .A4(n2567), .ZN(n2671)
         );
  INV_X1 U3765 ( .A(pmp_addr_i[465]), .ZN(n2665) );
  NOR2_X1 U3766 ( .A1(n5100), .A2(n2665), .ZN(n2570) );
  NAND2_X1 U3767 ( .A1(n6027), .A2(n3980), .ZN(n2667) );
  AOI22_X1 U3768 ( .A1(n2570), .A2(n2667), .B1(n1996), .B2(pmp_addr_i[466]), 
        .ZN(n2577) );
  INV_X1 U3769 ( .A(pmp_addr_i[468]), .ZN(n2571) );
  NAND2_X1 U3770 ( .A1(n4836), .A2(n2571), .ZN(n2574) );
  INV_X1 U3771 ( .A(pmp_addr_i[467]), .ZN(n2573) );
  NAND2_X1 U3772 ( .A1(n4533), .A2(n2573), .ZN(n2572) );
  NAND2_X1 U3773 ( .A1(n2574), .A2(n2572), .ZN(n2664) );
  NOR2_X1 U3774 ( .A1(n5191), .A2(n2573), .ZN(n2575) );
  AOI22_X1 U3775 ( .A1(n2575), .A2(n2574), .B1(n5192), .B2(pmp_addr_i[468]), 
        .ZN(n2576) );
  OAI21_X1 U3776 ( .B1(n2577), .B2(n2664), .A(n2576), .ZN(n2578) );
  INV_X1 U3777 ( .A(n2578), .ZN(n2607) );
  NOR2_X1 U3778 ( .A1(n5208), .A2(n2579), .ZN(n2581) );
  AOI22_X1 U3779 ( .A1(n2582), .A2(n2581), .B1(n2580), .B2(pmp_addr_i[470]), 
        .ZN(n2587) );
  INV_X1 U3780 ( .A(pmp_addr_i[471]), .ZN(n2583) );
  NOR2_X1 U3781 ( .A1(n5202), .A2(n2583), .ZN(n2584) );
  AOI22_X1 U3782 ( .A1(n2585), .A2(n2584), .B1(n3806), .B2(pmp_addr_i[472]), 
        .ZN(n2586) );
  OAI21_X1 U3783 ( .B1(n2588), .B2(n2587), .A(n2586), .ZN(n2592) );
  NOR2_X1 U3784 ( .A1(pmp_addr_i[478]), .A2(pmp_addr_i[479]), .ZN(n2589) );
  OAI21_X1 U3785 ( .B1(n6018), .B2(n2590), .A(n2589), .ZN(n2591) );
  AOI21_X1 U3786 ( .B1(n2593), .B2(n2592), .A(n2591), .ZN(n2606) );
  INV_X1 U3787 ( .A(pmp_addr_i[473]), .ZN(n2594) );
  NOR2_X1 U3788 ( .A1(n5162), .A2(n2594), .ZN(n2595) );
  AOI22_X1 U3789 ( .A1(n2596), .A2(n2595), .B1(n4438), .B2(pmp_addr_i[474]), 
        .ZN(n2602) );
  INV_X1 U3790 ( .A(pmp_addr_i[475]), .ZN(n2597) );
  NOR2_X1 U3791 ( .A1(instr_addr_o_29_), .A2(n2597), .ZN(n2598) );
  AOI22_X1 U3792 ( .A1(n2599), .A2(n2598), .B1(n5115), .B2(pmp_addr_i[476]), 
        .ZN(n2600) );
  OAI21_X1 U3793 ( .B1(n2602), .B2(n2601), .A(n2600), .ZN(n2604) );
  NAND2_X1 U3794 ( .A1(n2604), .A2(n2603), .ZN(n2605) );
  OAI211_X1 U3795 ( .C1(n2671), .C2(n2607), .A(n2606), .B(n2605), .ZN(n2675)
         );
  INV_X1 U3796 ( .A(pmp_cfg_i[114]), .ZN(n2608) );
  NOR2_X1 U3797 ( .A1(n23), .A2(n2608), .ZN(n2674) );
  INV_X1 U3798 ( .A(pmp_addr_i[452]), .ZN(n2609) );
  NAND2_X1 U3799 ( .A1(instr_addr_o_6_), .A2(n2609), .ZN(n2617) );
  INV_X1 U3800 ( .A(pmp_addr_i[451]), .ZN(n2610) );
  NOR2_X1 U3801 ( .A1(n5280), .A2(n2610), .ZN(n2612) );
  AOI22_X1 U3802 ( .A1(n2617), .A2(n2612), .B1(n2611), .B2(pmp_addr_i[452]), 
        .ZN(n2621) );
  OR2_X1 U3803 ( .A1(pmp_addr_i[449]), .A2(pmp_addr_i[448]), .ZN(n2613) );
  NOR2_X1 U3804 ( .A1(n2613), .A2(pmp_addr_i[450]), .ZN(n2615) );
  INV_X1 U3805 ( .A(n2613), .ZN(n2614) );
  OAI22_X1 U3806 ( .A1(n5899), .A2(n2615), .B1(n2614), .B2(n2391), .ZN(n2616)
         );
  OAI211_X1 U3807 ( .C1(pmp_addr_i[451]), .C2(n3839), .A(n2617), .B(n2616), 
        .ZN(n2620) );
  NAND2_X1 U3808 ( .A1(n154), .A2(n3906), .ZN(n2627) );
  NAND2_X1 U3809 ( .A1(n205), .A2(n2400), .ZN(n2625) );
  NAND2_X1 U3810 ( .A1(n5270), .A2(n3903), .ZN(n2626) );
  INV_X1 U3811 ( .A(pmp_addr_i[453]), .ZN(n2624) );
  NAND2_X1 U3812 ( .A1(n5268), .A2(n2624), .ZN(n2618) );
  NAND4_X1 U3813 ( .A1(n2627), .A2(n2625), .A3(n2626), .A4(n2618), .ZN(n2619)
         );
  AOI21_X1 U3814 ( .B1(n2621), .B2(n2620), .A(n2619), .ZN(n2639) );
  NOR2_X1 U3815 ( .A1(n5040), .A2(n3906), .ZN(n2622) );
  AOI22_X1 U3816 ( .A1(n2622), .A2(n2626), .B1(n4602), .B2(pmp_addr_i[456]), 
        .ZN(n2630) );
  OAI22_X1 U3817 ( .A1(n5740), .A2(n2624), .B1(n6005), .B2(n2400), .ZN(n2628)
         );
  NAND4_X1 U3818 ( .A1(n2628), .A2(n2627), .A3(n2626), .A4(n2625), .ZN(n2629)
         );
  NAND2_X1 U3819 ( .A1(n2630), .A2(n2629), .ZN(n2638) );
  NAND2_X1 U3820 ( .A1(n5251), .A2(n3926), .ZN(n2652) );
  INV_X1 U3821 ( .A(pmp_addr_i[459]), .ZN(n2650) );
  NAND2_X1 U3822 ( .A1(n4061), .A2(n2650), .ZN(n2631) );
  NAND2_X1 U3823 ( .A1(n2652), .A2(n2631), .ZN(n2654) );
  OR2_X1 U3824 ( .A1(n2632), .A2(n7923), .ZN(n7927) );
  AND2_X1 U3825 ( .A1(n7927), .A2(pmp_addr_i[462]), .ZN(n7715) );
  INV_X1 U3826 ( .A(n7715), .ZN(n2633) );
  NAND2_X1 U3827 ( .A1(n5229), .A2(n2633), .ZN(n2658) );
  INV_X1 U3828 ( .A(pmp_addr_i[458]), .ZN(n2634) );
  NAND2_X1 U3829 ( .A1(n5245), .A2(n2634), .ZN(n2649) );
  INV_X1 U3830 ( .A(pmp_addr_i[463]), .ZN(n2641) );
  NAND2_X1 U3831 ( .A1(n12265), .A2(n2641), .ZN(n2640) );
  NAND2_X1 U3832 ( .A1(instr_addr_o_11_), .A2(n3933), .ZN(n2635) );
  NAND2_X1 U3833 ( .A1(instr_addr_o_15_), .A2(n3226), .ZN(n2656) );
  INV_X1 U3834 ( .A(pmp_addr_i[464]), .ZN(n2636) );
  NAND2_X1 U3835 ( .A1(n5047), .A2(n2636), .ZN(n2643) );
  NAND2_X1 U3836 ( .A1(n2656), .A2(n2643), .ZN(n2637) );
  AND2_X1 U3837 ( .A1(n2643), .A2(n2640), .ZN(n2659) );
  INV_X1 U3838 ( .A(n2659), .ZN(n2646) );
  NAND2_X1 U3839 ( .A1(n12217), .A2(n7715), .ZN(n2645) );
  NOR2_X1 U3840 ( .A1(n12156), .A2(n2641), .ZN(n2642) );
  AOI22_X1 U3841 ( .A1(n2643), .A2(n2642), .B1(n1922), .B2(pmp_addr_i[464]), 
        .ZN(n2644) );
  OAI21_X1 U3842 ( .B1(n2646), .B2(n2645), .A(n2644), .ZN(n2647) );
  INV_X1 U3843 ( .A(n2647), .ZN(n2662) );
  NOR2_X1 U3844 ( .A1(n3934), .A2(n3933), .ZN(n2648) );
  AOI22_X1 U3845 ( .A1(n2649), .A2(n2648), .B1(n5070), .B2(pmp_addr_i[458]), 
        .ZN(n2655) );
  NOR2_X1 U3846 ( .A1(n150), .A2(n2650), .ZN(n2651) );
  AOI22_X1 U3847 ( .A1(n2652), .A2(n2651), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[460]), .ZN(n2653) );
  OAI21_X1 U3848 ( .B1(n2655), .B2(n2654), .A(n2653), .ZN(n2657) );
  NAND4_X1 U3849 ( .A1(n2657), .A2(n2659), .A3(n2658), .A4(n2656), .ZN(n2661)
         );
  NAND4_X1 U3850 ( .A1(n2659), .A2(pmp_addr_i[461]), .A3(n6017), .A4(n2658), 
        .ZN(n2660) );
  NAND4_X1 U3851 ( .A1(n2663), .A2(n2662), .A3(n2661), .A4(n2660), .ZN(n2673)
         );
  INV_X1 U3852 ( .A(n2664), .ZN(n2669) );
  NAND2_X1 U3853 ( .A1(instr_addr_o_19_), .A2(n2665), .ZN(n2666) );
  AND2_X1 U3854 ( .A1(n2667), .A2(n2666), .ZN(n2668) );
  NAND3_X1 U3855 ( .A1(n2669), .A2(n2674), .A3(n2668), .ZN(n2670) );
  NOR2_X1 U3856 ( .A1(n2671), .A2(n2670), .ZN(n2672) );
  AOI22_X1 U3857 ( .A1(n2675), .A2(n2674), .B1(n2673), .B2(n2672), .ZN(n2930)
         );
  NAND2_X1 U3858 ( .A1(pmp_addr_i[33]), .A2(pmp_addr_i[32]), .ZN(n4995) );
  OR2_X1 U3859 ( .A1(n4995), .A2(n2683), .ZN(n11487) );
  INV_X1 U3860 ( .A(pmp_cfg_i[11]), .ZN(n2695) );
  OAI21_X1 U3861 ( .B1(n11487), .B2(n2695), .A(pmp_cfg_i[12]), .ZN(n2684) );
  NAND2_X1 U3862 ( .A1(n2693), .A2(pmp_cfg_i[12]), .ZN(n2677) );
  INV_X1 U3863 ( .A(pmp_addr_i[36]), .ZN(n2676) );
  AOI21_X1 U3864 ( .B1(n2684), .B2(n2677), .A(n2676), .ZN(n2679) );
  AND2_X1 U3865 ( .A1(n36), .A2(pmp_addr_i[4]), .ZN(n2678) );
  NAND2_X1 U3866 ( .A1(n36), .A2(pmp_addr_i[3]), .ZN(n2681) );
  OAI21_X1 U3867 ( .B1(n2684), .B2(n2693), .A(n2681), .ZN(n8222) );
  INV_X1 U3868 ( .A(n8222), .ZN(n8379) );
  NOR2_X1 U3869 ( .A1(n20), .A2(n8379), .ZN(n4970) );
  NAND2_X1 U3870 ( .A1(n36), .A2(pmp_addr_i[2]), .ZN(n2682) );
  OAI21_X1 U3871 ( .B1(n2684), .B2(n2683), .A(n2682), .ZN(n8219) );
  AND2_X1 U3872 ( .A1(pmp_cfg_i[11]), .A2(pmp_addr_i[32]), .ZN(n2687) );
  NAND2_X1 U3873 ( .A1(pmp_cfg_i[12]), .A2(pmp_addr_i[33]), .ZN(n2686) );
  NAND2_X1 U3874 ( .A1(n36), .A2(pmp_addr_i[1]), .ZN(n2685) );
  OAI21_X1 U3875 ( .B1(n2687), .B2(n2686), .A(n2685), .ZN(n8380) );
  NAND2_X1 U3876 ( .A1(n36), .A2(pmp_addr_i[0]), .ZN(n2689) );
  OR2_X1 U3877 ( .A1(n11482), .A2(pmp_cfg_i[11]), .ZN(n2688) );
  NAND2_X1 U3878 ( .A1(n2689), .A2(n2688), .ZN(n8381) );
  OR2_X1 U3879 ( .A1(n8380), .A2(n8381), .ZN(n2690) );
  NAND2_X1 U3880 ( .A1(n8219), .A2(n2690), .ZN(n2691) );
  INV_X1 U3881 ( .A(n8219), .ZN(n8334) );
  INV_X1 U3882 ( .A(n2690), .ZN(n4997) );
  AOI22_X1 U3883 ( .A1(n3836), .A2(n2691), .B1(n8334), .B2(n4997), .ZN(n2692)
         );
  NOR3_X1 U3884 ( .A1(n4958), .A2(n4970), .A3(n2692), .ZN(n2706) );
  NAND2_X1 U3885 ( .A1(instr_addr_o_5_), .A2(n8379), .ZN(n4993) );
  NAND2_X1 U3886 ( .A1(instr_addr_o_6_), .A2(n327), .ZN(n4932) );
  OAI21_X1 U3887 ( .B1(n4958), .B2(n4993), .A(n4932), .ZN(n2705) );
  NAND2_X1 U3888 ( .A1(n11476), .A2(pmp_addr_i[36]), .ZN(n11479) );
  INV_X1 U3889 ( .A(pmp_addr_i[37]), .ZN(n2694) );
  OR2_X1 U3890 ( .A1(n11479), .A2(n2694), .ZN(n11512) );
  OR2_X1 U3891 ( .A1(n11512), .A2(n2695), .ZN(n2734) );
  NAND2_X1 U3892 ( .A1(pmp_addr_i[39]), .A2(pmp_addr_i[38]), .ZN(n11493) );
  OAI21_X1 U3893 ( .B1(n2734), .B2(n11493), .A(pmp_cfg_i[12]), .ZN(n2730) );
  NAND2_X1 U3894 ( .A1(n36), .A2(pmp_addr_i[7]), .ZN(n2696) );
  OAI21_X1 U3895 ( .B1(n2730), .B2(n2697), .A(n2696), .ZN(n8236) );
  INV_X1 U3896 ( .A(n8236), .ZN(n8228) );
  NOR2_X1 U3897 ( .A1(n155), .A2(n8228), .ZN(n4949) );
  NAND2_X1 U3898 ( .A1(n36), .A2(pmp_addr_i[8]), .ZN(n2698) );
  OAI21_X1 U3899 ( .B1(n2730), .B2(n4937), .A(n2698), .ZN(n8235) );
  INV_X1 U3900 ( .A(n8235), .ZN(n8229) );
  INV_X1 U3901 ( .A(pmp_addr_i[5]), .ZN(n2701) );
  AND2_X1 U3902 ( .A1(pmp_cfg_i[12]), .A2(pmp_addr_i[37]), .ZN(n2699) );
  NAND2_X1 U3903 ( .A1(n2734), .A2(n2699), .ZN(n2700) );
  OAI21_X1 U3904 ( .B1(n160), .B2(n2701), .A(n2700), .ZN(n8231) );
  INV_X1 U3905 ( .A(n8231), .ZN(n4989) );
  NOR2_X1 U3906 ( .A1(n4605), .A2(n4989), .ZN(n4928) );
  INV_X1 U3907 ( .A(pmp_addr_i[6]), .ZN(n3655) );
  AND2_X1 U3908 ( .A1(pmp_cfg_i[12]), .A2(pmp_addr_i[38]), .ZN(n2702) );
  NAND2_X1 U3909 ( .A1(n2734), .A2(n2702), .ZN(n2703) );
  OAI21_X1 U3910 ( .B1(n160), .B2(n3655), .A(n2703), .ZN(n8230) );
  INV_X1 U3911 ( .A(n8230), .ZN(n8339) );
  NOR2_X1 U3912 ( .A1(n5342), .A2(n8339), .ZN(n4941) );
  NOR2_X1 U3913 ( .A1(n4928), .A2(n4941), .ZN(n2704) );
  OAI211_X1 U3914 ( .C1(n2706), .C2(n2705), .A(n2704), .B(n2711), .ZN(n2713)
         );
  NAND2_X1 U3915 ( .A1(n5268), .A2(n4989), .ZN(n2708) );
  OAI22_X1 U3916 ( .A1(n4941), .A2(n2708), .B1(n4606), .B2(n8230), .ZN(n2710)
         );
  NAND2_X1 U3917 ( .A1(n5040), .A2(n8228), .ZN(n4920) );
  NAND2_X1 U3918 ( .A1(n5270), .A2(n8229), .ZN(n4921) );
  OAI21_X1 U3919 ( .B1(n4920), .B2(n4965), .A(n4921), .ZN(n2709) );
  AOI21_X1 U3920 ( .B1(n2711), .B2(n2710), .A(n2709), .ZN(n2712) );
  NAND3_X1 U3921 ( .A1(pmp_addr_i[40]), .A2(pmp_addr_i[42]), .A3(
        pmp_addr_i[41]), .ZN(n2714) );
  OR2_X1 U3922 ( .A1(n11493), .A2(n2714), .ZN(n4933) );
  NAND2_X1 U3923 ( .A1(pmp_addr_i[44]), .A2(pmp_addr_i[43]), .ZN(n4967) );
  NOR2_X1 U3924 ( .A1(n4933), .A2(n4967), .ZN(n2722) );
  NAND2_X1 U3925 ( .A1(n2722), .A2(pmp_addr_i[45]), .ZN(n2715) );
  NOR2_X1 U3926 ( .A1(n11512), .A2(n2715), .ZN(n11473) );
  NAND2_X1 U3927 ( .A1(n11473), .A2(pmp_addr_i[46]), .ZN(n11510) );
  NAND2_X1 U3928 ( .A1(pmp_cfg_i[11]), .A2(pmp_addr_i[47]), .ZN(n2716) );
  INV_X1 U3929 ( .A(pmp_addr_i[48]), .ZN(n2718) );
  NAND2_X1 U3930 ( .A1(n36), .A2(pmp_addr_i[16]), .ZN(n2717) );
  OAI21_X1 U3931 ( .B1(n4996), .B2(n2718), .A(n2717), .ZN(n8366) );
  INV_X1 U3932 ( .A(n8366), .ZN(n2719) );
  NOR2_X1 U3933 ( .A1(n6019), .A2(n2719), .ZN(n2752) );
  INV_X1 U3934 ( .A(pmp_addr_i[47]), .ZN(n2721) );
  NAND2_X1 U3935 ( .A1(n36), .A2(pmp_addr_i[15]), .ZN(n2720) );
  OAI21_X1 U3936 ( .B1(n4996), .B2(n2721), .A(n2720), .ZN(n8254) );
  INV_X1 U3937 ( .A(n8254), .ZN(n5000) );
  OR2_X1 U3938 ( .A1(n2752), .A2(n4966), .ZN(n2749) );
  INV_X1 U3939 ( .A(n2722), .ZN(n11469) );
  OAI21_X1 U3940 ( .B1(n2734), .B2(n11469), .A(pmp_cfg_i[12]), .ZN(n2741) );
  NAND2_X1 U3941 ( .A1(n36), .A2(pmp_addr_i[13]), .ZN(n2723) );
  OAI21_X1 U3942 ( .B1(n2741), .B2(n2724), .A(n2723), .ZN(n8204) );
  INV_X1 U3943 ( .A(n8204), .ZN(n8326) );
  NOR2_X1 U3944 ( .A1(n208), .A2(n8326), .ZN(n4948) );
  NAND2_X1 U3945 ( .A1(n2724), .A2(pmp_cfg_i[12]), .ZN(n2725) );
  AOI21_X1 U3946 ( .B1(n2741), .B2(n2725), .A(n2891), .ZN(n2727) );
  AND2_X1 U3947 ( .A1(n36), .A2(pmp_addr_i[14]), .ZN(n2726) );
  NOR2_X1 U3948 ( .A1(n3100), .A2(n325), .ZN(n4976) );
  OR2_X1 U3949 ( .A1(n4948), .A2(n4976), .ZN(n2728) );
  NOR2_X1 U3950 ( .A1(n2749), .A2(n2728), .ZN(n2747) );
  NAND2_X1 U3951 ( .A1(n4937), .A2(pmp_cfg_i[12]), .ZN(n2729) );
  AOI21_X1 U3952 ( .B1(n2730), .B2(n2729), .A(n4981), .ZN(n2732) );
  AND2_X1 U3953 ( .A1(n36), .A2(pmp_addr_i[9]), .ZN(n2731) );
  NOR2_X1 U3954 ( .A1(n6002), .A2(n326), .ZN(n4940) );
  INV_X1 U3955 ( .A(n2733), .ZN(n4494) );
  OAI21_X1 U3956 ( .B1(n2734), .B2(n4933), .A(pmp_cfg_i[12]), .ZN(n2738) );
  INV_X1 U3957 ( .A(pmp_addr_i[42]), .ZN(n2736) );
  NAND2_X1 U3958 ( .A1(n36), .A2(pmp_addr_i[10]), .ZN(n2735) );
  OAI21_X1 U3959 ( .B1(n2738), .B2(n2736), .A(n2735), .ZN(n8208) );
  INV_X1 U3960 ( .A(n8208), .ZN(n8341) );
  NOR2_X1 U3961 ( .A1(n4940), .A2(n2743), .ZN(n2742) );
  INV_X1 U3962 ( .A(pmp_addr_i[43]), .ZN(n4934) );
  NAND2_X1 U3963 ( .A1(n36), .A2(pmp_addr_i[11]), .ZN(n2737) );
  OAI21_X1 U3964 ( .B1(n2738), .B2(n4934), .A(n2737), .ZN(n8210) );
  INV_X1 U3965 ( .A(n8210), .ZN(n8340) );
  NOR2_X1 U3966 ( .A1(n5997), .A2(n8340), .ZN(n4957) );
  NAND2_X1 U3968 ( .A1(n36), .A2(pmp_addr_i[12]), .ZN(n2740) );
  OAI21_X1 U3969 ( .B1(n2741), .B2(n2889), .A(n2740), .ZN(n8211) );
  INV_X1 U3970 ( .A(n8211), .ZN(n8325) );
  NOR2_X1 U3971 ( .A1(n12180), .A2(n8325), .ZN(n4929) );
  NOR2_X1 U3972 ( .A1(n4957), .A2(n4929), .ZN(n2744) );
  AND2_X1 U3973 ( .A1(n6002), .A2(n326), .ZN(n4939) );
  INV_X1 U3974 ( .A(n2743), .ZN(n4977) );
  AND2_X1 U3975 ( .A1(n5245), .A2(n8341), .ZN(n4980) );
  AOI21_X1 U3976 ( .B1(n4939), .B2(n4977), .A(n4980), .ZN(n2746) );
  INV_X1 U3977 ( .A(n2744), .ZN(n2745) );
  NAND2_X1 U3978 ( .A1(instr_addr_o_13_), .A2(n8340), .ZN(n4955) );
  NAND2_X1 U3979 ( .A1(n5251), .A2(n8325), .ZN(n4936) );
  OAI21_X1 U3980 ( .B1(n4929), .B2(n4955), .A(n4936), .ZN(n2748) );
  INV_X1 U3981 ( .A(n2749), .ZN(n2755) );
  NAND2_X1 U3982 ( .A1(instr_addr_o_15_), .A2(n8326), .ZN(n4956) );
  NAND2_X1 U3983 ( .A1(n12203), .A2(n325), .ZN(n4979) );
  OAI21_X1 U3984 ( .B1(n4976), .B2(n4956), .A(n4979), .ZN(n2754) );
  NAND2_X1 U3985 ( .A1(n12265), .A2(n5000), .ZN(n2751) );
  BUF_X1 U3986 ( .A(n3000), .Z(n2750) );
  OAI22_X1 U3987 ( .A1(n2752), .A2(n2751), .B1(n2750), .B2(n8366), .ZN(n2753)
         );
  AOI21_X1 U3988 ( .B1(n2755), .B2(n2754), .A(n2753), .ZN(n2756) );
  INV_X1 U3989 ( .A(pmp_addr_i[29]), .ZN(n2759) );
  OR2_X1 U3990 ( .A1(n4996), .A2(n2758), .ZN(n12075) );
  OAI21_X1 U3991 ( .B1(n160), .B2(n2759), .A(n12075), .ZN(n8276) );
  INV_X1 U3992 ( .A(n8276), .ZN(n8385) );
  INV_X1 U3993 ( .A(pmp_addr_i[31]), .ZN(n2760) );
  NOR2_X1 U3994 ( .A1(pmp_addr_i[30]), .A2(pmp_addr_i[31]), .ZN(n2761) );
  OAI21_X1 U3995 ( .B1(n6018), .B2(n8385), .A(n2761), .ZN(n2837) );
  INV_X1 U3996 ( .A(n2837), .ZN(n2771) );
  NAND2_X1 U3997 ( .A1(n36), .A2(pmp_addr_i[28]), .ZN(n2762) );
  OAI21_X1 U3998 ( .B1(n4996), .B2(n2839), .A(n2762), .ZN(n8361) );
  INV_X1 U3999 ( .A(n8361), .ZN(n2830) );
  NOR2_X1 U4000 ( .A1(n4560), .A2(n2830), .ZN(n2833) );
  INV_X1 U4001 ( .A(pmp_addr_i[59]), .ZN(n2764) );
  NAND2_X1 U4002 ( .A1(n36), .A2(pmp_addr_i[27]), .ZN(n2763) );
  OAI21_X1 U4003 ( .B1(n4996), .B2(n2764), .A(n2763), .ZN(n8330) );
  INV_X1 U4004 ( .A(n8330), .ZN(n2829) );
  NOR2_X1 U4005 ( .A1(n5149), .A2(n2829), .ZN(n2765) );
  NOR2_X1 U4006 ( .A1(n2833), .A2(n2765), .ZN(n2836) );
  INV_X1 U4007 ( .A(pmp_addr_i[58]), .ZN(n2767) );
  NAND2_X1 U4008 ( .A1(n36), .A2(pmp_addr_i[26]), .ZN(n2766) );
  OAI21_X1 U4009 ( .B1(n4996), .B2(n2767), .A(n2766), .ZN(n8360) );
  OR2_X1 U4010 ( .A1(n5368), .A2(n8302), .ZN(n2825) );
  INV_X1 U4011 ( .A(pmp_addr_i[57]), .ZN(n2769) );
  NAND2_X1 U4012 ( .A1(n36), .A2(pmp_addr_i[25]), .ZN(n2768) );
  OAI21_X1 U4013 ( .B1(n4996), .B2(n2769), .A(n2768), .ZN(n8369) );
  NAND2_X1 U4014 ( .A1(n5094), .A2(n8369), .ZN(n2770) );
  NAND4_X1 U4015 ( .A1(n2771), .A2(n2836), .A3(n2825), .A4(n2770), .ZN(n2822)
         );
  INV_X1 U4016 ( .A(pmp_addr_i[49]), .ZN(n2773) );
  NAND2_X1 U4017 ( .A1(n36), .A2(pmp_addr_i[17]), .ZN(n2772) );
  OAI21_X1 U4018 ( .B1(n4996), .B2(n2773), .A(n2772), .ZN(n8348) );
  NAND2_X1 U4019 ( .A1(n12208), .A2(n8348), .ZN(n2783) );
  INV_X1 U4020 ( .A(pmp_addr_i[50]), .ZN(n2775) );
  NAND2_X1 U4021 ( .A1(n36), .A2(pmp_addr_i[18]), .ZN(n2774) );
  OAI21_X1 U4022 ( .B1(n4996), .B2(n2775), .A(n2774), .ZN(n8349) );
  INV_X1 U4023 ( .A(n8349), .ZN(n2776) );
  INV_X1 U4024 ( .A(pmp_addr_i[52]), .ZN(n2778) );
  NAND2_X1 U4025 ( .A1(n36), .A2(pmp_addr_i[20]), .ZN(n2777) );
  OAI21_X1 U4026 ( .B1(n4996), .B2(n2778), .A(n2777), .ZN(n8350) );
  INV_X1 U4027 ( .A(n8350), .ZN(n2779) );
  NOR2_X1 U4028 ( .A1(n4836), .A2(n2779), .ZN(n2803) );
  INV_X1 U4029 ( .A(pmp_addr_i[51]), .ZN(n2781) );
  NAND2_X1 U4030 ( .A1(n36), .A2(pmp_addr_i[19]), .ZN(n2780) );
  OAI21_X1 U4031 ( .B1(n4996), .B2(n2781), .A(n2780), .ZN(n8367) );
  INV_X1 U4032 ( .A(n8367), .ZN(n2801) );
  NOR2_X1 U4033 ( .A1(n5842), .A2(n2801), .ZN(n2782) );
  NOR2_X1 U4034 ( .A1(n2803), .A2(n2782), .ZN(n2806) );
  NOR2_X1 U4035 ( .A1(n2822), .A2(n2784), .ZN(n2797) );
  INV_X1 U4036 ( .A(pmp_addr_i[56]), .ZN(n2786) );
  NAND2_X1 U4037 ( .A1(n36), .A2(pmp_addr_i[24]), .ZN(n2785) );
  OAI21_X1 U4038 ( .B1(n4996), .B2(n2786), .A(n2785), .ZN(n8359) );
  INV_X1 U4039 ( .A(n8359), .ZN(n2787) );
  NOR2_X1 U4040 ( .A1(n210), .A2(n2787), .ZN(n2815) );
  INV_X1 U4041 ( .A(pmp_addr_i[55]), .ZN(n2789) );
  NAND2_X1 U4042 ( .A1(n36), .A2(pmp_addr_i[23]), .ZN(n2788) );
  OAI21_X1 U4043 ( .B1(n4996), .B2(n2789), .A(n2788), .ZN(n8358) );
  INV_X1 U4044 ( .A(n8358), .ZN(n2813) );
  OR2_X1 U4046 ( .A1(n2815), .A2(n12187), .ZN(n2808) );
  INV_X1 U4047 ( .A(pmp_addr_i[53]), .ZN(n2792) );
  NAND2_X1 U4048 ( .A1(n36), .A2(pmp_addr_i[21]), .ZN(n2791) );
  OAI21_X1 U4049 ( .B1(n4996), .B2(n2792), .A(n2791), .ZN(n8351) );
  INV_X1 U4050 ( .A(n8351), .ZN(n2810) );
  INV_X1 U4051 ( .A(pmp_addr_i[54]), .ZN(n2794) );
  NAND2_X1 U4052 ( .A1(n36), .A2(pmp_addr_i[22]), .ZN(n2793) );
  OAI21_X1 U4053 ( .B1(n4996), .B2(n2794), .A(n2793), .ZN(n8368) );
  INV_X1 U4054 ( .A(n8368), .ZN(n2795) );
  OR2_X1 U4055 ( .A1(n5330), .A2(n2795), .ZN(n2809) );
  OAI21_X1 U4056 ( .B1(n5208), .B2(n2810), .A(n2809), .ZN(n2796) );
  NOR2_X1 U4057 ( .A1(n2808), .A2(n2796), .ZN(n2807) );
  INV_X1 U4058 ( .A(n8348), .ZN(n2798) );
  NAND2_X1 U4059 ( .A1(n3793), .A2(n2798), .ZN(n2799) );
  OAI22_X1 U4060 ( .A1(n2800), .A2(n2799), .B1(n1996), .B2(n8349), .ZN(n2805)
         );
  NAND2_X1 U4061 ( .A1(n5191), .A2(n2801), .ZN(n2802) );
  OAI22_X1 U4062 ( .A1(n2803), .A2(n2802), .B1(n999), .B2(n8350), .ZN(n2804)
         );
  AOI21_X1 U4063 ( .B1(n2806), .B2(n2805), .A(n2804), .ZN(n2821) );
  INV_X1 U4064 ( .A(n2807), .ZN(n2820) );
  INV_X1 U4065 ( .A(n2808), .ZN(n2818) );
  INV_X1 U4066 ( .A(n2809), .ZN(n2812) );
  NAND2_X1 U4067 ( .A1(instr_addr_o_23_), .A2(n2810), .ZN(n2811) );
  OAI22_X1 U4068 ( .A1(n2812), .A2(n2811), .B1(n1269), .B2(n8368), .ZN(n2817)
         );
  NAND2_X1 U4069 ( .A1(n5365), .A2(n2813), .ZN(n2814) );
  OAI22_X1 U4070 ( .A1(n2815), .A2(n2814), .B1(n3806), .B2(n8359), .ZN(n2816)
         );
  AOI21_X1 U4071 ( .B1(n2818), .B2(n2817), .A(n2816), .ZN(n2819) );
  OAI21_X1 U4072 ( .B1(n2821), .B2(n2820), .A(n2819), .ZN(n2824) );
  INV_X1 U4073 ( .A(n2822), .ZN(n2823) );
  INV_X1 U4074 ( .A(n2825), .ZN(n2828) );
  INV_X1 U4075 ( .A(n8369), .ZN(n2826) );
  NAND2_X1 U4076 ( .A1(instr_addr_o_27_), .A2(n2826), .ZN(n2827) );
  OAI22_X1 U4077 ( .A1(n2828), .A2(n2827), .B1(n4438), .B2(n8360), .ZN(n2835)
         );
  NAND2_X1 U4078 ( .A1(n4900), .A2(n2829), .ZN(n2832) );
  AOI22_X1 U4079 ( .A1(n12161), .A2(n2830), .B1(n5154), .B2(n8385), .ZN(n2831)
         );
  OAI21_X1 U4080 ( .B1(n2833), .B2(n2832), .A(n2831), .ZN(n2834) );
  AOI21_X1 U4081 ( .B1(n2836), .B2(n2835), .A(n2834), .ZN(n2838) );
  NAND2_X1 U4082 ( .A1(n4866), .A2(n2758), .ZN(n2866) );
  INV_X1 U4083 ( .A(n1632), .ZN(n12263) );
  INV_X1 U4084 ( .A(pmp_addr_i[60]), .ZN(n2839) );
  NAND2_X1 U4085 ( .A1(n5980), .A2(n2839), .ZN(n2862) );
  OAI21_X1 U4086 ( .B1(n4406), .B2(pmp_addr_i[59]), .A(n2862), .ZN(n2864) );
  NAND2_X1 U4087 ( .A1(n210), .A2(n2786), .ZN(n2852) );
  OAI21_X1 U4088 ( .B1(n135), .B2(pmp_addr_i[55]), .A(n2852), .ZN(n2855) );
  INV_X1 U4089 ( .A(n2855), .ZN(n2841) );
  NAND2_X1 U4090 ( .A1(n4835), .A2(n2794), .ZN(n2850) );
  NAND2_X1 U4091 ( .A1(instr_addr_o_23_), .A2(n2792), .ZN(n2840) );
  NOR2_X1 U4092 ( .A1(n6020), .A2(n2773), .ZN(n2842) );
  NAND2_X1 U4093 ( .A1(n6027), .A2(n2775), .ZN(n2920) );
  AOI22_X1 U4094 ( .A1(n2842), .A2(n2920), .B1(n1996), .B2(pmp_addr_i[50]), 
        .ZN(n2847) );
  NAND2_X1 U4095 ( .A1(n4836), .A2(n2778), .ZN(n2844) );
  NAND2_X1 U4096 ( .A1(n4533), .A2(n2781), .ZN(n2843) );
  NAND2_X1 U4097 ( .A1(n2844), .A2(n2843), .ZN(n2918) );
  NOR2_X1 U4098 ( .A1(n5183), .A2(n2781), .ZN(n2845) );
  AOI22_X1 U4099 ( .A1(n2845), .A2(n2844), .B1(n999), .B2(pmp_addr_i[52]), 
        .ZN(n2846) );
  OAI21_X1 U4100 ( .B1(n2847), .B2(n2918), .A(n2846), .ZN(n2848) );
  INV_X1 U4101 ( .A(n2848), .ZN(n2870) );
  NOR2_X1 U4102 ( .A1(instr_addr_o_23_), .A2(n2792), .ZN(n2849) );
  AOI22_X1 U4103 ( .A1(n2850), .A2(n2849), .B1(n2580), .B2(pmp_addr_i[54]), 
        .ZN(n2854) );
  NOR2_X1 U4104 ( .A1(n12226), .A2(n2789), .ZN(n2851) );
  AOI22_X1 U4105 ( .A1(n2852), .A2(n2851), .B1(n3806), .B2(pmp_addr_i[56]), 
        .ZN(n2853) );
  OAI21_X1 U4106 ( .B1(n2855), .B2(n2854), .A(n2853), .ZN(n2857) );
  NOR2_X1 U4107 ( .A1(pmp_addr_i[62]), .A2(pmp_addr_i[63]), .ZN(n8193) );
  OAI21_X1 U4108 ( .B1(n4866), .B2(n2758), .A(n8193), .ZN(n2856) );
  AOI21_X1 U4109 ( .B1(n2858), .B2(n2857), .A(n2856), .ZN(n2869) );
  NOR2_X1 U4110 ( .A1(n5162), .A2(n2769), .ZN(n2859) );
  AOI22_X1 U4111 ( .A1(n2860), .A2(n2859), .B1(n4438), .B2(pmp_addr_i[58]), 
        .ZN(n2865) );
  NOR2_X1 U4112 ( .A1(n5149), .A2(n2764), .ZN(n2861) );
  AOI22_X1 U4113 ( .A1(n2862), .A2(n2861), .B1(n4658), .B2(pmp_addr_i[60]), 
        .ZN(n2863) );
  OAI21_X1 U4114 ( .B1(n2865), .B2(n2864), .A(n2863), .ZN(n2867) );
  NAND2_X1 U4115 ( .A1(n2867), .A2(n2866), .ZN(n2868) );
  OAI211_X1 U4116 ( .C1(n2924), .C2(n2870), .A(n2869), .B(n2868), .ZN(n2928)
         );
  AND2_X1 U4117 ( .A1(n36), .A2(pmp_cfg_i[10]), .ZN(n2927) );
  NAND2_X1 U4118 ( .A1(instr_addr_o_6_), .A2(n2676), .ZN(n2876) );
  NOR2_X1 U4119 ( .A1(n5280), .A2(n2693), .ZN(n2871) );
  AOI22_X1 U4120 ( .A1(n2876), .A2(n2871), .B1(n2611), .B2(pmp_addr_i[36]), 
        .ZN(n2880) );
  OR2_X1 U4121 ( .A1(pmp_addr_i[33]), .A2(pmp_addr_i[32]), .ZN(n2872) );
  NOR2_X1 U4122 ( .A1(n2872), .A2(pmp_addr_i[34]), .ZN(n2874) );
  INV_X1 U4123 ( .A(n2872), .ZN(n2873) );
  OAI22_X1 U4124 ( .A1(n5899), .A2(n2874), .B1(n2873), .B2(n2683), .ZN(n2875)
         );
  OAI211_X1 U4125 ( .C1(pmp_addr_i[35]), .C2(n3839), .A(n2876), .B(n2875), 
        .ZN(n2879) );
  NAND2_X1 U4126 ( .A1(n154), .A2(n2697), .ZN(n2885) );
  NAND2_X1 U4127 ( .A1(n205), .A2(n1943), .ZN(n2883) );
  NAND2_X1 U4128 ( .A1(n5270), .A2(n4937), .ZN(n2884) );
  NAND2_X1 U4129 ( .A1(n5268), .A2(n2694), .ZN(n2877) );
  NAND4_X1 U4130 ( .A1(n2885), .A2(n2883), .A3(n2884), .A4(n2877), .ZN(n2878)
         );
  AOI21_X1 U4131 ( .B1(n2880), .B2(n2879), .A(n2878), .ZN(n2894) );
  NOR2_X1 U4132 ( .A1(n155), .A2(n2697), .ZN(n2882) );
  AOI22_X1 U4133 ( .A1(n2882), .A2(n2884), .B1(n4602), .B2(pmp_addr_i[40]), 
        .ZN(n2888) );
  OAI22_X1 U4134 ( .A1(n5740), .A2(n2694), .B1(n6005), .B2(n1943), .ZN(n2886)
         );
  NAND4_X1 U4135 ( .A1(n2886), .A2(n2885), .A3(n2884), .A4(n2883), .ZN(n2887)
         );
  NAND2_X1 U4136 ( .A1(n2888), .A2(n2887), .ZN(n2893) );
  INV_X1 U4137 ( .A(pmp_addr_i[44]), .ZN(n2889) );
  NAND2_X1 U4138 ( .A1(n5251), .A2(n2889), .ZN(n2906) );
  NAND2_X1 U4139 ( .A1(n4061), .A2(n4934), .ZN(n2890) );
  NAND2_X1 U4140 ( .A1(n2906), .A2(n2890), .ZN(n2908) );
  INV_X1 U4141 ( .A(pmp_addr_i[46]), .ZN(n2891) );
  NAND2_X1 U4142 ( .A1(n5250), .A2(n2736), .ZN(n2904) );
  NAND2_X1 U4143 ( .A1(n12265), .A2(n2721), .ZN(n2895) );
  NAND2_X1 U4144 ( .A1(n208), .A2(n2724), .ZN(n2910) );
  NAND2_X1 U4145 ( .A1(gte_x_382_A_16_), .A2(n2718), .ZN(n2898) );
  NAND2_X1 U4146 ( .A1(n2910), .A2(n2898), .ZN(n2892) );
  NAND2_X1 U4147 ( .A1(n12217), .A2(pmp_addr_i[46]), .ZN(n2900) );
  NOR2_X1 U4148 ( .A1(n12156), .A2(n2721), .ZN(n2897) );
  AOI22_X1 U4149 ( .A1(n2898), .A2(n2897), .B1(n1922), .B2(pmp_addr_i[48]), 
        .ZN(n2899) );
  OAI21_X1 U4150 ( .B1(n2901), .B2(n2900), .A(n2899), .ZN(n2902) );
  INV_X1 U4151 ( .A(n2902), .ZN(n2916) );
  NOR2_X1 U4152 ( .A1(n5069), .A2(n4981), .ZN(n2903) );
  AOI22_X1 U4153 ( .A1(n2904), .A2(n2903), .B1(n5070), .B2(pmp_addr_i[42]), 
        .ZN(n2909) );
  NOR2_X1 U4154 ( .A1(n5997), .A2(n4934), .ZN(n2905) );
  AOI22_X1 U4155 ( .A1(n2906), .A2(n2905), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[44]), .ZN(n2907) );
  OAI21_X1 U4156 ( .B1(n2909), .B2(n2908), .A(n2907), .ZN(n2911) );
  NAND4_X1 U4157 ( .A1(n2911), .A2(n2913), .A3(n2912), .A4(n2910), .ZN(n2915)
         );
  NAND4_X1 U4158 ( .A1(n2913), .A2(pmp_addr_i[45]), .A3(n6017), .A4(n2912), 
        .ZN(n2914) );
  NAND4_X1 U4159 ( .A1(n2917), .A2(n2916), .A3(n2915), .A4(n2914), .ZN(n2926)
         );
  INV_X1 U4160 ( .A(n2918), .ZN(n2922) );
  NAND2_X1 U4161 ( .A1(instr_addr_o_19_), .A2(n2773), .ZN(n2919) );
  AND2_X1 U4162 ( .A1(n2920), .A2(n2919), .ZN(n2921) );
  NAND3_X1 U4163 ( .A1(n2922), .A2(n2927), .A3(n2921), .ZN(n2923) );
  NOR2_X1 U4164 ( .A1(n2924), .A2(n2923), .ZN(n2925) );
  AOI22_X1 U4165 ( .A1(n2928), .A2(n2927), .B1(n2926), .B2(n2925), .ZN(n2929)
         );
  INV_X1 U4166 ( .A(pmp_cfg_i[91]), .ZN(n2993) );
  NOR2_X1 U4167 ( .A1(n2993), .A2(pmp_cfg_i[92]), .ZN(n10256) );
  INV_X1 U4168 ( .A(n10256), .ZN(n2949) );
  NAND2_X1 U4169 ( .A1(pmp_addr_i[355]), .A2(pmp_addr_i[356]), .ZN(n5933) );
  INV_X1 U4170 ( .A(n5933), .ZN(n2931) );
  INV_X1 U4171 ( .A(pmp_cfg_i[92]), .ZN(n2952) );
  NAND3_X1 U4172 ( .A1(pmp_addr_i[352]), .A2(pmp_addr_i[354]), .A3(
        pmp_addr_i[353]), .ZN(n12042) );
  OAI21_X1 U4173 ( .B1(n12042), .B2(n2993), .A(pmp_cfg_i[92]), .ZN(n2951) );
  OAI21_X1 U4174 ( .B1(n2931), .B2(n2952), .A(n2951), .ZN(n2955) );
  NAND2_X1 U4175 ( .A1(n2955), .A2(pmp_addr_i[356]), .ZN(n2932) );
  OAI21_X1 U4176 ( .B1(n3050), .B2(n2933), .A(n2932), .ZN(n10139) );
  INV_X1 U4177 ( .A(n10139), .ZN(n10306) );
  NOR2_X1 U4178 ( .A1(n5277), .A2(n10306), .ZN(n2945) );
  INV_X1 U4179 ( .A(pmp_addr_i[355]), .ZN(n5935) );
  NAND2_X1 U4180 ( .A1(n10256), .A2(pmp_addr_i[323]), .ZN(n2934) );
  OAI21_X1 U4181 ( .B1(n2951), .B2(n5935), .A(n2934), .ZN(n10307) );
  INV_X1 U4182 ( .A(n10307), .ZN(n6014) );
  NOR2_X1 U4183 ( .A1(n5280), .A2(n6014), .ZN(n2935) );
  NOR2_X1 U4184 ( .A1(n2945), .A2(n2935), .ZN(n2948) );
  NAND2_X1 U4185 ( .A1(n10256), .A2(pmp_addr_i[322]), .ZN(n2936) );
  OAI21_X1 U4186 ( .B1(n2951), .B2(n2937), .A(n2936), .ZN(n10134) );
  INV_X1 U4187 ( .A(n10134), .ZN(n12059) );
  NOR2_X1 U4188 ( .A1(n5291), .A2(n12059), .ZN(n2943) );
  AND2_X1 U4189 ( .A1(pmp_cfg_i[91]), .A2(pmp_addr_i[352]), .ZN(n2940) );
  NAND2_X1 U4190 ( .A1(pmp_cfg_i[92]), .A2(pmp_addr_i[353]), .ZN(n2939) );
  NAND2_X1 U4191 ( .A1(n10256), .A2(pmp_addr_i[321]), .ZN(n2938) );
  OAI21_X1 U4192 ( .B1(n2940), .B2(n2939), .A(n2938), .ZN(n12027) );
  INV_X1 U4193 ( .A(n12027), .ZN(n10319) );
  OR2_X1 U4194 ( .A1(n2952), .A2(pmp_cfg_i[91]), .ZN(n5963) );
  NAND2_X1 U4195 ( .A1(n10256), .A2(pmp_addr_i[320]), .ZN(n2941) );
  OAI21_X1 U4196 ( .B1(n5963), .B2(n5949), .A(n2941), .ZN(n10308) );
  INV_X1 U4197 ( .A(n10308), .ZN(n6012) );
  NAND2_X1 U4198 ( .A1(n10319), .A2(n6012), .ZN(n2942) );
  NAND2_X1 U4199 ( .A1(n12150), .A2(n12059), .ZN(n5964) );
  OAI21_X1 U4200 ( .B1(n2943), .B2(n2942), .A(n5964), .ZN(n2947) );
  NAND2_X1 U4201 ( .A1(n5280), .A2(n6014), .ZN(n2944) );
  NAND2_X1 U4202 ( .A1(n12152), .A2(n10306), .ZN(n5932) );
  OAI21_X1 U4203 ( .B1(n2945), .B2(n2944), .A(n5932), .ZN(n2946) );
  AOI21_X1 U4204 ( .B1(n2948), .B2(n2947), .A(n2946), .ZN(n2972) );
  NAND2_X1 U4205 ( .A1(pmp_addr_i[358]), .A2(pmp_addr_i[357]), .ZN(n2950) );
  OAI21_X1 U4206 ( .B1(n12021), .B2(n2952), .A(n2951), .ZN(n2961) );
  NAND2_X1 U4207 ( .A1(n2961), .A2(pmp_addr_i[358]), .ZN(n2953) );
  OAI21_X1 U4208 ( .B1(n2949), .B2(n2954), .A(n2953), .ZN(n10145) );
  INV_X1 U4209 ( .A(n10145), .ZN(n10322) );
  NOR2_X1 U4210 ( .A1(n2623), .A2(n10322), .ZN(n2966) );
  NAND2_X1 U4211 ( .A1(n2955), .A2(pmp_addr_i[357]), .ZN(n2956) );
  OAI21_X1 U4212 ( .B1(n3050), .B2(n2957), .A(n2956), .ZN(n10146) );
  INV_X1 U4213 ( .A(n10146), .ZN(n10309) );
  NOR2_X1 U4214 ( .A1(n4605), .A2(n10309), .ZN(n2958) );
  NOR2_X1 U4215 ( .A1(n2966), .A2(n2958), .ZN(n2965) );
  OR2_X1 U4216 ( .A1(n12009), .A2(n2993), .ZN(n2973) );
  NAND3_X1 U4217 ( .A1(n2973), .A2(pmp_cfg_i[92]), .A3(pmp_addr_i[360]), .ZN(
        n2960) );
  OAI21_X1 U4218 ( .B1(n2949), .B2(n1077), .A(n2960), .ZN(n10149) );
  INV_X1 U4219 ( .A(n10149), .ZN(n10317) );
  NOR2_X1 U4220 ( .A1(instr_addr_o_10_), .A2(n10317), .ZN(n2967) );
  NAND2_X1 U4221 ( .A1(n2961), .A2(pmp_addr_i[359]), .ZN(n2962) );
  OAI21_X1 U4222 ( .B1(n2949), .B2(n2963), .A(n2962), .ZN(n10148) );
  INV_X1 U4223 ( .A(n10148), .ZN(n10305) );
  NOR2_X1 U4224 ( .A1(n154), .A2(n10305), .ZN(n2964) );
  NOR2_X1 U4225 ( .A1(n2967), .A2(n2964), .ZN(n2970) );
  NAND2_X1 U4226 ( .A1(n2965), .A2(n2970), .ZN(n2971) );
  NAND2_X1 U4227 ( .A1(n5268), .A2(n10309), .ZN(n5968) );
  NAND2_X1 U4228 ( .A1(n205), .A2(n10322), .ZN(n5958) );
  OAI21_X1 U4229 ( .B1(n2966), .B2(n5968), .A(n5958), .ZN(n2969) );
  NAND2_X1 U4230 ( .A1(n5040), .A2(n10305), .ZN(n5931) );
  NAND2_X1 U4231 ( .A1(n213), .A2(n10317), .ZN(n5965) );
  OAI21_X1 U4232 ( .B1(n2967), .B2(n5931), .A(n5965), .ZN(n2968) );
  OR2_X1 U4233 ( .A1(n2973), .A2(n3127), .ZN(n2981) );
  NAND2_X1 U4234 ( .A1(pmp_addr_i[362]), .A2(pmp_addr_i[361]), .ZN(n2977) );
  NAND2_X1 U4235 ( .A1(pmp_addr_i[364]), .A2(pmp_addr_i[363]), .ZN(n2974) );
  OR2_X1 U4236 ( .A1(n2977), .A2(n2974), .ZN(n2975) );
  OAI21_X1 U4237 ( .B1(n2981), .B2(n2975), .A(pmp_cfg_i[92]), .ZN(n2989) );
  INV_X1 U4238 ( .A(pmp_addr_i[364]), .ZN(n2992) );
  NAND2_X1 U4239 ( .A1(n10256), .A2(pmp_addr_i[332]), .ZN(n2976) );
  OAI21_X1 U4240 ( .B1(n2989), .B2(n2992), .A(n2976), .ZN(n10170) );
  INV_X1 U4241 ( .A(n10170), .ZN(n10314) );
  NOR2_X1 U4242 ( .A1(n206), .A2(n10314), .ZN(n3006) );
  OAI21_X1 U4243 ( .B1(n2981), .B2(n2977), .A(pmp_cfg_i[92]), .ZN(n2985) );
  INV_X1 U4244 ( .A(pmp_addr_i[363]), .ZN(n2991) );
  NAND2_X1 U4245 ( .A1(n10256), .A2(pmp_addr_i[331]), .ZN(n2978) );
  OAI21_X1 U4246 ( .B1(n2985), .B2(n2991), .A(n2978), .ZN(n10169) );
  INV_X1 U4247 ( .A(n10169), .ZN(n10315) );
  NOR2_X1 U4248 ( .A1(n150), .A2(n10315), .ZN(n2979) );
  NOR2_X1 U4249 ( .A1(n3006), .A2(n2979), .ZN(n3009) );
  AND2_X1 U4250 ( .A1(pmp_cfg_i[92]), .A2(pmp_addr_i[361]), .ZN(n2980) );
  NAND2_X1 U4251 ( .A1(n2981), .A2(n2980), .ZN(n2982) );
  OAI21_X1 U4252 ( .B1(n2949), .B2(n1041), .A(n2982), .ZN(n10166) );
  INV_X1 U4253 ( .A(n10166), .ZN(n10318) );
  NOR2_X1 U4254 ( .A1(n5069), .A2(n10318), .ZN(n2986) );
  INV_X1 U4255 ( .A(pmp_addr_i[362]), .ZN(n2984) );
  NAND2_X1 U4256 ( .A1(n10256), .A2(pmp_addr_i[330]), .ZN(n2983) );
  OAI21_X1 U4257 ( .B1(n2985), .B2(n2984), .A(n2983), .ZN(n10167) );
  INV_X1 U4258 ( .A(n10167), .ZN(n10316) );
  NOR2_X1 U4259 ( .A1(instr_addr_o_12_), .A2(n10316), .ZN(n3005) );
  NOR2_X1 U4260 ( .A1(n2986), .A2(n3005), .ZN(n2987) );
  NAND2_X1 U4261 ( .A1(n3009), .A2(n2987), .ZN(n3004) );
  NAND2_X1 U4262 ( .A1(n10256), .A2(pmp_addr_i[333]), .ZN(n2988) );
  OAI21_X1 U4263 ( .B1(n2989), .B2(n116), .A(n2988), .ZN(n10280) );
  INV_X1 U4264 ( .A(n10280), .ZN(n3010) );
  NOR2_X1 U4265 ( .A1(instr_addr_o_15_), .A2(n3010), .ZN(n2995) );
  INV_X1 U4266 ( .A(pmp_addr_i[361]), .ZN(n2990) );
  NAND2_X1 U4267 ( .A1(n12018), .A2(pmp_addr_i[362]), .ZN(n12008) );
  OR2_X1 U4268 ( .A1(n12008), .A2(n2991), .ZN(n12041) );
  OAI211_X1 U4269 ( .C1(n115), .C2(n2993), .A(pmp_addr_i[366]), .B(
        pmp_cfg_i[92]), .ZN(n2994) );
  OAI21_X1 U4270 ( .B1(n2949), .B2(n1048), .A(n2994), .ZN(n12051) );
  INV_X1 U4271 ( .A(n12051), .ZN(n6003) );
  NOR2_X1 U4272 ( .A1(n3100), .A2(n6003), .ZN(n3012) );
  NOR2_X1 U4273 ( .A1(n2995), .A2(n3012), .ZN(n3003) );
  INV_X1 U4274 ( .A(pmp_addr_i[366]), .ZN(n2996) );
  INV_X1 U4275 ( .A(pmp_addr_i[367]), .ZN(n2997) );
  AND2_X1 U4276 ( .A1(pmp_cfg_i[91]), .A2(pmp_cfg_i[92]), .ZN(n5948) );
  NAND2_X1 U4277 ( .A1(n6011), .A2(pmp_addr_i[367]), .ZN(n2998) );
  OAI21_X1 U4278 ( .B1(n2999), .B2(n3050), .A(n2998), .ZN(n10290) );
  INV_X1 U4279 ( .A(n10290), .ZN(n5973) );
  NAND2_X1 U4281 ( .A1(n6011), .A2(pmp_addr_i[368]), .ZN(n3001) );
  OAI21_X1 U4282 ( .B1(n2949), .B2(n1050), .A(n3001), .ZN(n10298) );
  NOR2_X1 U4283 ( .A1(n3002), .A2(n3014), .ZN(n3017) );
  NAND2_X1 U4284 ( .A1(n3003), .A2(n3017), .ZN(n3019) );
  NOR2_X1 U4285 ( .A1(n3004), .A2(n3019), .ZN(n3022) );
  NAND2_X1 U4286 ( .A1(instr_addr_o_11_), .A2(n10318), .ZN(n5960) );
  NAND2_X1 U4287 ( .A1(n5250), .A2(n10316), .ZN(n5957) );
  OAI21_X1 U4288 ( .B1(n3005), .B2(n5960), .A(n5957), .ZN(n3008) );
  NAND2_X1 U4289 ( .A1(n5997), .A2(n10315), .ZN(n5967) );
  NAND2_X1 U4290 ( .A1(n5251), .A2(n10314), .ZN(n5959) );
  OAI21_X1 U4291 ( .B1(n3006), .B2(n5967), .A(n5959), .ZN(n3007) );
  AOI21_X1 U4292 ( .B1(n3009), .B2(n3008), .A(n3007), .ZN(n3020) );
  NAND2_X1 U4293 ( .A1(n208), .A2(n3010), .ZN(n3011) );
  NAND2_X1 U4294 ( .A1(n3100), .A2(n6003), .ZN(n5993) );
  OAI21_X1 U4295 ( .B1(n3012), .B2(n3011), .A(n5993), .ZN(n3016) );
  NAND2_X1 U4296 ( .A1(n5974), .A2(n5973), .ZN(n5966) );
  OAI21_X1 U4297 ( .B1(n3014), .B2(n5966), .A(n3013), .ZN(n3015) );
  AOI21_X1 U4298 ( .B1(n3016), .B2(n3017), .A(n3015), .ZN(n3018) );
  OAI21_X1 U4299 ( .B1(n3020), .B2(n3019), .A(n3018), .ZN(n3021) );
  AOI21_X1 U4300 ( .B1(n3023), .B2(n3022), .A(n3021), .ZN(n3098) );
  NAND2_X1 U4301 ( .A1(n6011), .A2(pmp_addr_i[370]), .ZN(n3024) );
  OAI21_X1 U4302 ( .B1(n2949), .B2(n1063), .A(n3024), .ZN(n10296) );
  NOR2_X1 U4303 ( .A1(n6027), .A2(n10195), .ZN(n3058) );
  NAND2_X1 U4304 ( .A1(n6011), .A2(pmp_addr_i[369]), .ZN(n3026) );
  OAI21_X1 U4305 ( .B1(n2949), .B2(n1105), .A(n3026), .ZN(n10261) );
  NOR2_X1 U4306 ( .A1(n4907), .A2(n10194), .ZN(n3027) );
  NOR2_X1 U4307 ( .A1(n3058), .A2(n3027), .ZN(n3031) );
  INV_X1 U4308 ( .A(n2103), .ZN(n4836) );
  NAND2_X1 U4309 ( .A1(n6011), .A2(pmp_addr_i[372]), .ZN(n3028) );
  OAI21_X1 U4310 ( .B1(n2949), .B2(n1061), .A(n3028), .ZN(n10270) );
  NOR2_X1 U4311 ( .A1(n12157), .A2(n10203), .ZN(n3061) );
  NAND2_X1 U4312 ( .A1(n6011), .A2(pmp_addr_i[371]), .ZN(n3029) );
  OAI21_X1 U4313 ( .B1(n2949), .B2(n1108), .A(n3029), .ZN(n10260) );
  NOR2_X1 U4314 ( .A1(n5842), .A2(n34), .ZN(n3030) );
  NOR2_X1 U4315 ( .A1(n3061), .A2(n3030), .ZN(n3064) );
  NAND2_X1 U4316 ( .A1(n3031), .A2(n3064), .ZN(n3039) );
  NAND2_X1 U4317 ( .A1(n6011), .A2(pmp_addr_i[374]), .ZN(n3032) );
  OAI21_X1 U4318 ( .B1(n3050), .B2(n1059), .A(n3032), .ZN(n10259) );
  NOR2_X1 U4319 ( .A1(n4835), .A2(n10208), .ZN(n3067) );
  NAND2_X1 U4320 ( .A1(n6011), .A2(pmp_addr_i[373]), .ZN(n3033) );
  OAI21_X1 U4321 ( .B1(n3050), .B2(n1127), .A(n3033), .ZN(n10279) );
  NOR2_X1 U4322 ( .A1(n4859), .A2(n10207), .ZN(n3034) );
  NOR2_X1 U4323 ( .A1(n3067), .A2(n3034), .ZN(n3038) );
  NAND2_X1 U4325 ( .A1(n6011), .A2(pmp_addr_i[376]), .ZN(n3035) );
  OAI21_X1 U4326 ( .B1(n3050), .B2(n1057), .A(n3035), .ZN(n10268) );
  NOR2_X1 U4327 ( .A1(n4909), .A2(n10230), .ZN(n3070) );
  NAND2_X1 U4329 ( .A1(n6011), .A2(pmp_addr_i[375]), .ZN(n3036) );
  OAI21_X1 U4330 ( .B1(n3050), .B2(n1130), .A(n3036), .ZN(n10269) );
  NOR2_X1 U4331 ( .A1(n5365), .A2(n10229), .ZN(n3037) );
  NOR2_X1 U4332 ( .A1(n3070), .A2(n3037), .ZN(n3073) );
  NAND2_X1 U4333 ( .A1(n3038), .A2(n3073), .ZN(n3075) );
  NOR2_X1 U4334 ( .A1(n3039), .A2(n3075), .ZN(n3055) );
  NAND2_X1 U4335 ( .A1(n6011), .A2(pmp_addr_i[380]), .ZN(n3040) );
  OAI21_X1 U4336 ( .B1(n3050), .B2(n1055), .A(n3040), .ZN(n10258) );
  NOR2_X1 U4337 ( .A1(n4753), .A2(n10242), .ZN(n3083) );
  NAND2_X1 U4338 ( .A1(n6011), .A2(pmp_addr_i[379]), .ZN(n3042) );
  OAI21_X1 U4339 ( .B1(n3050), .B2(n1117), .A(n3042), .ZN(n10277) );
  NOR2_X1 U4340 ( .A1(n4900), .A2(n10241), .ZN(n3043) );
  NOR2_X1 U4341 ( .A1(n3083), .A2(n3043), .ZN(n3086) );
  NAND2_X1 U4342 ( .A1(n6011), .A2(pmp_addr_i[377]), .ZN(n3044) );
  OAI21_X1 U4343 ( .B1(n3050), .B2(n1114), .A(n3044), .ZN(n10278) );
  NOR2_X1 U4344 ( .A1(instr_addr_o_27_), .A2(n10234), .ZN(n3048) );
  INV_X1 U4345 ( .A(n3045), .ZN(n4901) );
  INV_X1 U4346 ( .A(pmp_addr_i[346]), .ZN(n3047) );
  NAND2_X1 U4347 ( .A1(n6011), .A2(pmp_addr_i[378]), .ZN(n3046) );
  OAI21_X1 U4348 ( .B1(n3050), .B2(n3047), .A(n3046), .ZN(n10266) );
  INV_X1 U4349 ( .A(n10266), .ZN(n3077) );
  NOR2_X1 U4350 ( .A1(n3048), .A2(n3080), .ZN(n3049) );
  NAND2_X1 U4351 ( .A1(n3086), .A2(n3049), .ZN(n3054) );
  NAND2_X1 U4352 ( .A1(n6011), .A2(pmp_addr_i[381]), .ZN(n12066) );
  OAI21_X1 U4353 ( .B1(n3050), .B2(n1138), .A(n12066), .ZN(n10304) );
  INV_X1 U4354 ( .A(n10304), .ZN(n3087) );
  NOR2_X1 U4355 ( .A1(n4866), .A2(n3087), .ZN(n3051) );
  NOR2_X1 U4356 ( .A1(n3051), .A2(pmp_addr_i[350]), .ZN(n3053) );
  INV_X1 U4357 ( .A(pmp_addr_i[351]), .ZN(n3052) );
  NAND2_X1 U4358 ( .A1(n3053), .A2(n3052), .ZN(n3091) );
  NOR2_X1 U4359 ( .A1(n3054), .A2(n3091), .ZN(n3094) );
  NAND2_X1 U4360 ( .A1(n3055), .A2(n3094), .ZN(n3097) );
  NAND2_X1 U4361 ( .A1(n4907), .A2(n10194), .ZN(n3057) );
  NAND2_X1 U4362 ( .A1(n6027), .A2(n10195), .ZN(n3056) );
  OAI21_X1 U4363 ( .B1(n3058), .B2(n3057), .A(n3056), .ZN(n3063) );
  NAND2_X1 U4364 ( .A1(n5842), .A2(n34), .ZN(n3060) );
  NAND2_X1 U4365 ( .A1(n4836), .A2(n10203), .ZN(n3059) );
  OAI21_X1 U4366 ( .B1(n3061), .B2(n3060), .A(n3059), .ZN(n3062) );
  AOI21_X1 U4367 ( .B1(n3064), .B2(n3063), .A(n3062), .ZN(n3076) );
  NAND2_X1 U4368 ( .A1(n4859), .A2(n10207), .ZN(n3066) );
  NAND2_X1 U4369 ( .A1(n4835), .A2(n10208), .ZN(n3065) );
  OAI21_X1 U4370 ( .B1(n3067), .B2(n3066), .A(n3065), .ZN(n3072) );
  NAND2_X1 U4371 ( .A1(instr_addr_o_25_), .A2(n10229), .ZN(n3069) );
  NAND2_X1 U4372 ( .A1(n4909), .A2(n10230), .ZN(n3068) );
  OAI21_X1 U4373 ( .B1(n3070), .B2(n3069), .A(n3068), .ZN(n3071) );
  AOI21_X1 U4374 ( .B1(n3073), .B2(n3072), .A(n3071), .ZN(n3074) );
  OAI21_X1 U4375 ( .B1(n3076), .B2(n3075), .A(n3074), .ZN(n3095) );
  NAND2_X1 U4376 ( .A1(n12195), .A2(n10234), .ZN(n3079) );
  NAND2_X1 U4377 ( .A1(n4901), .A2(n3077), .ZN(n3078) );
  OAI21_X1 U4378 ( .B1(n3080), .B2(n3079), .A(n3078), .ZN(n3085) );
  NAND2_X1 U4379 ( .A1(n4900), .A2(n10241), .ZN(n3082) );
  NAND2_X1 U4380 ( .A1(n5980), .A2(n10242), .ZN(n3081) );
  OAI21_X1 U4381 ( .B1(n3083), .B2(n3082), .A(n3081), .ZN(n3084) );
  AOI21_X1 U4382 ( .B1(n3086), .B2(n3085), .A(n3084), .ZN(n3092) );
  NAND2_X1 U4383 ( .A1(n6018), .A2(n3087), .ZN(n3088) );
  NOR2_X1 U4384 ( .A1(n3088), .A2(pmp_addr_i[350]), .ZN(n3089) );
  NAND2_X1 U4385 ( .A1(n3089), .A2(n3052), .ZN(n3090) );
  OAI21_X1 U4386 ( .B1(n3092), .B2(n3091), .A(n3090), .ZN(n3093) );
  AOI21_X1 U4387 ( .B1(n3095), .B2(n3094), .A(n3093), .ZN(n3096) );
  INV_X1 U4388 ( .A(pmp_addr_i[368]), .ZN(n3099) );
  NAND2_X1 U4389 ( .A1(n5047), .A2(n3099), .ZN(n3111) );
  NAND2_X1 U4390 ( .A1(n5229), .A2(n2996), .ZN(n3109) );
  OAI21_X1 U4391 ( .B1(n6017), .B2(pmp_addr_i[365]), .A(n3109), .ZN(n3101) );
  NOR2_X1 U4392 ( .A1(n3113), .A2(n3101), .ZN(n3144) );
  NAND2_X1 U4393 ( .A1(n5245), .A2(n2984), .ZN(n3135) );
  NOR2_X1 U4394 ( .A1(n5069), .A2(n2990), .ZN(n3102) );
  AOI22_X1 U4395 ( .A1(n3135), .A2(n3102), .B1(n5070), .B2(pmp_addr_i[362]), 
        .ZN(n3107) );
  NAND2_X1 U4396 ( .A1(n4788), .A2(n2992), .ZN(n3105) );
  NAND2_X1 U4397 ( .A1(n4061), .A2(n2991), .ZN(n3103) );
  NAND2_X1 U4398 ( .A1(n3105), .A2(n3103), .ZN(n3137) );
  NOR2_X1 U4399 ( .A1(n150), .A2(n2991), .ZN(n3104) );
  AOI22_X1 U4400 ( .A1(n3105), .A2(n3104), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[364]), .ZN(n3106) );
  OAI21_X1 U4401 ( .B1(n3107), .B2(n3137), .A(n3106), .ZN(n3116) );
  NOR2_X1 U4402 ( .A1(instr_addr_o_15_), .A2(n116), .ZN(n3108) );
  AOI22_X1 U4403 ( .A1(n3109), .A2(n3108), .B1(n5058), .B2(pmp_addr_i[366]), 
        .ZN(n3114) );
  AOI22_X1 U4405 ( .A1(n3111), .A2(n3110), .B1(n1922), .B2(pmp_addr_i[368]), 
        .ZN(n3112) );
  OAI21_X1 U4406 ( .B1(n3114), .B2(n3113), .A(n3112), .ZN(n3115) );
  AOI21_X1 U4407 ( .B1(n3144), .B2(n3116), .A(n3115), .ZN(n3162) );
  INV_X1 U4408 ( .A(pmp_addr_i[356]), .ZN(n3122) );
  NOR2_X1 U4409 ( .A1(instr_addr_o_6_), .A2(n3122), .ZN(n3126) );
  NOR2_X1 U4410 ( .A1(pmp_addr_i[353]), .A2(pmp_addr_i[352]), .ZN(n3117) );
  OAI22_X1 U4411 ( .A1(n6015), .A2(n5935), .B1(n3117), .B2(n2937), .ZN(n3121)
         );
  INV_X1 U4412 ( .A(n3117), .ZN(n3118) );
  NOR2_X1 U4413 ( .A1(n3118), .A2(pmp_addr_i[354]), .ZN(n3119) );
  NOR2_X1 U4414 ( .A1(n5291), .A2(n3119), .ZN(n3120) );
  NOR3_X1 U4415 ( .A1(n3126), .A2(n3121), .A3(n3120), .ZN(n3134) );
  NAND2_X1 U4416 ( .A1(n5293), .A2(n5935), .ZN(n3125) );
  INV_X1 U4417 ( .A(pmp_addr_i[357]), .ZN(n3129) );
  AOI22_X1 U4418 ( .A1(instr_addr_o_6_), .A2(n3122), .B1(n4605), .B2(n3129), 
        .ZN(n3124) );
  INV_X1 U4419 ( .A(pmp_addr_i[358]), .ZN(n3123) );
  NAND2_X1 U4420 ( .A1(instr_addr_o_8_), .A2(n3123), .ZN(n3131) );
  OAI211_X1 U4421 ( .C1(n3126), .C2(n3125), .A(n3124), .B(n3131), .ZN(n3133)
         );
  NOR2_X1 U4422 ( .A1(n153), .A2(n2959), .ZN(n3128) );
  INV_X1 U4423 ( .A(pmp_addr_i[360]), .ZN(n3127) );
  NAND2_X1 U4424 ( .A1(n5262), .A2(n3127), .ZN(n3139) );
  AOI22_X1 U4425 ( .A1(n3128), .A2(n3139), .B1(n4602), .B2(pmp_addr_i[360]), 
        .ZN(n3141) );
  NOR2_X1 U4426 ( .A1(n4605), .A2(n3129), .ZN(n3130) );
  AOI22_X1 U4427 ( .A1(n3131), .A2(n3130), .B1(n4606), .B2(pmp_addr_i[358]), 
        .ZN(n3132) );
  OAI211_X1 U4428 ( .C1(n3134), .C2(n3133), .A(n3141), .B(n3132), .ZN(n3145)
         );
  OAI21_X1 U4429 ( .B1(n5052), .B2(pmp_addr_i[361]), .A(n3135), .ZN(n3136) );
  NOR2_X1 U4430 ( .A1(n3137), .A2(n3136), .ZN(n3143) );
  NAND2_X1 U4431 ( .A1(n154), .A2(n2959), .ZN(n3138) );
  NAND2_X1 U4432 ( .A1(n3139), .A2(n3138), .ZN(n3140) );
  NAND2_X1 U4433 ( .A1(n3141), .A2(n3140), .ZN(n3142) );
  NAND4_X1 U4434 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), .ZN(n3161)
         );
  INV_X1 U4435 ( .A(pmp_addr_i[378]), .ZN(n3146) );
  INV_X1 U4436 ( .A(pmp_addr_i[376]), .ZN(n3147) );
  NAND2_X1 U4437 ( .A1(n210), .A2(n3147), .ZN(n3181) );
  INV_X1 U4438 ( .A(pmp_addr_i[375]), .ZN(n3179) );
  NAND2_X1 U4439 ( .A1(n5202), .A2(n3179), .ZN(n3148) );
  NAND2_X1 U4440 ( .A1(n3181), .A2(n3148), .ZN(n3183) );
  NOR2_X1 U4441 ( .A1(n3183), .A2(n3163), .ZN(n3159) );
  BUF_X1 U4442 ( .A(n3192), .Z(n4406) );
  INV_X1 U4443 ( .A(pmp_addr_i[380]), .ZN(n3149) );
  NAND2_X1 U4444 ( .A1(n12161), .A2(n3149), .ZN(n3193) );
  NAND2_X1 U4445 ( .A1(n5136), .A2(n1499), .ZN(n3194) );
  INV_X1 U4446 ( .A(pmp_addr_i[370]), .ZN(n3150) );
  NAND2_X1 U4447 ( .A1(n5187), .A2(n3150), .ZN(n3167) );
  OAI211_X1 U4448 ( .C1(n5313), .C2(pmp_addr_i[369]), .A(n3194), .B(n3167), 
        .ZN(n3151) );
  NOR2_X1 U4449 ( .A1(n3188), .A2(n3151), .ZN(n3158) );
  INV_X1 U4450 ( .A(pmp_addr_i[371]), .ZN(n3169) );
  NAND2_X1 U4451 ( .A1(n3152), .A2(n3169), .ZN(n3154) );
  INV_X1 U4452 ( .A(pmp_addr_i[372]), .ZN(n3153) );
  INV_X1 U4455 ( .A(pmp_addr_i[374]), .ZN(n3155) );
  NAND2_X1 U4456 ( .A1(instr_addr_o_24_), .A2(n3155), .ZN(n3178) );
  INV_X1 U4457 ( .A(pmp_addr_i[373]), .ZN(n3176) );
  NAND2_X1 U4458 ( .A1(n5208), .A2(n3176), .ZN(n3156) );
  AND2_X1 U4459 ( .A1(n3178), .A2(n3156), .ZN(n3174) );
  NAND4_X1 U4460 ( .A1(n3159), .A2(n3158), .A3(n3157), .A4(n3174), .ZN(n3160)
         );
  AOI21_X1 U4461 ( .B1(n3162), .B2(n3161), .A(n3160), .ZN(n3204) );
  INV_X1 U4462 ( .A(n3163), .ZN(n3164) );
  AND3_X1 U4463 ( .A1(n3164), .A2(n3165), .A3(n3194), .ZN(n3186) );
  INV_X1 U4464 ( .A(n3183), .ZN(n3175) );
  INV_X1 U4465 ( .A(pmp_addr_i[369]), .ZN(n3166) );
  NOR2_X1 U4466 ( .A1(n5100), .A2(n3166), .ZN(n3168) );
  AOI22_X1 U4467 ( .A1(n3168), .A2(n3167), .B1(n4631), .B2(pmp_addr_i[370]), 
        .ZN(n3173) );
  NOR2_X1 U4468 ( .A1(n5842), .A2(n3169), .ZN(n3171) );
  NOR2_X1 U4469 ( .A1(n5208), .A2(n3176), .ZN(n3177) );
  AOI22_X1 U4470 ( .A1(n3178), .A2(n3177), .B1(n2580), .B2(pmp_addr_i[374]), 
        .ZN(n3184) );
  NOR2_X1 U4471 ( .A1(n12226), .A2(n3179), .ZN(n3180) );
  AOI22_X1 U4472 ( .A1(n3181), .A2(n3180), .B1(n3806), .B2(pmp_addr_i[376]), 
        .ZN(n3182) );
  OAI21_X1 U4473 ( .B1(n3184), .B2(n3183), .A(n3182), .ZN(n3185) );
  NAND2_X1 U4474 ( .A1(n139), .A2(n3185), .ZN(n3201) );
  INV_X1 U4475 ( .A(n3194), .ZN(n3187) );
  NOR2_X1 U4476 ( .A1(n3188), .A2(n3187), .ZN(n3199) );
  NAND3_X1 U4477 ( .A1(n3189), .A2(pmp_addr_i[377]), .A3(n4147), .ZN(n3191) );
  NAND2_X1 U4478 ( .A1(n4438), .A2(pmp_addr_i[378]), .ZN(n3190) );
  NAND2_X1 U4479 ( .A1(n3191), .A2(n3190), .ZN(n3198) );
  BUF_X1 U4480 ( .A(n3192), .Z(n4623) );
  NAND4_X1 U4481 ( .A1(n3193), .A2(n3194), .A3(pmp_addr_i[379]), .A4(n4623), 
        .ZN(n3197) );
  NAND3_X1 U4482 ( .A1(n3194), .A2(pmp_addr_i[380]), .A3(n4658), .ZN(n3196) );
  NAND2_X1 U4483 ( .A1(n4660), .A2(pmp_addr_i[381]), .ZN(n3195) );
  NAND3_X1 U4484 ( .A1(n3202), .A2(n3201), .A3(n3200), .ZN(n3203) );
  OR2_X1 U4485 ( .A1(n3204), .A2(n3203), .ZN(n3205) );
  INV_X1 U4486 ( .A(n3206), .ZN(n11098) );
  OR2_X1 U4487 ( .A1(n3208), .A2(n3207), .ZN(n11120) );
  OAI21_X1 U4488 ( .B1(n3209), .B2(n11098), .A(n11120), .ZN(n3216) );
  NOR2_X1 U4489 ( .A1(n3229), .A2(n3903), .ZN(n11090) );
  NOR2_X1 U4490 ( .A1(n7791), .A2(n11090), .ZN(n3211) );
  NAND2_X1 U4491 ( .A1(n11090), .A2(pmp_addr_i[457]), .ZN(n3217) );
  OR2_X1 U4492 ( .A1(n3217), .A2(n2634), .ZN(n11115) );
  NOR2_X1 U4493 ( .A1(n11115), .A2(n2650), .ZN(n11114) );
  NOR2_X1 U4494 ( .A1(n11114), .A2(n7793), .ZN(n3210) );
  AOI22_X1 U4495 ( .A1(n3934), .A2(n3211), .B1(n12180), .B2(n3210), .ZN(n3215)
         );
  INV_X1 U4496 ( .A(n11120), .ZN(n3212) );
  NAND2_X1 U4497 ( .A1(n3212), .A2(pmp_addr_i[451]), .ZN(n11087) );
  NAND3_X1 U4498 ( .A1(n12152), .A2(n7656), .A3(n11087), .ZN(n3214) );
  INV_X1 U4499 ( .A(n11106), .ZN(n3231) );
  NAND3_X1 U4500 ( .A1(n4605), .A2(n7648), .A3(n3231), .ZN(n3213) );
  NAND4_X1 U4501 ( .A1(n3216), .A2(n3215), .A3(n3214), .A4(n3213), .ZN(n3224)
         );
  INV_X1 U4502 ( .A(n11094), .ZN(n3218) );
  INV_X1 U4503 ( .A(n3217), .ZN(n11125) );
  OAI22_X1 U4504 ( .A1(n3218), .A2(n3248), .B1(n3247), .B2(n11125), .ZN(n3223)
         );
  NAND2_X1 U4505 ( .A1(n12150), .A2(n11103), .ZN(n3251) );
  INV_X1 U4506 ( .A(n3219), .ZN(n11100) );
  NAND2_X1 U4507 ( .A1(n11114), .A2(pmp_addr_i[460]), .ZN(n11109) );
  NAND3_X1 U4508 ( .A1(n208), .A2(n7651), .A3(n11109), .ZN(n3221) );
  NAND3_X1 U4509 ( .A1(instr_addr_o_13_), .A2(n7647), .A3(n11115), .ZN(n3220)
         );
  OAI211_X1 U4510 ( .C1(n3251), .C2(n11100), .A(n3221), .B(n3220), .ZN(n3222)
         );
  NOR3_X1 U4511 ( .A1(n3224), .A2(n3223), .A3(n3222), .ZN(n3259) );
  OR2_X1 U4512 ( .A1(n11109), .A2(n3226), .ZN(n11134) );
  INV_X1 U4513 ( .A(n11134), .ZN(n3227) );
  NAND2_X1 U4514 ( .A1(n3227), .A2(n7715), .ZN(n3236) );
  AND2_X1 U4515 ( .A1(pmp_addr_i[454]), .A2(pmp_addr_i[453]), .ZN(n3234) );
  INV_X1 U4516 ( .A(n3228), .ZN(n4743) );
  AND2_X1 U4518 ( .A1(n11134), .A2(n7655), .ZN(n11138) );
  INV_X1 U4519 ( .A(n3229), .ZN(n11111) );
  NOR2_X1 U4520 ( .A1(n7821), .A2(n11111), .ZN(n3230) );
  AOI22_X1 U4521 ( .A1(n12203), .A2(n11138), .B1(n214), .B2(n3230), .ZN(n3233)
         );
  NAND3_X1 U4522 ( .A1(instr_addr_o_9_), .A2(n7667), .A3(n3231), .ZN(n3232) );
  OAI211_X1 U4523 ( .C1(n3238), .C2(n3234), .A(n3233), .B(n3232), .ZN(n3235)
         );
  AOI21_X1 U4524 ( .B1(n3237), .B2(n3236), .A(n3235), .ZN(n3258) );
  NAND4_X1 U4525 ( .A1(n3243), .A2(n3242), .A3(n3241), .A4(n3240), .ZN(n3244)
         );
  NOR2_X1 U4526 ( .A1(n3245), .A2(n3244), .ZN(n3257) );
  NAND4_X1 U4527 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3255)
         );
  INV_X1 U4528 ( .A(n3250), .ZN(n7658) );
  NAND4_X1 U4529 ( .A1(n3253), .A2(n3252), .A3(n3251), .A4(n7658), .ZN(n3254)
         );
  NOR2_X1 U4530 ( .A1(n3255), .A2(n3254), .ZN(n3256) );
  AOI22_X1 U4531 ( .A1(n3259), .A2(n3258), .B1(n3257), .B2(n3256), .ZN(n3408)
         );
  NOR2_X1 U4532 ( .A1(n3261), .A2(n3260), .ZN(n3265) );
  XNOR2_X1 U4533 ( .A(n6020), .B(n7862), .ZN(n3264) );
  XNOR2_X1 U4534 ( .A(n5550), .B(n7870), .ZN(n3263) );
  XNOR2_X1 U4535 ( .A(n5985), .B(n7856), .ZN(n3262) );
  NAND4_X1 U4536 ( .A1(n3265), .A2(n3264), .A3(n3263), .A4(n3262), .ZN(n3274)
         );
  OAI211_X1 U4537 ( .C1(n12150), .C2(n11103), .A(n3266), .B(pmp_cfg_i[114]), 
        .ZN(n3267) );
  NOR2_X1 U4538 ( .A1(n3268), .A2(n3267), .ZN(n3272) );
  XNOR2_X1 U4539 ( .A(n6019), .B(n7786), .ZN(n3271) );
  XNOR2_X1 U4540 ( .A(n4533), .B(n7859), .ZN(n3270) );
  INV_X1 U4541 ( .A(n1632), .ZN(n5980) );
  XNOR2_X1 U4542 ( .A(n5980), .B(n7871), .ZN(n3269) );
  NAND4_X1 U4543 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n3273)
         );
  NOR2_X1 U4544 ( .A1(n3274), .A2(n3273), .ZN(n3307) );
  XNOR2_X1 U4545 ( .A(n5162), .B(n7867), .ZN(n3279) );
  XNOR2_X1 U4546 ( .A(n6028), .B(n7853), .ZN(n3276) );
  NAND4_X1 U4547 ( .A1(n3279), .A2(n3278), .A3(n12227), .A4(n3276), .ZN(n3283)
         );
  INV_X1 U4548 ( .A(n3045), .ZN(n5979) );
  XNOR2_X1 U4549 ( .A(n146), .B(n7868), .ZN(n3281) );
  XNOR2_X1 U4550 ( .A(instr_addr_o_25_), .B(n7855), .ZN(n3280) );
  NAND2_X1 U4551 ( .A1(n3281), .A2(n3280), .ZN(n3282) );
  NOR2_X1 U4552 ( .A1(n3283), .A2(n3282), .ZN(n3306) );
  NAND4_X1 U4553 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3294)
         );
  INV_X2 U4554 ( .A(n3288), .ZN(instr_addr_o_22_) );
  XNOR2_X1 U4555 ( .A(instr_addr_o_22_), .B(n3289), .ZN(n3293) );
  INV_X2 U4556 ( .A(n3290), .ZN(n6027) );
  XNOR2_X1 U4557 ( .A(n4802), .B(n3291), .ZN(n3292) );
  NOR3_X1 U4558 ( .A1(n3294), .A2(n3293), .A3(n3292), .ZN(n3305) );
  INV_X1 U4559 ( .A(n3295), .ZN(instr_addr_o_31_) );
  XNOR2_X1 U4560 ( .A(instr_addr_o_31_), .B(n7874), .ZN(n3296) );
  NAND3_X1 U4561 ( .A1(n3298), .A2(n3297), .A3(n3296), .ZN(n3303) );
  XNOR2_X1 U4562 ( .A(n6025), .B(n7852), .ZN(n3299) );
  NAND3_X1 U4563 ( .A1(n3301), .A2(n3300), .A3(n3299), .ZN(n3302) );
  NOR2_X1 U4564 ( .A1(n3303), .A2(n3302), .ZN(n3304) );
  NAND4_X1 U4565 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .ZN(n3407)
         );
  INV_X1 U4566 ( .A(n3308), .ZN(n3312) );
  XNOR2_X1 U4567 ( .A(n4859), .B(n9260), .ZN(n3311) );
  INV_X1 U4568 ( .A(n3309), .ZN(n3310) );
  INV_X1 U4569 ( .A(n3313), .ZN(n3319) );
  INV_X1 U4570 ( .A(n3314), .ZN(n3318) );
  INV_X1 U4571 ( .A(n3315), .ZN(n3317) );
  AND4_X1 U4572 ( .A1(n3319), .A2(n3318), .A3(n3317), .A4(n3316), .ZN(n3327)
         );
  XNOR2_X1 U4573 ( .A(n6020), .B(n9270), .ZN(n3326) );
  NOR2_X1 U4574 ( .A1(n3324), .A2(n334), .ZN(n3325) );
  NAND4_X1 U4575 ( .A1(n3328), .A2(n3327), .A3(n3326), .A4(n3325), .ZN(n3349)
         );
  INV_X1 U4576 ( .A(n3329), .ZN(n3333) );
  XNOR2_X1 U4577 ( .A(n6028), .B(n9261), .ZN(n3332) );
  INV_X1 U4578 ( .A(n3330), .ZN(n3331) );
  AND3_X1 U4579 ( .A1(n3333), .A2(n3332), .A3(n3331), .ZN(n3339) );
  XNOR2_X1 U4580 ( .A(instr_addr_o_28_), .B(n9276), .ZN(n3338) );
  XNOR2_X1 U4581 ( .A(n4644), .B(n9263), .ZN(n3337) );
  XNOR2_X1 U4582 ( .A(instr_addr_o_22_), .B(n9268), .ZN(n3335) );
  XNOR2_X1 U4583 ( .A(n6027), .B(n9271), .ZN(n3334) );
  OAI21_X1 U4586 ( .B1(n5976), .B2(n9059), .A(n3340), .ZN(n3341) );
  NOR2_X1 U4587 ( .A1(n3342), .A2(n3341), .ZN(n3346) );
  XNOR2_X1 U4588 ( .A(n5985), .B(n9264), .ZN(n3345) );
  XNOR2_X1 U4589 ( .A(instr_addr_o_21_), .B(n9267), .ZN(n3344) );
  XNOR2_X1 U4590 ( .A(n134), .B(n9275), .ZN(n3343) );
  NAND4_X1 U4591 ( .A1(n3346), .A2(n3345), .A3(n3344), .A4(n3343), .ZN(n3347)
         );
  NOR3_X1 U4592 ( .A1(n3349), .A2(n3348), .A3(n3347), .ZN(n3406) );
  INV_X1 U4593 ( .A(n3384), .ZN(n3354) );
  INV_X1 U4594 ( .A(n3396), .ZN(n3353) );
  AND2_X1 U4595 ( .A1(n3373), .A2(pmp_addr_i[322]), .ZN(n3372) );
  NAND2_X1 U4596 ( .A1(n3350), .A2(n3372), .ZN(n11644) );
  OR2_X1 U4597 ( .A1(n11644), .A2(n1077), .ZN(n11676) );
  INV_X1 U4598 ( .A(n3351), .ZN(n3352) );
  NOR2_X1 U4599 ( .A1(n11676), .A2(n3352), .ZN(n3376) );
  NAND2_X1 U4600 ( .A1(n3376), .A2(pmp_addr_i[331]), .ZN(n11668) );
  AOI22_X1 U4601 ( .A1(n3354), .A2(n11648), .B1(n3353), .B2(n11668), .ZN(n3355) );
  XNOR2_X1 U4602 ( .A(n5136), .B(n9282), .ZN(n3400) );
  XNOR2_X1 U4603 ( .A(n5550), .B(n9278), .ZN(n3399) );
  XNOR2_X1 U4604 ( .A(n5980), .B(n9279), .ZN(n3398) );
  NAND4_X1 U4605 ( .A1(n3355), .A2(n3400), .A3(n3399), .A4(n3398), .ZN(n3405)
         );
  NAND3_X1 U4606 ( .A1(instr_addr_o_11_), .A2(n9073), .A3(n11676), .ZN(n3363)
         );
  INV_X1 U4607 ( .A(n3372), .ZN(n11686) );
  INV_X1 U4608 ( .A(pmp_addr_i[323]), .ZN(n3356) );
  OR2_X1 U4609 ( .A1(n11686), .A2(n3356), .ZN(n3358) );
  INV_X1 U4610 ( .A(n3358), .ZN(n3357) );
  NAND2_X1 U4611 ( .A1(n3357), .A2(pmp_addr_i[324]), .ZN(n11653) );
  NAND3_X1 U4612 ( .A1(n4605), .A2(n9058), .A3(n11653), .ZN(n3362) );
  NAND3_X1 U4613 ( .A1(instr_addr_o_6_), .A2(n9071), .A3(n3358), .ZN(n3361) );
  INV_X1 U4614 ( .A(n11653), .ZN(n3359) );
  NAND2_X1 U4615 ( .A1(n3359), .A2(pmp_addr_i[325]), .ZN(n11655) );
  NAND3_X1 U4616 ( .A1(instr_addr_o_8_), .A2(n9075), .A3(n11655), .ZN(n3360)
         );
  NAND4_X1 U4617 ( .A1(n3363), .A2(n3362), .A3(n3361), .A4(n3360), .ZN(n3371)
         );
  INV_X1 U4618 ( .A(n11644), .ZN(n3364) );
  NAND3_X1 U4619 ( .A1(n3364), .A2(pmp_addr_i[328]), .A3(pmp_addr_i[329]), 
        .ZN(n3365) );
  NAND3_X1 U4620 ( .A1(n5245), .A2(n9072), .A3(n3365), .ZN(n3370) );
  NAND3_X1 U4621 ( .A1(n12156), .A2(n9077), .A3(n11689), .ZN(n3369) );
  NAND3_X1 U4622 ( .A1(n5262), .A2(n9074), .A3(n11644), .ZN(n3368) );
  NOR2_X1 U4623 ( .A1(n11681), .A2(n3366), .ZN(n11680) );
  NAND2_X1 U4624 ( .A1(n5226), .A2(n11680), .ZN(n3367) );
  NOR2_X1 U4625 ( .A1(n9221), .A2(n3372), .ZN(n3375) );
  INV_X1 U4626 ( .A(n3373), .ZN(n11662) );
  OR2_X1 U4627 ( .A1(n3374), .A2(n9329), .ZN(n9333) );
  NAND3_X1 U4628 ( .A1(n9333), .A2(pmp_cfg_i[84]), .A3(pmp_cfg_i[82]), .ZN(
        n3385) );
  AOI211_X1 U4629 ( .C1(n6015), .C2(n3375), .A(n11662), .B(n3385), .ZN(n3380)
         );
  INV_X1 U4630 ( .A(n3390), .ZN(n3377) );
  INV_X1 U4631 ( .A(n3376), .ZN(n11650) );
  NAND2_X1 U4632 ( .A1(n3377), .A2(n11650), .ZN(n3379) );
  INV_X1 U4633 ( .A(n3846), .ZN(n4204) );
  OAI211_X1 U4634 ( .C1(n11642), .C2(n11686), .A(n4204), .B(n9070), .ZN(n3378)
         );
  AND4_X1 U4635 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(n3393)
         );
  AOI21_X1 U4636 ( .B1(n5976), .B2(n9059), .A(n3385), .ZN(n3392) );
  AND4_X1 U4637 ( .A1(n3389), .A2(n3388), .A3(n3387), .A4(n3386), .ZN(n3391)
         );
  NAND4_X1 U4638 ( .A1(n3393), .A2(n3392), .A3(n3391), .A4(n3390), .ZN(n3403)
         );
  AND4_X1 U4639 ( .A1(n3397), .A2(n3396), .A3(n3395), .A4(n3394), .ZN(n3401)
         );
  NAND4_X1 U4640 ( .A1(n3401), .A2(n3400), .A3(n3399), .A4(n3398), .ZN(n3402)
         );
  NOR2_X1 U4641 ( .A1(n3410), .A2(n3409), .ZN(n3416) );
  NOR2_X1 U4642 ( .A1(n3412), .A2(n3411), .ZN(n3415) );
  XNOR2_X1 U4643 ( .A(n4909), .B(n8636), .ZN(n3414) );
  XNOR2_X1 U4644 ( .A(instr_addr_o_21_), .B(n8642), .ZN(n3413) );
  NAND4_X1 U4645 ( .A1(n3416), .A2(n3415), .A3(n3414), .A4(n3413), .ZN(n3425)
         );
  XNOR2_X1 U4646 ( .A(n6018), .B(n8584), .ZN(n3417) );
  OAI21_X1 U4647 ( .B1(n3418), .B2(n11420), .A(n3417), .ZN(n3424) );
  NAND2_X1 U4648 ( .A1(n11420), .A2(pmp_addr_i[388]), .ZN(n11423) );
  INV_X1 U4649 ( .A(pmp_addr_i[389]), .ZN(n3518) );
  OR2_X1 U4650 ( .A1(n11423), .A2(n3518), .ZN(n11406) );
  NOR2_X1 U4651 ( .A1(n11406), .A2(n1577), .ZN(n11411) );
  INV_X1 U4652 ( .A(n3419), .ZN(n3422) );
  NAND2_X1 U4653 ( .A1(n11411), .A2(pmp_addr_i[391]), .ZN(n11410) );
  OR2_X1 U4654 ( .A1(n11410), .A2(n1586), .ZN(n3437) );
  NOR2_X1 U4655 ( .A1(n3437), .A2(n3420), .ZN(n11438) );
  AND2_X1 U4656 ( .A1(n11438), .A2(pmp_addr_i[394]), .ZN(n11450) );
  OAI22_X1 U4657 ( .A1(n11411), .A2(n3422), .B1(n3421), .B2(n11450), .ZN(n3423) );
  NOR3_X1 U4658 ( .A1(n3425), .A2(n3424), .A3(n3423), .ZN(n3496) );
  NOR2_X1 U4659 ( .A1(n3427), .A2(n3426), .ZN(n3436) );
  XNOR2_X1 U4660 ( .A(n6025), .B(n8643), .ZN(n3435) );
  INV_X1 U4661 ( .A(n3428), .ZN(n3430) );
  INV_X1 U4662 ( .A(n11438), .ZN(n3429) );
  NAND2_X1 U4663 ( .A1(n3430), .A2(n3429), .ZN(n3434) );
  INV_X1 U4664 ( .A(n3431), .ZN(n3432) );
  NAND2_X1 U4665 ( .A1(n3432), .A2(n11406), .ZN(n3433) );
  NAND4_X1 U4666 ( .A1(n3436), .A2(n3435), .A3(n3434), .A4(n3433), .ZN(n3449)
         );
  INV_X1 U4667 ( .A(n3437), .ZN(n11435) );
  INV_X1 U4668 ( .A(n3438), .ZN(n3440) );
  OAI211_X1 U4669 ( .C1(n11435), .C2(n3441), .A(n3440), .B(n3439), .ZN(n3448)
         );
  INV_X1 U4670 ( .A(n11423), .ZN(n3446) );
  INV_X1 U4671 ( .A(n3442), .ZN(n3443) );
  OAI211_X1 U4672 ( .C1(n3446), .C2(n3445), .A(n3444), .B(n3443), .ZN(n3447)
         );
  NOR3_X1 U4673 ( .A1(n3449), .A2(n3448), .A3(n3447), .ZN(n3495) );
  NOR2_X1 U4674 ( .A1(n3451), .A2(n3450), .ZN(n3460) );
  XNOR2_X1 U4675 ( .A(n4835), .B(n8635), .ZN(n3459) );
  INV_X1 U4676 ( .A(n3452), .ZN(n3456) );
  INV_X1 U4677 ( .A(n3463), .ZN(n3453) );
  NAND2_X1 U4678 ( .A1(n3453), .A2(pmp_addr_i[396]), .ZN(n3454) );
  OR2_X1 U4679 ( .A1(n11410), .A2(n3454), .ZN(n11442) );
  NOR2_X1 U4680 ( .A1(n11442), .A2(n3455), .ZN(n3462) );
  NAND2_X1 U4681 ( .A1(n3462), .A2(pmp_addr_i[398]), .ZN(n11448) );
  NAND2_X1 U4682 ( .A1(n3456), .A2(n11448), .ZN(n3458) );
  XNOR2_X1 U4683 ( .A(n4836), .B(n8634), .ZN(n3457) );
  NAND4_X1 U4684 ( .A1(n3460), .A2(n3459), .A3(n3458), .A4(n3457), .ZN(n3473)
         );
  INV_X1 U4685 ( .A(n3461), .ZN(n11434) );
  INV_X1 U4686 ( .A(n3462), .ZN(n11446) );
  NAND3_X1 U4687 ( .A1(instr_addr_o_16_), .A2(n11409), .A3(n11446), .ZN(n3465)
         );
  OR2_X1 U4688 ( .A1(n11410), .A2(n3463), .ZN(n11453) );
  NAND3_X1 U4689 ( .A1(n12181), .A2(n8679), .A3(n11453), .ZN(n3464) );
  OAI211_X1 U4690 ( .C1(n3466), .C2(n11434), .A(n3465), .B(n3464), .ZN(n3472)
         );
  INV_X1 U4691 ( .A(n3467), .ZN(n3470) );
  XNOR2_X1 U4692 ( .A(n4802), .B(n8641), .ZN(n3469) );
  NAND3_X1 U4693 ( .A1(n208), .A2(n8678), .A3(n11442), .ZN(n3468) );
  NAND3_X1 U4694 ( .A1(n3470), .A2(n3469), .A3(n3468), .ZN(n3471) );
  NOR3_X1 U4695 ( .A1(n3473), .A2(n3472), .A3(n3471), .ZN(n3494) );
  NAND3_X1 U4696 ( .A1(n5270), .A2(n8670), .A3(n11410), .ZN(n3481) );
  INV_X1 U4697 ( .A(n3474), .ZN(n11425) );
  NOR2_X1 U4698 ( .A1(n8530), .A2(n11425), .ZN(n3479) );
  NAND2_X1 U4699 ( .A1(n3476), .A2(n3475), .ZN(n8706) );
  NAND4_X1 U4700 ( .A1(n8706), .A2(n3477), .A3(pmp_cfg_i[100]), .A4(
        pmp_cfg_i[98]), .ZN(n3478) );
  AOI21_X1 U4701 ( .B1(n5976), .B2(n3479), .A(n3478), .ZN(n3480) );
  OAI211_X1 U4702 ( .C1(n12150), .C2(n8661), .A(n3481), .B(n3480), .ZN(n3482)
         );
  INV_X1 U4703 ( .A(n3482), .ZN(n3486) );
  XNOR2_X1 U4704 ( .A(n5980), .B(n8651), .ZN(n3485) );
  XNOR2_X1 U4705 ( .A(n5365), .B(n8653), .ZN(n3484) );
  XNOR2_X1 U4706 ( .A(n4901), .B(n8654), .ZN(n3483) );
  NAND4_X1 U4707 ( .A1(n3486), .A2(n3485), .A3(n3484), .A4(n3483), .ZN(n3492)
         );
  XNOR2_X1 U4708 ( .A(n4900), .B(n8659), .ZN(n3490) );
  XNOR2_X1 U4709 ( .A(n4908), .B(n8652), .ZN(n3489) );
  XNOR2_X1 U4710 ( .A(n12195), .B(n8644), .ZN(n3488) );
  XNOR2_X1 U4711 ( .A(n6020), .B(n8633), .ZN(n3487) );
  NAND4_X1 U4712 ( .A1(n3490), .A2(n3489), .A3(n3488), .A4(n3487), .ZN(n3491)
         );
  NOR2_X1 U4713 ( .A1(n3492), .A2(n3491), .ZN(n3493) );
  NAND2_X1 U4714 ( .A1(pmp_addr_i[416]), .A2(pmp_addr_i[417]), .ZN(n11975) );
  AND2_X1 U4715 ( .A1(pmp_addr_i[420]), .A2(pmp_addr_i[419]), .ZN(n11954) );
  NAND4_X1 U4716 ( .A1(n3511), .A2(n11954), .A3(pmp_addr_i[421]), .A4(
        pmp_addr_i[422]), .ZN(n11988) );
  OR2_X1 U4717 ( .A1(n11988), .A2(n3549), .ZN(n11985) );
  OR2_X1 U4718 ( .A1(n11985), .A2(n3522), .ZN(n11989) );
  INV_X1 U4719 ( .A(pmp_cfg_i[107]), .ZN(n3536) );
  OAI21_X1 U4720 ( .B1(n11989), .B2(n3536), .A(pmp_cfg_i[108]), .ZN(n3523) );
  INV_X1 U4721 ( .A(pmp_addr_i[425]), .ZN(n3499) );
  NAND2_X1 U4722 ( .A1(n9911), .A2(pmp_addr_i[393]), .ZN(n3498) );
  OAI21_X1 U4723 ( .B1(n3523), .B2(n3499), .A(n3498), .ZN(n9819) );
  INV_X1 U4724 ( .A(n9819), .ZN(n9965) );
  NAND2_X1 U4725 ( .A1(n6002), .A2(n9965), .ZN(n4504) );
  OAI21_X1 U4726 ( .B1(n3535), .B2(n3536), .A(pmp_cfg_i[108]), .ZN(n3534) );
  INV_X1 U4727 ( .A(pmp_addr_i[428]), .ZN(n3501) );
  NAND2_X1 U4728 ( .A1(n9911), .A2(pmp_addr_i[396]), .ZN(n3500) );
  OAI21_X1 U4729 ( .B1(n3534), .B2(n3501), .A(n3500), .ZN(n9940) );
  INV_X1 U4730 ( .A(n9940), .ZN(n9988) );
  NAND2_X1 U4731 ( .A1(n11992), .A2(pmp_addr_i[426]), .ZN(n11952) );
  OR2_X1 U4732 ( .A1(n11952), .A2(n4582), .ZN(n11950) );
  AOI22_X1 U4733 ( .A1(n3503), .A2(n11989), .B1(n3502), .B2(n11950), .ZN(n3530) );
  INV_X1 U4734 ( .A(pmp_cfg_i[108]), .ZN(n3570) );
  NOR2_X1 U4735 ( .A1(n3570), .A2(pmp_cfg_i[107]), .ZN(n3574) );
  AOI21_X1 U4736 ( .B1(n11988), .B2(pmp_cfg_i[108]), .A(n3574), .ZN(n3550) );
  INV_X1 U4737 ( .A(pmp_addr_i[422]), .ZN(n3505) );
  NAND2_X1 U4738 ( .A1(n9911), .A2(pmp_addr_i[390]), .ZN(n3504) );
  OAI21_X1 U4739 ( .B1(n3550), .B2(n3505), .A(n3504), .ZN(n9798) );
  INV_X1 U4740 ( .A(n9798), .ZN(n9979) );
  AND2_X1 U4741 ( .A1(n5269), .A2(n9979), .ZN(n3561) );
  INV_X1 U4742 ( .A(pmp_addr_i[429]), .ZN(n3533) );
  OR2_X1 U4743 ( .A1(n3535), .A2(n3533), .ZN(n11963) );
  NAND2_X1 U4744 ( .A1(pmp_cfg_i[107]), .A2(pmp_cfg_i[108]), .ZN(n3515) );
  AOI21_X1 U4745 ( .B1(n11947), .B2(pmp_addr_i[431]), .A(n3515), .ZN(n3539) );
  NAND2_X1 U4746 ( .A1(n3539), .A2(n3511), .ZN(n11958) );
  INV_X1 U4747 ( .A(n11954), .ZN(n3506) );
  OR3_X1 U4748 ( .A1(n11958), .A2(n3506), .A3(n4604), .ZN(n11972) );
  NAND2_X1 U4749 ( .A1(n3533), .A2(pmp_cfg_i[108]), .ZN(n3508) );
  AOI21_X1 U4750 ( .B1(n3534), .B2(n3508), .A(n3507), .ZN(n3510) );
  AND2_X1 U4751 ( .A1(n9911), .A2(pmp_addr_i[398]), .ZN(n3509) );
  OR2_X1 U4752 ( .A1(n3510), .A2(n3509), .ZN(n11966) );
  INV_X1 U4753 ( .A(n11966), .ZN(n9986) );
  AND2_X1 U4754 ( .A1(n4743), .A2(n9986), .ZN(n3560) );
  AOI22_X1 U4755 ( .A1(n3561), .A2(n11972), .B1(n3560), .B2(n11963), .ZN(n3529) );
  INV_X1 U4756 ( .A(n9911), .ZN(n3629) );
  INV_X1 U4757 ( .A(n3574), .ZN(n9972) );
  OAI21_X1 U4758 ( .B1(n3511), .B2(n3570), .A(n9972), .ZN(n3524) );
  NAND2_X1 U4759 ( .A1(n3524), .A2(pmp_addr_i[419]), .ZN(n3512) );
  OAI21_X1 U4760 ( .B1(n3629), .B2(n3513), .A(n3512), .ZN(n9980) );
  INV_X1 U4761 ( .A(n9980), .ZN(n9971) );
  AND2_X1 U4762 ( .A1(n5293), .A2(n9971), .ZN(n3564) );
  OR2_X1 U4763 ( .A1(n12267), .A2(n3515), .ZN(n3520) );
  NOR2_X1 U4764 ( .A1(n11958), .A2(n3514), .ZN(n11969) );
  INV_X1 U4765 ( .A(n3515), .ZN(n11979) );
  NOR2_X1 U4766 ( .A1(n11954), .A2(n3570), .ZN(n3516) );
  OR2_X1 U4767 ( .A1(n3524), .A2(n3516), .ZN(n3551) );
  NAND2_X1 U4768 ( .A1(n3551), .A2(pmp_addr_i[421]), .ZN(n3517) );
  OAI21_X1 U4769 ( .B1(n3629), .B2(n3518), .A(n3517), .ZN(n9799) );
  AOI22_X1 U4770 ( .A1(n11969), .A2(pmp_addr_i[420]), .B1(n11979), .B2(n9799), 
        .ZN(n3519) );
  AOI22_X1 U4771 ( .A1(n3564), .A2(n11958), .B1(n3520), .B2(n3519), .ZN(n3528)
         );
  NAND2_X1 U4772 ( .A1(n9911), .A2(pmp_addr_i[392]), .ZN(n3521) );
  OAI21_X1 U4773 ( .B1(n3523), .B2(n3522), .A(n3521), .ZN(n9802) );
  INV_X1 U4774 ( .A(n9802), .ZN(n9966) );
  AND2_X1 U4775 ( .A1(n5262), .A2(n9966), .ZN(n3558) );
  NAND2_X1 U4776 ( .A1(n3524), .A2(pmp_addr_i[418]), .ZN(n3525) );
  OAI21_X1 U4777 ( .B1(n3629), .B2(n3526), .A(n3525), .ZN(n9787) );
  INV_X1 U4778 ( .A(n9787), .ZN(n9974) );
  AND2_X1 U4779 ( .A1(n12150), .A2(n9974), .ZN(n3563) );
  AOI22_X1 U4780 ( .A1(n3558), .A2(n11985), .B1(n3563), .B2(n11975), .ZN(n3527) );
  NAND4_X1 U4781 ( .A1(n3530), .A2(n3529), .A3(n3528), .A4(n3527), .ZN(n3569)
         );
  INV_X1 U4782 ( .A(n207), .ZN(n4498) );
  NAND2_X1 U4783 ( .A1(n9911), .A2(pmp_addr_i[397]), .ZN(n3532) );
  OAI21_X1 U4784 ( .B1(n3534), .B2(n3533), .A(n3532), .ZN(n9942) );
  INV_X1 U4785 ( .A(n9942), .ZN(n4497) );
  INV_X1 U4786 ( .A(n3535), .ZN(n11990) );
  OAI21_X1 U4787 ( .B1(n11952), .B2(n3536), .A(pmp_cfg_i[108]), .ZN(n3545) );
  NAND2_X1 U4788 ( .A1(n9911), .A2(pmp_addr_i[394]), .ZN(n3537) );
  OAI21_X1 U4789 ( .B1(n3545), .B2(n3538), .A(n3537), .ZN(n9948) );
  NOR2_X1 U4790 ( .A1(n9948), .A2(n11992), .ZN(n3543) );
  NAND2_X1 U4791 ( .A1(n3626), .A2(pmp_addr_i[431]), .ZN(n3540) );
  OAI21_X1 U4792 ( .B1(n3629), .B2(n3541), .A(n3540), .ZN(n9842) );
  NOR2_X1 U4793 ( .A1(n9842), .A2(n11947), .ZN(n3542) );
  AOI22_X1 U4794 ( .A1(instr_addr_o_12_), .A2(n3543), .B1(n12265), .B2(n3542), 
        .ZN(n3547) );
  NAND2_X1 U4795 ( .A1(n9911), .A2(pmp_addr_i[395]), .ZN(n3544) );
  OAI21_X1 U4796 ( .B1(n3545), .B2(n4582), .A(n3544), .ZN(n9946) );
  INV_X1 U4797 ( .A(n9946), .ZN(n9982) );
  NAND3_X1 U4798 ( .A1(instr_addr_o_13_), .A2(n9982), .A3(n11952), .ZN(n3546)
         );
  OAI211_X1 U4799 ( .C1(n4514), .C2(n11990), .A(n3547), .B(n3546), .ZN(n3557)
         );
  INV_X1 U4800 ( .A(n11988), .ZN(n3555) );
  NAND2_X1 U4801 ( .A1(n9911), .A2(pmp_addr_i[391]), .ZN(n3548) );
  OAI21_X1 U4802 ( .B1(n3550), .B2(n3549), .A(n3548), .ZN(n9801) );
  INV_X1 U4803 ( .A(n9801), .ZN(n9978) );
  NAND2_X1 U4804 ( .A1(n3551), .A2(pmp_addr_i[420]), .ZN(n3552) );
  OAI21_X1 U4805 ( .B1(n3629), .B2(n3553), .A(n3552), .ZN(n9790) );
  INV_X1 U4806 ( .A(n9790), .ZN(n3554) );
  NAND2_X1 U4807 ( .A1(n5277), .A2(n3554), .ZN(n4473) );
  OAI22_X1 U4808 ( .A1(n3555), .A2(n4484), .B1(n4473), .B2(n11969), .ZN(n3556)
         );
  OR2_X1 U4809 ( .A1(n3557), .A2(n3556), .ZN(n3568) );
  NAND2_X1 U4810 ( .A1(n937), .A2(n9982), .ZN(n4507) );
  INV_X1 U4811 ( .A(n4507), .ZN(n3559) );
  INV_X1 U4812 ( .A(n9799), .ZN(n4476) );
  NAND2_X1 U4813 ( .A1(n5740), .A2(n4476), .ZN(n4481) );
  INV_X1 U4814 ( .A(n9948), .ZN(n9983) );
  NAND2_X1 U4815 ( .A1(n4494), .A2(n9983), .ZN(n4503) );
  NAND4_X1 U4816 ( .A1(n4481), .A2(n4470), .A3(n4474), .A4(n4503), .ZN(n3565)
         );
  NOR2_X1 U4817 ( .A1(n3566), .A2(n3565), .ZN(n3567) );
  NOR2_X1 U4818 ( .A1(n4204), .A2(n9978), .ZN(n4478) );
  NOR2_X1 U4819 ( .A1(n3570), .A2(pmp_addr_i[416]), .ZN(n3571) );
  OAI21_X1 U4820 ( .B1(n3574), .B2(n3571), .A(pmp_addr_i[417]), .ZN(n3573) );
  NAND2_X1 U4821 ( .A1(n9911), .A2(pmp_addr_i[385]), .ZN(n3572) );
  NAND2_X1 U4822 ( .A1(n3573), .A2(n3572), .ZN(n9784) );
  NAND2_X1 U4823 ( .A1(n9911), .A2(pmp_addr_i[384]), .ZN(n3576) );
  NAND2_X1 U4824 ( .A1(n3574), .A2(pmp_addr_i[416]), .ZN(n3575) );
  NAND2_X1 U4825 ( .A1(n3576), .A2(n3575), .ZN(n9783) );
  INV_X1 U4826 ( .A(pmp_cfg_i[106]), .ZN(n3577) );
  NOR3_X1 U4827 ( .A1(n9784), .A2(n9783), .A3(n3577), .ZN(n3578) );
  OR2_X1 U4828 ( .A1(n3626), .A2(n9911), .ZN(n9994) );
  OAI211_X1 U4829 ( .C1(n6015), .C2(n9971), .A(n3578), .B(n9994), .ZN(n3579)
         );
  NOR2_X1 U4830 ( .A1(n4478), .A2(n3579), .ZN(n3587) );
  NAND2_X1 U4831 ( .A1(n3626), .A2(pmp_addr_i[435]), .ZN(n3580) );
  OAI21_X1 U4832 ( .B1(n3629), .B2(n3581), .A(n3580), .ZN(n9914) );
  XNOR2_X1 U4833 ( .A(n5842), .B(n9914), .ZN(n3586) );
  NAND2_X1 U4834 ( .A1(n3626), .A2(pmp_addr_i[433]), .ZN(n3582) );
  OAI21_X1 U4835 ( .B1(n3629), .B2(n3583), .A(n3582), .ZN(n9934) );
  XNOR2_X1 U4836 ( .A(n6020), .B(n9934), .ZN(n3585) );
  NAND2_X1 U4837 ( .A1(n3626), .A2(pmp_addr_i[445]), .ZN(n12006) );
  OAI21_X1 U4838 ( .B1(n3629), .B2(n12085), .A(n12006), .ZN(n9964) );
  XNOR2_X1 U4839 ( .A(n4866), .B(n9964), .ZN(n3584) );
  NAND4_X1 U4840 ( .A1(n3587), .A2(n3586), .A3(n3585), .A4(n3584), .ZN(n3599)
         );
  NAND2_X1 U4841 ( .A1(n3626), .A2(pmp_addr_i[432]), .ZN(n3588) );
  OAI21_X1 U4842 ( .B1(n3629), .B2(n3589), .A(n3588), .ZN(n9939) );
  XNOR2_X1 U4843 ( .A(n4908), .B(n9939), .ZN(n3597) );
  NAND2_X1 U4844 ( .A1(n3626), .A2(pmp_addr_i[440]), .ZN(n3590) );
  OAI21_X1 U4845 ( .B1(n3629), .B2(n3591), .A(n3590), .ZN(n9925) );
  XNOR2_X1 U4846 ( .A(n5985), .B(n9925), .ZN(n3596) );
  NAND2_X1 U4847 ( .A1(n3626), .A2(pmp_addr_i[444]), .ZN(n3592) );
  OAI21_X1 U4848 ( .B1(n3629), .B2(n1598), .A(n3592), .ZN(n9957) );
  XNOR2_X1 U4849 ( .A(n12207), .B(n9957), .ZN(n3595) );
  NAND2_X1 U4850 ( .A1(n3626), .A2(pmp_addr_i[443]), .ZN(n3593) );
  OAI21_X1 U4851 ( .B1(n3629), .B2(n1631), .A(n3593), .ZN(n9956) );
  XNOR2_X1 U4852 ( .A(n5550), .B(n9956), .ZN(n3594) );
  NAND4_X1 U4853 ( .A1(n3597), .A2(n3596), .A3(n3595), .A4(n3594), .ZN(n3598)
         );
  NOR2_X1 U4854 ( .A1(n3599), .A2(n3598), .ZN(n3637) );
  NAND2_X1 U4855 ( .A1(n3626), .A2(pmp_addr_i[437]), .ZN(n3600) );
  OAI21_X1 U4856 ( .B1(n3629), .B2(n3601), .A(n3600), .ZN(n9917) );
  XNOR2_X1 U4857 ( .A(n6025), .B(n9917), .ZN(n3611) );
  NAND2_X1 U4858 ( .A1(n3626), .A2(pmp_addr_i[436]), .ZN(n3602) );
  OAI21_X1 U4859 ( .B1(n3629), .B2(n3603), .A(n3602), .ZN(n9916) );
  XNOR2_X1 U4860 ( .A(n12157), .B(n9916), .ZN(n3610) );
  NAND2_X1 U4861 ( .A1(n3626), .A2(pmp_addr_i[438]), .ZN(n3604) );
  OAI21_X1 U4862 ( .B1(n3629), .B2(n3605), .A(n3604), .ZN(n9918) );
  XNOR2_X1 U4863 ( .A(n4835), .B(n9918), .ZN(n3609) );
  NAND2_X1 U4864 ( .A1(n3626), .A2(pmp_addr_i[434]), .ZN(n3606) );
  OAI21_X1 U4865 ( .B1(n3629), .B2(n3607), .A(n3606), .ZN(n9936) );
  XNOR2_X1 U4866 ( .A(instr_addr_o_20_), .B(n9936), .ZN(n3608) );
  AND4_X1 U4867 ( .A1(n3611), .A2(n3610), .A3(n3609), .A4(n3608), .ZN(n3618)
         );
  OAI22_X1 U4868 ( .A1(n6002), .A2(n9965), .B1(n12180), .B2(n9988), .ZN(n3613)
         );
  OAI22_X1 U4869 ( .A1(n205), .A2(n9979), .B1(n5229), .B2(n9986), .ZN(n3612)
         );
  NOR2_X1 U4870 ( .A1(n3613), .A2(n3612), .ZN(n3617) );
  OAI22_X1 U4871 ( .A1(n5997), .A2(n9982), .B1(n12179), .B2(n4497), .ZN(n3615)
         );
  OAI22_X1 U4872 ( .A1(instr_addr_o_6_), .A2(n3554), .B1(n12267), .B2(n4476), 
        .ZN(n3614) );
  NOR2_X1 U4873 ( .A1(n3615), .A2(n3614), .ZN(n3616) );
  NAND3_X1 U4874 ( .A1(n3617), .A2(n3618), .A3(n3616), .ZN(n3635) );
  INV_X1 U4875 ( .A(n9842), .ZN(n4516) );
  OAI22_X1 U4876 ( .A1(instr_addr_o_12_), .A2(n9983), .B1(n5974), .B2(n4516), 
        .ZN(n3621) );
  OAI22_X1 U4877 ( .A1(n12202), .A2(n9966), .B1(n5976), .B2(n9974), .ZN(n3620)
         );
  NOR2_X1 U4878 ( .A1(n3621), .A2(n3620), .ZN(n3633) );
  NAND2_X1 U4879 ( .A1(n3626), .A2(pmp_addr_i[442]), .ZN(n3622) );
  OAI21_X1 U4880 ( .B1(n3629), .B2(n3623), .A(n3622), .ZN(n9927) );
  XNOR2_X1 U4881 ( .A(n4901), .B(n9927), .ZN(n3632) );
  NAND2_X1 U4882 ( .A1(n3626), .A2(pmp_addr_i[441]), .ZN(n3624) );
  OAI21_X1 U4883 ( .B1(n3629), .B2(n3625), .A(n3624), .ZN(n9926) );
  XNOR2_X1 U4884 ( .A(instr_addr_o_27_), .B(n9926), .ZN(n3631) );
  NAND2_X1 U4885 ( .A1(n3626), .A2(pmp_addr_i[439]), .ZN(n3627) );
  OAI21_X1 U4886 ( .B1(n3629), .B2(n3628), .A(n3627), .ZN(n9924) );
  XNOR2_X1 U4887 ( .A(n12226), .B(n9924), .ZN(n3630) );
  NAND4_X1 U4888 ( .A1(n3633), .A2(n3632), .A3(n3631), .A4(n3630), .ZN(n3634)
         );
  NOR2_X1 U4889 ( .A1(n3635), .A2(n3634), .ZN(n3636) );
  NAND2_X1 U4891 ( .A1(pmp_privil_mode_i[1]), .A2(pmp_privil_mode_i[0]), .ZN(
        n8081) );
  NAND2_X1 U4892 ( .A1(pmp_addr_i[0]), .A2(pmp_addr_i[1]), .ZN(n3691) );
  INV_X1 U4893 ( .A(pmp_addr_i[2]), .ZN(n3690) );
  OR2_X1 U4894 ( .A1(n3691), .A2(n3690), .ZN(n3642) );
  NAND2_X1 U4895 ( .A1(pmp_cfg_i[3]), .A2(pmp_addr_i[3]), .ZN(n3639) );
  NOR2_X1 U4896 ( .A1(n3642), .A2(n3639), .ZN(n3675) );
  NAND2_X1 U4897 ( .A1(pmp_addr_i[4]), .A2(pmp_addr_i[5]), .ZN(n3674) );
  NAND2_X1 U4898 ( .A1(pmp_addr_i[6]), .A2(pmp_addr_i[7]), .ZN(n3640) );
  NOR2_X1 U4899 ( .A1(n3674), .A2(n3640), .ZN(n3643) );
  NAND2_X1 U4900 ( .A1(n3675), .A2(n3643), .ZN(n3665) );
  INV_X1 U4901 ( .A(pmp_addr_i[8]), .ZN(n3641) );
  NOR2_X1 U4902 ( .A1(n3665), .A2(n3641), .ZN(n3672) );
  NAND2_X1 U4903 ( .A1(n3672), .A2(pmp_addr_i[9]), .ZN(n3684) );
  NAND2_X1 U4904 ( .A1(pmp_addr_i[10]), .A2(pmp_addr_i[11]), .ZN(n3645) );
  NOR2_X1 U4905 ( .A1(n3684), .A2(n3645), .ZN(n3661) );
  INV_X1 U4906 ( .A(pmp_addr_i[11]), .ZN(n3652) );
  INV_X1 U4907 ( .A(n3642), .ZN(n3663) );
  NAND4_X1 U4908 ( .A1(n3663), .A2(pmp_addr_i[3]), .A3(pmp_addr_i[8]), .A4(
        n3643), .ZN(n3648) );
  NAND2_X1 U4909 ( .A1(pmp_addr_i[13]), .A2(pmp_addr_i[12]), .ZN(n3644) );
  OR2_X1 U4910 ( .A1(n3645), .A2(n3644), .ZN(n3650) );
  INV_X1 U4911 ( .A(n3650), .ZN(n3646) );
  NAND4_X1 U4912 ( .A1(n3646), .A2(pmp_addr_i[15]), .A3(pmp_addr_i[14]), .A4(
        pmp_addr_i[9]), .ZN(n3647) );
  AND2_X1 U4913 ( .A1(pmp_cfg_i[3]), .A2(pmp_cfg_i[4]), .ZN(n11230) );
  OAI21_X1 U4914 ( .B1(n3648), .B2(n3647), .A(n11230), .ZN(n3688) );
  OR2_X1 U4915 ( .A1(n3688), .A2(n3648), .ZN(n11206) );
  INV_X1 U4916 ( .A(pmp_addr_i[9]), .ZN(n3649) );
  NOR2_X1 U4917 ( .A1(n11206), .A2(n3649), .ZN(n11210) );
  NAND2_X1 U4918 ( .A1(n11210), .A2(pmp_addr_i[10]), .ZN(n11215) );
  NAND3_X1 U4919 ( .A1(instr_addr_o_13_), .A2(n330), .A3(n11215), .ZN(n3659)
         );
  NOR2_X1 U4920 ( .A1(n3684), .A2(n3650), .ZN(n3683) );
  INV_X1 U4921 ( .A(pmp_addr_i[13]), .ZN(n3651) );
  NOR2_X1 U4922 ( .A1(n11215), .A2(n3652), .ZN(n11209) );
  NAND2_X1 U4923 ( .A1(n11209), .A2(pmp_addr_i[12]), .ZN(n3682) );
  NAND3_X1 U4924 ( .A1(instr_addr_o_15_), .A2(n329), .A3(n3682), .ZN(n3658) );
  NAND2_X1 U4925 ( .A1(n3663), .A2(pmp_addr_i[3]), .ZN(n3653) );
  OR2_X1 U4926 ( .A1(n3688), .A2(n3653), .ZN(n11234) );
  INV_X1 U4927 ( .A(pmp_addr_i[4]), .ZN(n3654) );
  NOR2_X1 U4928 ( .A1(n11234), .A2(n3654), .ZN(n11218) );
  NAND2_X1 U4929 ( .A1(n11218), .A2(pmp_addr_i[5]), .ZN(n11220) );
  OR2_X1 U4930 ( .A1(n11220), .A2(n3655), .ZN(n11207) );
  NAND3_X1 U4931 ( .A1(n155), .A2(n158), .A3(n11207), .ZN(n3657) );
  NAND3_X1 U4932 ( .A1(instr_addr_o_6_), .A2(n324), .A3(n11234), .ZN(n3656) );
  AND4_X1 U4933 ( .A1(n3659), .A2(n3658), .A3(n3657), .A4(n3656), .ZN(n3671)
         );
  INV_X1 U4934 ( .A(pmp_addr_i[12]), .ZN(n3660) );
  NOR2_X1 U4935 ( .A1(n3661), .A2(n3660), .ZN(n11333) );
  INV_X1 U4936 ( .A(n11333), .ZN(n11208) );
  OAI22_X1 U4937 ( .A1(n5997), .A2(n330), .B1(n12181), .B2(n11208), .ZN(n3708)
         );
  INV_X1 U4938 ( .A(n3708), .ZN(n3670) );
  INV_X1 U4939 ( .A(pmp_addr_i[3]), .ZN(n3662) );
  NOR2_X1 U4940 ( .A1(n3675), .A2(n3662), .ZN(n11290) );
  NOR2_X1 U4941 ( .A1(n11290), .A2(n3663), .ZN(n11233) );
  INV_X1 U4942 ( .A(n11230), .ZN(n3664) );
  AOI21_X1 U4943 ( .B1(n6015), .B2(n11233), .A(n3664), .ZN(n3669) );
  AND2_X1 U4944 ( .A1(n3665), .A2(pmp_addr_i[8]), .ZN(n11213) );
  INV_X1 U4945 ( .A(pmp_addr_i[7]), .ZN(n3666) );
  NOR2_X1 U4946 ( .A1(n11207), .A2(n3666), .ZN(n11214) );
  OAI21_X1 U4947 ( .B1(n11213), .B2(n11214), .A(n12202), .ZN(n3667) );
  OAI21_X1 U4948 ( .B1(n12202), .B2(n11213), .A(n3667), .ZN(n3668) );
  NAND4_X1 U4949 ( .A1(n3671), .A2(n3670), .A3(n3669), .A4(n3668), .ZN(n3715)
         );
  NOR2_X1 U4950 ( .A1(n3672), .A2(n3649), .ZN(n3698) );
  INV_X1 U4951 ( .A(n11206), .ZN(n3673) );
  NOR2_X1 U4952 ( .A1(n3698), .A2(n3673), .ZN(n3678) );
  INV_X1 U4953 ( .A(n3674), .ZN(n3676) );
  NAND2_X1 U4954 ( .A1(n3676), .A2(n3675), .ZN(n3679) );
  AND2_X1 U4955 ( .A1(n3679), .A2(pmp_addr_i[5]), .ZN(n3699) );
  NOR2_X1 U4956 ( .A1(n11218), .A2(n3699), .ZN(n3677) );
  AOI22_X1 U4957 ( .A1(n3934), .A2(n3678), .B1(n4605), .B2(n3677), .ZN(n3697)
         );
  NOR2_X1 U4958 ( .A1(n11209), .A2(n11333), .ZN(n3681) );
  AND2_X1 U4959 ( .A1(n11220), .A2(n159), .ZN(n3680) );
  AOI22_X1 U4960 ( .A1(n12181), .A2(n3681), .B1(n6005), .B2(n3680), .ZN(n3696)
         );
  INV_X1 U4961 ( .A(n3682), .ZN(n11237) );
  NAND2_X1 U4962 ( .A1(n11237), .A2(pmp_addr_i[13]), .ZN(n11226) );
  INV_X1 U4963 ( .A(pmp_addr_i[14]), .ZN(n3687) );
  AND2_X1 U4964 ( .A1(n11226), .A2(n328), .ZN(n3686) );
  AND2_X1 U4965 ( .A1(n3684), .A2(pmp_addr_i[10]), .ZN(n3700) );
  NOR2_X1 U4966 ( .A1(n3700), .A2(n11210), .ZN(n3685) );
  AOI22_X1 U4967 ( .A1(n12203), .A2(n3686), .B1(n5245), .B2(n3685), .ZN(n3695)
         );
  NOR2_X1 U4968 ( .A1(n11226), .A2(n3687), .ZN(n11241) );
  INV_X1 U4969 ( .A(pmp_cfg_i[4]), .ZN(n3865) );
  OR2_X1 U4970 ( .A1(n3865), .A2(pmp_cfg_i[3]), .ZN(n11250) );
  NAND2_X1 U4971 ( .A1(n3688), .A2(n11250), .ZN(n3745) );
  INV_X1 U4972 ( .A(pmp_cfg_i[3]), .ZN(n3689) );
  NOR2_X1 U4973 ( .A1(n3689), .A2(pmp_cfg_i[4]), .ZN(n8079) );
  AND2_X1 U4974 ( .A1(n3758), .A2(pmp_addr_i[15]), .ZN(n7994) );
  NOR2_X1 U4975 ( .A1(n11241), .A2(n7994), .ZN(n3693) );
  NOR2_X1 U4976 ( .A1(n3691), .A2(n3689), .ZN(n3735) );
  NOR2_X1 U4977 ( .A1(n3735), .A2(n3690), .ZN(n3732) );
  INV_X1 U4978 ( .A(n3691), .ZN(n3692) );
  NOR2_X1 U4979 ( .A1(n3732), .A2(n3692), .ZN(n11229) );
  AOI22_X1 U4980 ( .A1(n5062), .A2(n3693), .B1(n5899), .B2(n11229), .ZN(n3694)
         );
  NAND4_X1 U4981 ( .A1(n3697), .A2(n3696), .A3(n3695), .A4(n3694), .ZN(n3714)
         );
  INV_X1 U4982 ( .A(n3698), .ZN(n11335) );
  INV_X1 U4983 ( .A(n3699), .ZN(n11345) );
  AOI22_X1 U4984 ( .A1(n6002), .A2(n11335), .B1(n5740), .B2(n11345), .ZN(n3704) );
  AOI22_X1 U4985 ( .A1(instr_addr_o_9_), .A2(n158), .B1(instr_addr_o_6_), .B2(
        n324), .ZN(n3703) );
  AOI22_X1 U4986 ( .A1(n12181), .A2(n11208), .B1(n6005), .B2(n159), .ZN(n3702)
         );
  INV_X1 U4987 ( .A(n3700), .ZN(n11336) );
  AOI22_X1 U4988 ( .A1(n5229), .A2(n328), .B1(n5245), .B2(n11336), .ZN(n3701)
         );
  AND4_X1 U4989 ( .A1(n3703), .A2(n3702), .A3(n3704), .A4(n3701), .ZN(n3712)
         );
  AOI22_X1 U4990 ( .A1(n5997), .A2(n330), .B1(n12179), .B2(n329), .ZN(n3711)
         );
  INV_X1 U4991 ( .A(n11290), .ZN(n11254) );
  AOI21_X1 U4992 ( .B1(n6015), .B2(n11254), .A(n11250), .ZN(n3706) );
  INV_X1 U4993 ( .A(n7994), .ZN(n3733) );
  NAND2_X1 U4994 ( .A1(n5974), .A2(n3733), .ZN(n3705) );
  OAI211_X1 U4995 ( .C1(n3876), .C2(n3732), .A(n3706), .B(n3705), .ZN(n3707)
         );
  NOR2_X1 U4996 ( .A1(n3708), .A2(n3707), .ZN(n3710) );
  XNOR2_X1 U4997 ( .A(n12202), .B(n11213), .ZN(n3709) );
  NAND4_X1 U4998 ( .A1(n3712), .A2(n3711), .A3(n3710), .A4(n3709), .ZN(n3713)
         );
  OAI21_X1 U4999 ( .B1(n3715), .B2(n3714), .A(n3713), .ZN(n3753) );
  XNOR2_X1 U5000 ( .A(instr_addr_o_21_), .B(pmp_addr_i[19]), .ZN(n3719) );
  XNOR2_X1 U5001 ( .A(n5985), .B(pmp_addr_i[24]), .ZN(n3718) );
  AND2_X1 U5002 ( .A1(n3745), .A2(pmp_addr_i[16]), .ZN(n11297) );
  XNOR2_X1 U5003 ( .A(n4908), .B(n11297), .ZN(n3717) );
  XNOR2_X1 U5004 ( .A(n5550), .B(pmp_addr_i[27]), .ZN(n3716) );
  NAND4_X1 U5005 ( .A1(n3719), .A2(n3718), .A3(n3717), .A4(n3716), .ZN(n3725)
         );
  AND2_X1 U5006 ( .A1(n3745), .A2(pmp_addr_i[17]), .ZN(n11282) );
  XNOR2_X1 U5007 ( .A(n6020), .B(n11282), .ZN(n3723) );
  XNOR2_X1 U5008 ( .A(n4866), .B(pmp_addr_i[29]), .ZN(n3722) );
  AND2_X1 U5009 ( .A1(n3745), .A2(pmp_addr_i[21]), .ZN(n11295) );
  XNOR2_X1 U5010 ( .A(n6025), .B(n11295), .ZN(n3721) );
  XNOR2_X1 U5011 ( .A(n12213), .B(pmp_addr_i[20]), .ZN(n3720) );
  NAND4_X1 U5012 ( .A1(n3723), .A2(n3722), .A3(n3721), .A4(n3720), .ZN(n3724)
         );
  NOR2_X1 U5013 ( .A1(n3725), .A2(n3724), .ZN(n3752) );
  OAI22_X1 U5014 ( .A1(n155), .A2(n158), .B1(n12179), .B2(n329), .ZN(n3727) );
  OAI22_X1 U5015 ( .A1(instr_addr_o_6_), .A2(n324), .B1(n4605), .B2(n11345), 
        .ZN(n3726) );
  NOR2_X1 U5016 ( .A1(n3727), .A2(n3726), .ZN(n3744) );
  OAI22_X1 U5017 ( .A1(n6002), .A2(n11335), .B1(n6005), .B2(n159), .ZN(n3729)
         );
  OAI22_X1 U5018 ( .A1(n5226), .A2(n328), .B1(n5245), .B2(n11336), .ZN(n3728)
         );
  NOR2_X1 U5019 ( .A1(n3729), .A2(n3728), .ZN(n3743) );
  AND2_X1 U5020 ( .A1(n3745), .A2(pmp_addr_i[18]), .ZN(n11284) );
  XNOR2_X1 U5021 ( .A(instr_addr_o_20_), .B(n11284), .ZN(n3731) );
  XNOR2_X1 U5022 ( .A(n4835), .B(pmp_addr_i[22]), .ZN(n3730) );
  AND2_X1 U5023 ( .A1(n3731), .A2(n3730), .ZN(n3742) );
  INV_X1 U5024 ( .A(n3732), .ZN(n11287) );
  OAI22_X1 U5025 ( .A1(n12265), .A2(n3733), .B1(n5976), .B2(n11287), .ZN(n3740) );
  INV_X1 U5026 ( .A(pmp_addr_i[1]), .ZN(n3734) );
  NOR2_X1 U5027 ( .A1(n3735), .A2(n3734), .ZN(n11228) );
  INV_X1 U5028 ( .A(pmp_addr_i[0]), .ZN(n11258) );
  NOR2_X1 U5029 ( .A1(n11250), .A2(n11258), .ZN(n3737) );
  INV_X1 U5030 ( .A(pmp_cfg_i[2]), .ZN(n3736) );
  NOR3_X1 U5031 ( .A1(n11228), .A2(n3737), .A3(n3736), .ZN(n3738) );
  OAI211_X1 U5032 ( .C1(n6015), .C2(n11254), .A(n3738), .B(n3758), .ZN(n3739)
         );
  NOR2_X1 U5033 ( .A1(n3740), .A2(n3739), .ZN(n3741) );
  NAND4_X1 U5034 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3751)
         );
  XNOR2_X1 U5035 ( .A(n12226), .B(pmp_addr_i[23]), .ZN(n3749) );
  AND2_X1 U5036 ( .A1(n3745), .A2(pmp_addr_i[26]), .ZN(n11318) );
  XNOR2_X1 U5037 ( .A(n4901), .B(n11318), .ZN(n3748) );
  AND2_X1 U5038 ( .A1(n3745), .A2(pmp_addr_i[28]), .ZN(n11304) );
  XNOR2_X1 U5039 ( .A(n4753), .B(n11304), .ZN(n3747) );
  AND2_X1 U5040 ( .A1(n3745), .A2(pmp_addr_i[25]), .ZN(n11321) );
  XNOR2_X1 U5041 ( .A(instr_addr_o_27_), .B(n11321), .ZN(n3746) );
  NAND4_X1 U5042 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .ZN(n3750)
         );
  AND2_X1 U5043 ( .A1(n3758), .A2(pmp_addr_i[16]), .ZN(n7996) );
  INV_X1 U5044 ( .A(n7996), .ZN(n3759) );
  NAND2_X1 U5045 ( .A1(n6019), .A2(n3759), .ZN(n3776) );
  OAI21_X1 U5046 ( .B1(n4234), .B2(n7994), .A(n3776), .ZN(n3778) );
  AND2_X1 U5047 ( .A1(n3758), .A2(pmp_addr_i[13]), .ZN(n7988) );
  AND2_X1 U5048 ( .A1(n3758), .A2(pmp_addr_i[14]), .ZN(n7989) );
  INV_X1 U5049 ( .A(n7989), .ZN(n3760) );
  NAND2_X1 U5050 ( .A1(n5229), .A2(n3760), .ZN(n3774) );
  OAI21_X1 U5051 ( .B1(n4578), .B2(n7988), .A(n3774), .ZN(n3761) );
  NOR2_X1 U5052 ( .A1(n3778), .A2(n3761), .ZN(n3859) );
  AND2_X1 U5053 ( .A1(n3758), .A2(pmp_addr_i[10]), .ZN(n7975) );
  INV_X1 U5054 ( .A(n7975), .ZN(n3762) );
  NAND2_X1 U5055 ( .A1(instr_addr_o_12_), .A2(n3762), .ZN(n3855) );
  AND2_X1 U5056 ( .A1(n3758), .A2(pmp_addr_i[9]), .ZN(n7974) );
  INV_X1 U5057 ( .A(n7974), .ZN(n3763) );
  NOR2_X1 U5058 ( .A1(n3934), .A2(n3763), .ZN(n3764) );
  AOI22_X1 U5059 ( .A1(n3855), .A2(n3764), .B1(n5070), .B2(n7975), .ZN(n3771)
         );
  AND2_X1 U5060 ( .A1(n3758), .A2(pmp_addr_i[12]), .ZN(n7981) );
  INV_X1 U5061 ( .A(n7981), .ZN(n3765) );
  NAND2_X1 U5062 ( .A1(instr_addr_o_14_), .A2(n3765), .ZN(n3769) );
  AND2_X1 U5063 ( .A1(n3758), .A2(pmp_addr_i[11]), .ZN(n7980) );
  INV_X1 U5064 ( .A(n7980), .ZN(n3767) );
  NAND2_X1 U5065 ( .A1(n4061), .A2(n3767), .ZN(n3766) );
  NAND2_X1 U5066 ( .A1(n3769), .A2(n3766), .ZN(n3857) );
  NOR2_X1 U5067 ( .A1(n149), .A2(n3767), .ZN(n3768) );
  AOI22_X1 U5068 ( .A1(n3769), .A2(n3768), .B1(instr_addr_o_14__BAR), .B2(
        n7981), .ZN(n3770) );
  OAI21_X1 U5069 ( .B1(n3771), .B2(n3857), .A(n3770), .ZN(n3781) );
  INV_X1 U5070 ( .A(n7988), .ZN(n3772) );
  NOR2_X1 U5071 ( .A1(instr_addr_o_15_), .A2(n3772), .ZN(n3773) );
  AOI22_X1 U5072 ( .A1(n3774), .A2(n3773), .B1(n5058), .B2(n7989), .ZN(n3779)
         );
  NOR2_X1 U5073 ( .A1(n4069), .A2(n3733), .ZN(n3775) );
  AOI22_X1 U5074 ( .A1(n3776), .A2(n3775), .B1(n2082), .B2(n7996), .ZN(n3777)
         );
  OAI21_X1 U5075 ( .B1(n3779), .B2(n3778), .A(n3777), .ZN(n3780) );
  AOI21_X1 U5076 ( .B1(n3859), .B2(n3781), .A(n3780), .ZN(n3828) );
  AND2_X1 U5077 ( .A1(n3758), .A2(pmp_addr_i[27]), .ZN(n8054) );
  AND2_X1 U5078 ( .A1(n3758), .A2(pmp_addr_i[28]), .ZN(n8055) );
  INV_X1 U5079 ( .A(n8055), .ZN(n3782) );
  NAND2_X1 U5080 ( .A1(n12263), .A2(n3782), .ZN(n3799) );
  OAI21_X1 U5081 ( .B1(n4656), .B2(n8054), .A(n3799), .ZN(n3798) );
  AND2_X1 U5082 ( .A1(n3758), .A2(pmp_addr_i[26]), .ZN(n8050) );
  INV_X1 U5083 ( .A(n8050), .ZN(n3783) );
  NAND2_X1 U5084 ( .A1(instr_addr_o_28_), .A2(n3783), .ZN(n3796) );
  AND2_X1 U5085 ( .A1(n3758), .A2(pmp_addr_i[29]), .ZN(n8062) );
  INV_X1 U5086 ( .A(n8062), .ZN(n3784) );
  NAND2_X1 U5087 ( .A1(n191), .A2(n3784), .ZN(n3800) );
  AND2_X1 U5088 ( .A1(n3758), .A2(pmp_addr_i[25]), .ZN(n8049) );
  INV_X1 U5089 ( .A(n8049), .ZN(n3785) );
  NAND2_X1 U5090 ( .A1(n12195), .A2(n3785), .ZN(n3786) );
  NAND3_X1 U5091 ( .A1(n3796), .A2(n3800), .A3(n3786), .ZN(n3787) );
  NOR2_X1 U5092 ( .A1(n3798), .A2(n3787), .ZN(n3825) );
  AND2_X1 U5093 ( .A1(n3758), .A2(pmp_addr_i[23]), .ZN(n8038) );
  AND2_X1 U5094 ( .A1(n3758), .A2(pmp_addr_i[24]), .ZN(n8039) );
  INV_X1 U5095 ( .A(n8039), .ZN(n3788) );
  NAND2_X1 U5096 ( .A1(n12158), .A2(n3788), .ZN(n3808) );
  OAI21_X1 U5097 ( .B1(n135), .B2(n8038), .A(n3808), .ZN(n3810) );
  AND2_X1 U5098 ( .A1(n3758), .A2(pmp_addr_i[21]), .ZN(n8033) );
  AND2_X1 U5099 ( .A1(n3758), .A2(pmp_addr_i[22]), .ZN(n8034) );
  INV_X1 U5100 ( .A(n8034), .ZN(n3789) );
  NAND2_X1 U5101 ( .A1(n6028), .A2(n3789), .ZN(n3804) );
  OAI21_X1 U5102 ( .B1(n5086), .B2(n8033), .A(n3804), .ZN(n3790) );
  NOR2_X1 U5103 ( .A1(n3810), .A2(n3790), .ZN(n3824) );
  AND2_X1 U5104 ( .A1(n3758), .A2(pmp_addr_i[19]), .ZN(n8025) );
  INV_X1 U5105 ( .A(n8025), .ZN(n3791) );
  NAND2_X1 U5106 ( .A1(instr_addr_o_21_), .A2(n3791), .ZN(n3817) );
  AND2_X1 U5107 ( .A1(n3758), .A2(pmp_addr_i[20]), .ZN(n8026) );
  INV_X1 U5108 ( .A(n8026), .ZN(n3792) );
  NAND2_X1 U5109 ( .A1(n4836), .A2(n3792), .ZN(n3818) );
  AND2_X1 U5110 ( .A1(n3758), .A2(pmp_addr_i[18]), .ZN(n8021) );
  INV_X1 U5111 ( .A(n8021), .ZN(n3813) );
  NAND2_X1 U5112 ( .A1(instr_addr_o_20_), .A2(n3813), .ZN(n3815) );
  AND2_X1 U5113 ( .A1(n3758), .A2(pmp_addr_i[17]), .ZN(n8020) );
  INV_X1 U5114 ( .A(n8020), .ZN(n3814) );
  NAND2_X1 U5115 ( .A1(instr_addr_o_19_), .A2(n3814), .ZN(n3794) );
  AND4_X1 U5116 ( .A1(n3817), .A2(n3818), .A3(n3815), .A4(n3794), .ZN(n3795)
         );
  NAND3_X1 U5117 ( .A1(n12197), .A2(n3824), .A3(n3795), .ZN(n3863) );
  NAND2_X1 U5118 ( .A1(n5111), .A2(n8050), .ZN(n3797) );
  AND2_X1 U5119 ( .A1(n3758), .A2(pmp_addr_i[30]), .ZN(n8063) );
  AND2_X1 U5120 ( .A1(n3758), .A2(pmp_addr_i[31]), .ZN(n8066) );
  INV_X1 U5121 ( .A(n8033), .ZN(n3802) );
  NOR2_X1 U5122 ( .A1(n5208), .A2(n3802), .ZN(n3803) );
  INV_X1 U5123 ( .A(n8038), .ZN(n3805) );
  NOR2_X1 U5124 ( .A1(n4644), .A2(n3805), .ZN(n3807) );
  AOI22_X1 U5125 ( .A1(n3808), .A2(n3807), .B1(n3806), .B2(n8039), .ZN(n3809)
         );
  NAND2_X1 U5126 ( .A1(n3825), .A2(n3811), .ZN(n3812) );
  OAI22_X1 U5127 ( .A1(n5100), .A2(n3814), .B1(n4802), .B2(n3813), .ZN(n3816)
         );
  NAND4_X1 U5128 ( .A1(n3817), .A2(n3816), .A3(n3818), .A4(n3815), .ZN(n3822)
         );
  NAND3_X1 U5129 ( .A1(n3819), .A2(n3818), .A3(n8025), .ZN(n3821) );
  NAND2_X1 U5130 ( .A1(n999), .A2(n8026), .ZN(n3820) );
  NAND3_X1 U5131 ( .A1(n3822), .A2(n3821), .A3(n3820), .ZN(n3823) );
  NAND3_X1 U5132 ( .A1(n3825), .A2(n3824), .A3(n3823), .ZN(n3826) );
  OAI211_X1 U5133 ( .C1(n3828), .C2(n3863), .A(n3827), .B(n3826), .ZN(n3867)
         );
  AND2_X1 U5134 ( .A1(n3758), .A2(pmp_addr_i[4]), .ZN(n7947) );
  INV_X1 U5135 ( .A(n7947), .ZN(n3829) );
  NAND2_X1 U5136 ( .A1(instr_addr_o_6_), .A2(n3829), .ZN(n3838) );
  AND2_X1 U5137 ( .A1(n3758), .A2(pmp_addr_i[3]), .ZN(n7946) );
  INV_X1 U5138 ( .A(n7946), .ZN(n3830) );
  NOR2_X1 U5139 ( .A1(n5280), .A2(n3830), .ZN(n3831) );
  AOI22_X1 U5140 ( .A1(n3838), .A2(n3831), .B1(n2611), .B2(n7947), .ZN(n3843)
         );
  AND2_X1 U5141 ( .A1(n3758), .A2(pmp_addr_i[1]), .ZN(n7938) );
  AND2_X1 U5142 ( .A1(n3758), .A2(pmp_addr_i[0]), .ZN(n7937) );
  OR2_X1 U5143 ( .A1(n7938), .A2(n7937), .ZN(n3832) );
  AND2_X1 U5144 ( .A1(n3758), .A2(pmp_addr_i[2]), .ZN(n7942) );
  NOR2_X1 U5145 ( .A1(n3832), .A2(n7942), .ZN(n3835) );
  INV_X1 U5146 ( .A(n3832), .ZN(n3834) );
  INV_X1 U5147 ( .A(n7942), .ZN(n3833) );
  OAI22_X1 U5148 ( .A1(n3836), .A2(n3835), .B1(n3834), .B2(n3833), .ZN(n3837)
         );
  OAI211_X1 U5149 ( .C1(n7946), .C2(n3839), .A(n3838), .B(n3837), .ZN(n3842)
         );
  AND2_X1 U5150 ( .A1(n3758), .A2(pmp_addr_i[5]), .ZN(n7957) );
  AND2_X1 U5151 ( .A1(n3758), .A2(pmp_addr_i[6]), .ZN(n7958) );
  INV_X1 U5152 ( .A(n7958), .ZN(n3840) );
  NAND2_X1 U5153 ( .A1(instr_addr_o_8_), .A2(n3840), .ZN(n3845) );
  OAI21_X1 U5154 ( .B1(n3844), .B2(n7957), .A(n3845), .ZN(n3841) );
  AOI21_X1 U5155 ( .B1(n3843), .B2(n3842), .A(n3841), .ZN(n3862) );
  NAND3_X1 U5156 ( .A1(n3845), .A2(n3844), .A3(n7957), .ZN(n3850) );
  AND2_X1 U5157 ( .A1(n3758), .A2(pmp_addr_i[8]), .ZN(n7963) );
  INV_X1 U5158 ( .A(n7963), .ZN(n3851) );
  NOR2_X1 U5159 ( .A1(n213), .A2(n3851), .ZN(n3853) );
  INV_X1 U5160 ( .A(n3853), .ZN(n3849) );
  NAND2_X1 U5161 ( .A1(n4606), .A2(n7958), .ZN(n3848) );
  AND2_X1 U5162 ( .A1(n3758), .A2(pmp_addr_i[7]), .ZN(n7962) );
  NAND2_X1 U5163 ( .A1(n3846), .A2(n7962), .ZN(n3847) );
  NAND4_X1 U5164 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(n3861)
         );
  INV_X1 U5165 ( .A(n7962), .ZN(n3852) );
  AOI22_X1 U5166 ( .A1(instr_addr_o_9_), .A2(n3852), .B1(instr_addr_o_10_), 
        .B2(n3851), .ZN(n3854) );
  NOR2_X1 U5167 ( .A1(n3854), .A2(n3853), .ZN(n3858) );
  OAI21_X1 U5168 ( .B1(n5052), .B2(n7974), .A(n3855), .ZN(n3856) );
  NOR3_X1 U5169 ( .A1(n3858), .A2(n3857), .A3(n3856), .ZN(n3860) );
  OAI211_X1 U5170 ( .C1(n3862), .C2(n3861), .A(n3860), .B(n3859), .ZN(n3864)
         );
  NOR2_X1 U5171 ( .A1(n3864), .A2(n3863), .ZN(n3866) );
  OAI211_X1 U5172 ( .C1(n3867), .C2(n3866), .A(pmp_cfg_i[2]), .B(n3865), .ZN(
        n3868) );
  NOR2_X1 U5173 ( .A1(n12131), .A2(n12229), .ZN(n6049) );
  NAND2_X1 U5174 ( .A1(pmp_addr_i[480]), .A2(pmp_addr_i[481]), .ZN(n3877) );
  NOR2_X1 U5175 ( .A1(n3877), .A2(n4077), .ZN(n4673) );
  NAND2_X1 U5176 ( .A1(n4673), .A2(pmp_addr_i[483]), .ZN(n11785) );
  INV_X1 U5177 ( .A(pmp_cfg_i[123]), .ZN(n3895) );
  OAI21_X1 U5178 ( .B1(n11785), .B2(n3895), .A(pmp_cfg_i[124]), .ZN(n3874) );
  NAND2_X1 U5179 ( .A1(n6624), .A2(pmp_addr_i[452]), .ZN(n3871) );
  OAI21_X1 U5180 ( .B1(n3874), .B2(n4083), .A(n3871), .ZN(n6510) );
  INV_X1 U5181 ( .A(n6510), .ZN(n3888) );
  NOR2_X1 U5182 ( .A1(instr_addr_o_6_), .A2(n3888), .ZN(n3890) );
  INV_X1 U5183 ( .A(pmp_addr_i[483]), .ZN(n3873) );
  NAND2_X1 U5184 ( .A1(n6624), .A2(pmp_addr_i[451]), .ZN(n3872) );
  OAI21_X1 U5185 ( .B1(n3874), .B2(n3873), .A(n3872), .ZN(n6509) );
  INV_X1 U5186 ( .A(n6509), .ZN(n3887) );
  NOR2_X1 U5187 ( .A1(n5280), .A2(n3887), .ZN(n3875) );
  NOR2_X1 U5188 ( .A1(n3890), .A2(n3875), .ZN(n3893) );
  OAI21_X1 U5189 ( .B1(n3877), .B2(n3895), .A(pmp_cfg_i[124]), .ZN(n3881) );
  NAND2_X1 U5190 ( .A1(n6624), .A2(pmp_addr_i[450]), .ZN(n3878) );
  OAI21_X1 U5191 ( .B1(n3881), .B2(n4077), .A(n3878), .ZN(n6506) );
  INV_X1 U5192 ( .A(n6506), .ZN(n6674) );
  NOR2_X1 U5193 ( .A1(n5976), .A2(n6674), .ZN(n3886) );
  INV_X1 U5194 ( .A(pmp_addr_i[481]), .ZN(n3880) );
  NAND2_X1 U5195 ( .A1(n6624), .A2(pmp_addr_i[449]), .ZN(n3879) );
  OAI21_X1 U5196 ( .B1(n3881), .B2(n3880), .A(n3879), .ZN(n6503) );
  INV_X1 U5197 ( .A(n6503), .ZN(n6677) );
  NAND2_X1 U5198 ( .A1(n6624), .A2(pmp_addr_i[448]), .ZN(n3883) );
  NAND2_X1 U5199 ( .A1(n3895), .A2(pmp_addr_i[480]), .ZN(n3882) );
  NAND2_X1 U5200 ( .A1(n6677), .A2(n323), .ZN(n3885) );
  NAND2_X1 U5201 ( .A1(n5899), .A2(n6674), .ZN(n3884) );
  OAI21_X1 U5202 ( .B1(n3886), .B2(n3885), .A(n3884), .ZN(n3892) );
  NAND2_X1 U5203 ( .A1(n4596), .A2(n3887), .ZN(n3889) );
  NAND2_X1 U5204 ( .A1(n5277), .A2(n3888), .ZN(n4697) );
  OAI21_X1 U5205 ( .B1(n3890), .B2(n3889), .A(n4697), .ZN(n3891) );
  AOI21_X1 U5206 ( .B1(n3893), .B2(n3892), .A(n3891), .ZN(n3921) );
  NAND4_X1 U5207 ( .A1(n4673), .A2(pmp_addr_i[485]), .A3(pmp_addr_i[483]), 
        .A4(pmp_addr_i[484]), .ZN(n11779) );
  OAI21_X1 U5208 ( .B1(n11779), .B2(n3895), .A(pmp_cfg_i[124]), .ZN(n3900) );
  INV_X1 U5209 ( .A(pmp_addr_i[486]), .ZN(n3922) );
  NAND2_X1 U5210 ( .A1(n6624), .A2(pmp_addr_i[454]), .ZN(n3896) );
  OAI21_X1 U5211 ( .B1(n3900), .B2(n3922), .A(n3896), .ZN(n6518) );
  INV_X1 U5212 ( .A(n6518), .ZN(n3909) );
  NOR2_X1 U5213 ( .A1(n5269), .A2(n3909), .ZN(n3911) );
  INV_X1 U5214 ( .A(pmp_addr_i[485]), .ZN(n3898) );
  NAND2_X1 U5215 ( .A1(n6624), .A2(pmp_addr_i[453]), .ZN(n3897) );
  OAI21_X1 U5216 ( .B1(n3900), .B2(n3898), .A(n3897), .ZN(n6519) );
  INV_X1 U5217 ( .A(n6519), .ZN(n3908) );
  NOR2_X1 U5218 ( .A1(n5268), .A2(n3908), .ZN(n3899) );
  NOR2_X1 U5219 ( .A1(n3911), .A2(n3899), .ZN(n3907) );
  INV_X1 U5220 ( .A(n6624), .ZN(n4006) );
  AND2_X1 U5221 ( .A1(pmp_addr_i[487]), .A2(pmp_addr_i[486]), .ZN(n3901) );
  INV_X1 U5222 ( .A(pmp_cfg_i[124]), .ZN(n6673) );
  OAI21_X1 U5223 ( .B1(n3901), .B2(n6673), .A(n3900), .ZN(n3904) );
  NAND2_X1 U5224 ( .A1(n3904), .A2(pmp_addr_i[488]), .ZN(n3902) );
  OAI21_X1 U5225 ( .B1(n4006), .B2(n3903), .A(n3902), .ZN(n6525) );
  INV_X1 U5226 ( .A(n6525), .ZN(n3912) );
  NOR2_X1 U5227 ( .A1(n214), .A2(n3912), .ZN(n3915) );
  NAND2_X1 U5228 ( .A1(n3904), .A2(pmp_addr_i[487]), .ZN(n3905) );
  OAI21_X1 U5229 ( .B1(n4006), .B2(n3906), .A(n3905), .ZN(n6672) );
  INV_X1 U5230 ( .A(n6672), .ZN(n6654) );
  NOR2_X1 U5231 ( .A1(n5040), .A2(n6654), .ZN(n4708) );
  NOR2_X1 U5232 ( .A1(n3915), .A2(n4708), .ZN(n3918) );
  NAND2_X1 U5233 ( .A1(n3907), .A2(n3918), .ZN(n3920) );
  NAND2_X1 U5234 ( .A1(n4605), .A2(n3908), .ZN(n4699) );
  NAND2_X1 U5235 ( .A1(n5342), .A2(n3909), .ZN(n3910) );
  OAI21_X1 U5236 ( .B1(n3911), .B2(n4699), .A(n3910), .ZN(n3917) );
  NAND2_X1 U5237 ( .A1(n5040), .A2(n6654), .ZN(n3914) );
  NAND2_X1 U5238 ( .A1(n214), .A2(n3912), .ZN(n3913) );
  OAI21_X1 U5239 ( .B1(n3915), .B2(n3914), .A(n3913), .ZN(n3916) );
  AOI21_X1 U5240 ( .B1(n3918), .B2(n3917), .A(n3916), .ZN(n3919) );
  OAI21_X1 U5241 ( .B1(n3921), .B2(n3920), .A(n3919), .ZN(n3978) );
  OR2_X1 U5242 ( .A1(n11779), .A2(n3922), .ZN(n11769) );
  NAND2_X1 U5243 ( .A1(pmp_addr_i[487]), .A2(pmp_addr_i[488]), .ZN(n3923) );
  NAND2_X1 U5244 ( .A1(n4681), .A2(pmp_cfg_i[123]), .ZN(n3931) );
  NAND2_X1 U5245 ( .A1(pmp_addr_i[489]), .A2(pmp_addr_i[490]), .ZN(n3927) );
  INV_X1 U5246 ( .A(pmp_addr_i[491]), .ZN(n3929) );
  NOR2_X1 U5247 ( .A1(n3927), .A2(n3929), .ZN(n3945) );
  INV_X1 U5248 ( .A(n3945), .ZN(n3924) );
  OR2_X1 U5249 ( .A1(n3931), .A2(n3924), .ZN(n3940) );
  NAND3_X1 U5250 ( .A1(n3940), .A2(pmp_addr_i[492]), .A3(pmp_cfg_i[124]), .ZN(
        n3925) );
  OAI21_X1 U5251 ( .B1(n4006), .B2(n3926), .A(n3925), .ZN(n6653) );
  INV_X1 U5252 ( .A(n6653), .ZN(n4733) );
  NOR2_X1 U5253 ( .A1(n4788), .A2(n4733), .ZN(n3961) );
  OAI21_X1 U5254 ( .B1(n3931), .B2(n3927), .A(pmp_cfg_i[124]), .ZN(n3936) );
  NAND2_X1 U5255 ( .A1(n6624), .A2(pmp_addr_i[459]), .ZN(n3928) );
  OAI21_X1 U5256 ( .B1(n3936), .B2(n3929), .A(n3928), .ZN(n6531) );
  INV_X1 U5257 ( .A(n6531), .ZN(n3959) );
  NOR2_X1 U5258 ( .A1(n5997), .A2(n3959), .ZN(n3930) );
  NOR2_X1 U5259 ( .A1(n3961), .A2(n3930), .ZN(n3964) );
  NAND3_X1 U5260 ( .A1(n3931), .A2(pmp_addr_i[489]), .A3(pmp_cfg_i[124]), .ZN(
        n3932) );
  OAI21_X1 U5261 ( .B1(n4006), .B2(n3933), .A(n3932), .ZN(n6527) );
  INV_X1 U5262 ( .A(n6527), .ZN(n3955) );
  NOR2_X1 U5263 ( .A1(n5069), .A2(n3955), .ZN(n3937) );
  INV_X1 U5264 ( .A(pmp_addr_i[490]), .ZN(n4685) );
  NAND2_X1 U5265 ( .A1(n6624), .A2(pmp_addr_i[458]), .ZN(n3935) );
  OAI21_X1 U5266 ( .B1(n3936), .B2(n4685), .A(n3935), .ZN(n6528) );
  NOR2_X1 U5267 ( .A1(n4494), .A2(n6683), .ZN(n3958) );
  NOR2_X1 U5268 ( .A1(n3937), .A2(n3958), .ZN(n3938) );
  NAND2_X1 U5269 ( .A1(n3964), .A2(n3938), .ZN(n3954) );
  NAND2_X1 U5270 ( .A1(pmp_addr_i[493]), .A2(pmp_addr_i[492]), .ZN(n3939) );
  OAI21_X1 U5271 ( .B1(n3940), .B2(n3939), .A(pmp_cfg_i[124]), .ZN(n3943) );
  INV_X1 U5272 ( .A(pmp_addr_i[493]), .ZN(n3947) );
  NAND2_X1 U5273 ( .A1(n6624), .A2(pmp_addr_i[461]), .ZN(n3941) );
  OAI21_X1 U5274 ( .B1(n3943), .B2(n3947), .A(n3941), .ZN(n6533) );
  NOR2_X1 U5275 ( .A1(n12178), .A2(n4730), .ZN(n3944) );
  INV_X1 U5276 ( .A(pmp_addr_i[494]), .ZN(n3948) );
  NAND2_X1 U5277 ( .A1(n6624), .A2(pmp_addr_i[462]), .ZN(n3942) );
  OAI21_X1 U5278 ( .B1(n3943), .B2(n3948), .A(n3942), .ZN(n6554) );
  INV_X1 U5279 ( .A(n6554), .ZN(n3965) );
  NOR2_X1 U5280 ( .A1(n4743), .A2(n3965), .ZN(n3967) );
  NOR2_X1 U5281 ( .A1(n3944), .A2(n3967), .ZN(n3953) );
  NAND2_X1 U5282 ( .A1(n4681), .A2(n3945), .ZN(n11762) );
  INV_X1 U5283 ( .A(pmp_addr_i[492]), .ZN(n3946) );
  OR2_X1 U5284 ( .A1(n11762), .A2(n3946), .ZN(n4684) );
  OR2_X1 U5285 ( .A1(n4684), .A2(n3947), .ZN(n11807) );
  AND2_X1 U5287 ( .A1(pmp_cfg_i[123]), .A2(pmp_addr_i[495]), .ZN(n3949) );
  AOI21_X2 U5288 ( .B1(n11790), .B2(n3949), .A(n6673), .ZN(n4674) );
  NAND2_X1 U5289 ( .A1(n4674), .A2(pmp_addr_i[495]), .ZN(n3950) );
  OAI21_X1 U5290 ( .B1(n2641), .B2(n4006), .A(n3950), .ZN(n11793) );
  INV_X1 U5291 ( .A(n11793), .ZN(n4719) );
  NAND2_X1 U5292 ( .A1(n4674), .A2(pmp_addr_i[496]), .ZN(n3951) );
  OAI21_X1 U5293 ( .B1(n2636), .B2(n4006), .A(n3951), .ZN(n6648) );
  NOR2_X1 U5294 ( .A1(n3952), .A2(n3969), .ZN(n3972) );
  NAND2_X1 U5295 ( .A1(n3972), .A2(n3953), .ZN(n3974) );
  NOR2_X1 U5296 ( .A1(n3954), .A2(n3974), .ZN(n3977) );
  NAND2_X1 U5297 ( .A1(n6002), .A2(n3955), .ZN(n3957) );
  NAND2_X1 U5298 ( .A1(instr_addr_o_12_), .A2(n6683), .ZN(n3956) );
  OAI21_X1 U5299 ( .B1(n3958), .B2(n3957), .A(n3956), .ZN(n3963) );
  NAND2_X1 U5300 ( .A1(n5997), .A2(n3959), .ZN(n4698) );
  AOI21_X1 U5301 ( .B1(n3964), .B2(n3963), .A(n3962), .ZN(n3975) );
  NAND2_X1 U5302 ( .A1(n4498), .A2(n4730), .ZN(n4694) );
  NAND2_X1 U5303 ( .A1(n5229), .A2(n3965), .ZN(n3966) );
  OAI21_X1 U5304 ( .B1(n3967), .B2(n4694), .A(n3966), .ZN(n3971) );
  NAND2_X1 U5305 ( .A1(n5974), .A2(n4719), .ZN(n4703) );
  OAI21_X1 U5306 ( .B1(n3969), .B2(n4703), .A(n3968), .ZN(n3970) );
  AOI21_X1 U5307 ( .B1(n3972), .B2(n3971), .A(n3970), .ZN(n3973) );
  OAI21_X1 U5308 ( .B1(n3975), .B2(n3974), .A(n3973), .ZN(n3976) );
  AOI21_X1 U5309 ( .B1(n3978), .B2(n3977), .A(n3976), .ZN(n4056) );
  INV_X1 U5310 ( .A(pmp_addr_i[466]), .ZN(n3980) );
  NAND2_X1 U5311 ( .A1(n4674), .A2(pmp_addr_i[498]), .ZN(n3979) );
  OAI21_X1 U5312 ( .B1(n3980), .B2(n4006), .A(n3979), .ZN(n6645) );
  INV_X1 U5313 ( .A(n6645), .ZN(n4013) );
  NOR2_X1 U5314 ( .A1(n5187), .A2(n4013), .ZN(n4016) );
  NAND2_X1 U5315 ( .A1(n4674), .A2(pmp_addr_i[497]), .ZN(n3981) );
  OAI21_X1 U5316 ( .B1(n2665), .B2(n4006), .A(n3981), .ZN(n6644) );
  NOR2_X1 U5317 ( .A1(n4907), .A2(n6558), .ZN(n3982) );
  NOR2_X1 U5318 ( .A1(n4016), .A2(n3982), .ZN(n3987) );
  NAND2_X1 U5319 ( .A1(n4674), .A2(pmp_addr_i[500]), .ZN(n3983) );
  OAI21_X1 U5320 ( .B1(n2571), .B2(n4006), .A(n3983), .ZN(n6627) );
  NOR2_X1 U5321 ( .A1(n5181), .A2(n6569), .ZN(n4019) );
  INV_X1 U5322 ( .A(n3984), .ZN(n4533) );
  NAND2_X1 U5323 ( .A1(n4674), .A2(pmp_addr_i[499]), .ZN(n3985) );
  OAI21_X1 U5324 ( .B1(n2573), .B2(n4006), .A(n3985), .ZN(n6626) );
  NOR2_X1 U5325 ( .A1(n4533), .A2(n6565), .ZN(n3986) );
  NOR2_X1 U5326 ( .A1(n4019), .A2(n3986), .ZN(n4022) );
  NAND2_X1 U5327 ( .A1(n3987), .A2(n4022), .ZN(n3996) );
  NAND2_X1 U5329 ( .A1(n4674), .A2(pmp_addr_i[502]), .ZN(n3988) );
  OAI21_X1 U5330 ( .B1(n2566), .B2(n4006), .A(n3988), .ZN(n6629) );
  NOR2_X1 U5331 ( .A1(instr_addr_o_24_), .A2(n6591), .ZN(n4025) );
  NAND2_X1 U5332 ( .A1(n4674), .A2(pmp_addr_i[501]), .ZN(n3989) );
  OAI21_X1 U5333 ( .B1(n2579), .B2(n4006), .A(n3989), .ZN(n6628) );
  NOR2_X1 U5334 ( .A1(n4859), .A2(n6570), .ZN(n3990) );
  NOR2_X1 U5335 ( .A1(n4025), .A2(n3990), .ZN(n3995) );
  NAND2_X1 U5336 ( .A1(n4674), .A2(pmp_addr_i[504]), .ZN(n3991) );
  OAI21_X1 U5337 ( .B1(n2565), .B2(n4006), .A(n3991), .ZN(n6635) );
  NOR2_X1 U5338 ( .A1(n4909), .A2(n6595), .ZN(n4029) );
  INV_X1 U5339 ( .A(n3992), .ZN(instr_addr_o_25_) );
  NAND2_X1 U5340 ( .A1(n4674), .A2(pmp_addr_i[503]), .ZN(n3993) );
  OAI21_X1 U5341 ( .B1(n2583), .B2(n4006), .A(n3993), .ZN(n6634) );
  INV_X1 U5342 ( .A(n6634), .ZN(n4026) );
  NOR2_X1 U5343 ( .A1(n5365), .A2(n4026), .ZN(n3994) );
  NOR2_X1 U5344 ( .A1(n4029), .A2(n3994), .ZN(n4032) );
  NAND2_X1 U5345 ( .A1(n3995), .A2(n4032), .ZN(n4034) );
  NOR2_X1 U5346 ( .A1(n3996), .A2(n4034), .ZN(n4012) );
  NAND2_X1 U5347 ( .A1(n4674), .A2(pmp_addr_i[508]), .ZN(n3997) );
  OAI21_X1 U5348 ( .B1(n2562), .B2(n4006), .A(n3997), .ZN(n6637) );
  NAND2_X1 U5349 ( .A1(n4674), .A2(pmp_addr_i[507]), .ZN(n3998) );
  OAI21_X1 U5350 ( .B1(n2597), .B2(n4006), .A(n3998), .ZN(n6664) );
  NOR2_X1 U5351 ( .A1(n4900), .A2(n6604), .ZN(n3999) );
  NOR2_X1 U5352 ( .A1(n4041), .A2(n3999), .ZN(n4044) );
  NAND2_X1 U5353 ( .A1(n4674), .A2(pmp_addr_i[505]), .ZN(n4001) );
  OAI21_X1 U5354 ( .B1(n2594), .B2(n4006), .A(n4001), .ZN(n6663) );
  NOR2_X1 U5355 ( .A1(n4556), .A2(n6596), .ZN(n4003) );
  NAND2_X1 U5356 ( .A1(n4674), .A2(pmp_addr_i[506]), .ZN(n4002) );
  OAI21_X1 U5357 ( .B1(n2563), .B2(n4006), .A(n4002), .ZN(n6636) );
  NOR2_X1 U5358 ( .A1(n5368), .A2(n6603), .ZN(n4038) );
  NOR2_X1 U5359 ( .A1(n4003), .A2(n4038), .ZN(n4004) );
  NAND2_X1 U5360 ( .A1(n4044), .A2(n4004), .ZN(n4011) );
  NAND2_X1 U5361 ( .A1(n4674), .A2(pmp_addr_i[509]), .ZN(n12103) );
  OAI21_X1 U5362 ( .B1(n4006), .B2(n2590), .A(n12103), .ZN(n6671) );
  INV_X1 U5363 ( .A(n6671), .ZN(n4045) );
  NOR2_X1 U5364 ( .A1(n147), .A2(n4045), .ZN(n4008) );
  INV_X1 U5365 ( .A(pmp_addr_i[478]), .ZN(n4007) );
  NOR2_X1 U5366 ( .A1(n4008), .A2(pmp_addr_i[478]), .ZN(n4010) );
  INV_X1 U5367 ( .A(pmp_addr_i[479]), .ZN(n4009) );
  NAND2_X1 U5368 ( .A1(n4010), .A2(n4009), .ZN(n4049) );
  NOR2_X1 U5369 ( .A1(n4011), .A2(n4049), .ZN(n4052) );
  NAND2_X1 U5370 ( .A1(n4012), .A2(n4052), .ZN(n4055) );
  NAND2_X1 U5371 ( .A1(n4907), .A2(n6558), .ZN(n4015) );
  NAND2_X1 U5372 ( .A1(n4802), .A2(n4013), .ZN(n4014) );
  OAI21_X1 U5373 ( .B1(n4016), .B2(n4015), .A(n4014), .ZN(n4021) );
  NAND2_X1 U5374 ( .A1(n4533), .A2(n6565), .ZN(n4018) );
  NAND2_X1 U5375 ( .A1(instr_addr_o_22_), .A2(n6569), .ZN(n4017) );
  OAI21_X1 U5376 ( .B1(n4019), .B2(n4018), .A(n4017), .ZN(n4020) );
  AOI21_X1 U5377 ( .B1(n4022), .B2(n4021), .A(n4020), .ZN(n4035) );
  NAND2_X1 U5378 ( .A1(n4859), .A2(n6570), .ZN(n4024) );
  NAND2_X1 U5379 ( .A1(instr_addr_o_24_), .A2(n6591), .ZN(n4023) );
  OAI21_X1 U5380 ( .B1(n4025), .B2(n4024), .A(n4023), .ZN(n4031) );
  NAND2_X1 U5381 ( .A1(instr_addr_o_25_), .A2(n4026), .ZN(n4028) );
  NAND2_X1 U5382 ( .A1(n4909), .A2(n6595), .ZN(n4027) );
  OAI21_X1 U5383 ( .B1(n4029), .B2(n4028), .A(n4027), .ZN(n4030) );
  AOI21_X1 U5384 ( .B1(n4032), .B2(n4031), .A(n4030), .ZN(n4033) );
  OAI21_X1 U5385 ( .B1(n4035), .B2(n4034), .A(n4033), .ZN(n4053) );
  NAND2_X1 U5386 ( .A1(n4556), .A2(n6596), .ZN(n4037) );
  NAND2_X1 U5387 ( .A1(n5979), .A2(n6603), .ZN(n4036) );
  OAI21_X1 U5388 ( .B1(n4038), .B2(n4037), .A(n4036), .ZN(n4043) );
  NAND2_X1 U5389 ( .A1(n4560), .A2(n6608), .ZN(n4039) );
  OAI21_X1 U5390 ( .B1(n4041), .B2(n4040), .A(n4039), .ZN(n4042) );
  AOI21_X1 U5391 ( .B1(n4044), .B2(n4043), .A(n4042), .ZN(n4050) );
  NAND2_X1 U5392 ( .A1(n147), .A2(n4045), .ZN(n4046) );
  NOR2_X1 U5393 ( .A1(n4046), .A2(pmp_addr_i[478]), .ZN(n4047) );
  NAND2_X1 U5394 ( .A1(n4047), .A2(n4009), .ZN(n4048) );
  OAI21_X1 U5395 ( .B1(n4050), .B2(n4049), .A(n4048), .ZN(n4051) );
  AOI21_X1 U5396 ( .B1(n4053), .B2(n4052), .A(n4051), .ZN(n4054) );
  OAI21_X1 U5397 ( .B1(n4056), .B2(n4055), .A(n4054), .ZN(n4166) );
  INV_X1 U5398 ( .A(pmp_addr_i[496]), .ZN(n4057) );
  NAND2_X1 U5399 ( .A1(n5047), .A2(n4057), .ZN(n4071) );
  OAI21_X1 U5400 ( .B1(n5048), .B2(pmp_addr_i[495]), .A(n4071), .ZN(n4073) );
  OAI21_X1 U5402 ( .B1(n6017), .B2(pmp_addr_i[493]), .A(n4068), .ZN(n4058) );
  NOR2_X1 U5403 ( .A1(n4073), .A2(n4058), .ZN(n4103) );
  NAND2_X1 U5404 ( .A1(n4494), .A2(n4685), .ZN(n4094) );
  INV_X1 U5405 ( .A(pmp_addr_i[489]), .ZN(n4059) );
  NOR2_X1 U5406 ( .A1(n4493), .A2(n4059), .ZN(n4060) );
  AOI22_X1 U5407 ( .A1(n4094), .A2(n4060), .B1(n5070), .B2(pmp_addr_i[490]), 
        .ZN(n4066) );
  NAND2_X1 U5408 ( .A1(n4788), .A2(n3946), .ZN(n4064) );
  NAND2_X1 U5409 ( .A1(n4061), .A2(n3929), .ZN(n4062) );
  NAND2_X1 U5410 ( .A1(n4064), .A2(n4062), .ZN(n4096) );
  NOR2_X1 U5411 ( .A1(n937), .A2(n3929), .ZN(n4063) );
  AOI22_X1 U5412 ( .A1(n4064), .A2(n4063), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[492]), .ZN(n4065) );
  OAI21_X1 U5413 ( .B1(n4066), .B2(n4096), .A(n4065), .ZN(n4076) );
  NOR2_X1 U5414 ( .A1(n5057), .A2(n3947), .ZN(n4067) );
  AOI22_X1 U5415 ( .A1(n4068), .A2(n4067), .B1(n5058), .B2(pmp_addr_i[494]), 
        .ZN(n4074) );
  AOI22_X1 U5416 ( .A1(n4071), .A2(n4070), .B1(n2750), .B2(pmp_addr_i[496]), 
        .ZN(n4072) );
  OAI21_X1 U5417 ( .B1(n4074), .B2(n4073), .A(n4072), .ZN(n4075) );
  AOI21_X1 U5418 ( .B1(n4103), .B2(n4076), .A(n4075), .ZN(n4118) );
  INV_X1 U5419 ( .A(pmp_addr_i[484]), .ZN(n4083) );
  NOR2_X1 U5420 ( .A1(n5277), .A2(n4083), .ZN(n4086) );
  NOR2_X1 U5421 ( .A1(pmp_addr_i[481]), .A2(pmp_addr_i[480]), .ZN(n4078) );
  INV_X1 U5422 ( .A(pmp_addr_i[482]), .ZN(n4077) );
  OAI22_X1 U5423 ( .A1(n6015), .A2(n3873), .B1(n4078), .B2(n4077), .ZN(n4082)
         );
  INV_X1 U5424 ( .A(n4078), .ZN(n4079) );
  NOR2_X1 U5425 ( .A1(n4079), .A2(pmp_addr_i[482]), .ZN(n4080) );
  NOR2_X1 U5426 ( .A1(n5291), .A2(n4080), .ZN(n4081) );
  NOR3_X1 U5427 ( .A1(n4086), .A2(n4082), .A3(n4081), .ZN(n4093) );
  NAND2_X1 U5428 ( .A1(n5293), .A2(n3873), .ZN(n4085) );
  AOI22_X1 U5429 ( .A1(instr_addr_o_6_), .A2(n4083), .B1(n12267), .B2(n3898), 
        .ZN(n4084) );
  NAND2_X1 U5430 ( .A1(instr_addr_o_8_), .A2(n3922), .ZN(n4090) );
  OAI211_X1 U5431 ( .C1(n4086), .C2(n4085), .A(n4084), .B(n4090), .ZN(n4092)
         );
  INV_X1 U5432 ( .A(pmp_addr_i[488]), .ZN(n4087) );
  NAND2_X1 U5433 ( .A1(n5262), .A2(n4087), .ZN(n4098) );
  NOR2_X1 U5434 ( .A1(n4605), .A2(n3898), .ZN(n4089) );
  AOI22_X1 U5435 ( .A1(n4090), .A2(n4089), .B1(n4606), .B2(pmp_addr_i[486]), 
        .ZN(n4091) );
  OAI211_X1 U5436 ( .C1(n4093), .C2(n4092), .A(n4100), .B(n4091), .ZN(n4104)
         );
  OAI21_X1 U5437 ( .B1(n5052), .B2(pmp_addr_i[489]), .A(n4094), .ZN(n4095) );
  NOR2_X1 U5438 ( .A1(n4096), .A2(n4095), .ZN(n4102) );
  NAND2_X1 U5439 ( .A1(instr_addr_o_9_), .A2(n11761), .ZN(n4097) );
  NAND2_X1 U5440 ( .A1(n4098), .A2(n4097), .ZN(n4099) );
  NAND2_X1 U5441 ( .A1(n4100), .A2(n4099), .ZN(n4101) );
  NAND4_X1 U5442 ( .A1(n4104), .A2(n4103), .A3(n4102), .A4(n4101), .ZN(n4117)
         );
  INV_X1 U5443 ( .A(pmp_addr_i[506]), .ZN(n4105) );
  NAND2_X1 U5444 ( .A1(n5979), .A2(n4105), .ZN(n4148) );
  OAI21_X1 U5445 ( .B1(n5094), .B2(pmp_addr_i[505]), .A(n4148), .ZN(n4120) );
  INV_X1 U5446 ( .A(pmp_addr_i[504]), .ZN(n4106) );
  NAND2_X1 U5447 ( .A1(n12158), .A2(n4106), .ZN(n4140) );
  INV_X1 U5448 ( .A(pmp_addr_i[503]), .ZN(n4138) );
  NAND2_X1 U5449 ( .A1(n137), .A2(n4138), .ZN(n4107) );
  NAND2_X1 U5450 ( .A1(n4140), .A2(n4107), .ZN(n4142) );
  NOR2_X1 U5451 ( .A1(n4120), .A2(n4142), .ZN(n4115) );
  OAI21_X1 U5452 ( .B1(n4406), .B2(pmp_addr_i[507]), .A(n4151), .ZN(n4146) );
  INV_X1 U5453 ( .A(pmp_addr_i[498]), .ZN(n4108) );
  NAND2_X1 U5454 ( .A1(n5187), .A2(n4108), .ZN(n4122) );
  OAI211_X1 U5455 ( .C1(n5313), .C2(pmp_addr_i[497]), .A(n4152), .B(n4122), 
        .ZN(n4109) );
  NOR2_X1 U5456 ( .A1(n4146), .A2(n4109), .ZN(n4114) );
  INV_X1 U5457 ( .A(pmp_addr_i[500]), .ZN(n4110) );
  NAND2_X1 U5458 ( .A1(n5181), .A2(n4110), .ZN(n4126) );
  INV_X1 U5459 ( .A(pmp_addr_i[499]), .ZN(n4125) );
  NAND2_X1 U5460 ( .A1(n5191), .A2(n4125), .ZN(n4111) );
  INV_X1 U5461 ( .A(pmp_addr_i[502]), .ZN(n4112) );
  NAND2_X1 U5462 ( .A1(n6028), .A2(n4112), .ZN(n4137) );
  INV_X1 U5463 ( .A(pmp_addr_i[501]), .ZN(n4134) );
  NAND2_X1 U5464 ( .A1(n5208), .A2(n4134), .ZN(n4113) );
  AND2_X1 U5465 ( .A1(n4137), .A2(n4113), .ZN(n4132) );
  NAND4_X1 U5466 ( .A1(n4115), .A2(n4114), .A3(n4124), .A4(n4132), .ZN(n4116)
         );
  AOI21_X1 U5467 ( .B1(n4118), .B2(n4117), .A(n4116), .ZN(n4163) );
  INV_X1 U5468 ( .A(n4152), .ZN(n4119) );
  INV_X1 U5469 ( .A(n4142), .ZN(n4133) );
  INV_X1 U5470 ( .A(pmp_addr_i[497]), .ZN(n4121) );
  NOR2_X1 U5471 ( .A1(n5100), .A2(n4121), .ZN(n4123) );
  AOI22_X1 U5472 ( .A1(n4123), .A2(n4122), .B1(n2569), .B2(pmp_addr_i[498]), 
        .ZN(n4130) );
  NOR2_X1 U5473 ( .A1(n5842), .A2(n4125), .ZN(n4127) );
  AOI22_X1 U5474 ( .A1(n4127), .A2(n4126), .B1(n5192), .B2(pmp_addr_i[500]), 
        .ZN(n4128) );
  OAI21_X1 U5475 ( .B1(n4130), .B2(n4129), .A(n4128), .ZN(n4131) );
  NAND4_X1 U5476 ( .A1(n4145), .A2(n4133), .A3(n4132), .A4(n4131), .ZN(n4161)
         );
  NOR2_X1 U5477 ( .A1(n4859), .A2(n4134), .ZN(n4136) );
  AOI22_X1 U5478 ( .A1(n4137), .A2(n4136), .B1(n1269), .B2(pmp_addr_i[502]), 
        .ZN(n4143) );
  NOR2_X1 U5479 ( .A1(n4644), .A2(n4138), .ZN(n4139) );
  AOI22_X1 U5480 ( .A1(n4140), .A2(n4139), .B1(n3806), .B2(pmp_addr_i[504]), 
        .ZN(n4141) );
  OAI21_X1 U5481 ( .B1(n4143), .B2(n4142), .A(n4141), .ZN(n4144) );
  NAND2_X1 U5482 ( .A1(n4145), .A2(n4144), .ZN(n4160) );
  NOR2_X1 U5483 ( .A1(n4146), .A2(n4119), .ZN(n4158) );
  NAND3_X1 U5484 ( .A1(n4148), .A2(pmp_addr_i[505]), .A3(n4147), .ZN(n4150) );
  NAND2_X1 U5485 ( .A1(n4438), .A2(pmp_addr_i[506]), .ZN(n4149) );
  NAND2_X1 U5486 ( .A1(n4150), .A2(n4149), .ZN(n4157) );
  NAND4_X1 U5487 ( .A1(n4151), .A2(n4152), .A3(pmp_addr_i[507]), .A4(n4656), 
        .ZN(n4155) );
  NOR2_X1 U5488 ( .A1(pmp_addr_i[510]), .A2(pmp_addr_i[511]), .ZN(n6484) );
  NAND3_X1 U5489 ( .A1(n4152), .A2(pmp_addr_i[508]), .A3(n4658), .ZN(n4154) );
  NAND2_X1 U5490 ( .A1(n4660), .A2(pmp_addr_i[509]), .ZN(n4153) );
  AOI21_X1 U5491 ( .B1(n4158), .B2(n4157), .A(n4156), .ZN(n4159) );
  OR2_X1 U5492 ( .A1(n4163), .A2(n4162), .ZN(n4165) );
  AND2_X1 U5493 ( .A1(n6624), .A2(pmp_cfg_i[122]), .ZN(n4164) );
  INV_X1 U5494 ( .A(pmp_cfg_i[27]), .ZN(n4194) );
  INV_X1 U5495 ( .A(n7551), .ZN(n4274) );
  INV_X1 U5496 ( .A(pmp_addr_i[68]), .ZN(n5676) );
  NAND2_X1 U5497 ( .A1(pmp_addr_i[96]), .A2(pmp_addr_i[97]), .ZN(n4787) );
  INV_X1 U5498 ( .A(pmp_addr_i[98]), .ZN(n4172) );
  OR2_X1 U5499 ( .A1(n4787), .A2(n4172), .ZN(n4759) );
  NAND2_X1 U5500 ( .A1(pmp_addr_i[100]), .A2(pmp_addr_i[99]), .ZN(n4167) );
  NOR2_X1 U5501 ( .A1(n4759), .A2(n4167), .ZN(n4187) );
  INV_X1 U5502 ( .A(pmp_cfg_i[28]), .ZN(n4229) );
  AOI21_X1 U5503 ( .B1(n4187), .B2(pmp_cfg_i[27]), .A(n4229), .ZN(n4189) );
  NAND2_X1 U5504 ( .A1(n4189), .A2(pmp_addr_i[100]), .ZN(n4168) );
  OAI21_X1 U5505 ( .B1(n4274), .B2(n5676), .A(n4168), .ZN(n7333) );
  INV_X1 U5506 ( .A(n7333), .ZN(n7563) );
  OAI21_X1 U5507 ( .B1(n4759), .B2(n4194), .A(pmp_cfg_i[28]), .ZN(n4173) );
  NAND2_X1 U5508 ( .A1(n7551), .A2(pmp_addr_i[67]), .ZN(n4169) );
  OAI21_X1 U5509 ( .B1(n4173), .B2(n4762), .A(n4169), .ZN(n7332) );
  INV_X1 U5510 ( .A(n7332), .ZN(n4182) );
  NOR2_X1 U5511 ( .A1(n20), .A2(n4182), .ZN(n4170) );
  NOR2_X1 U5512 ( .A1(n4183), .A2(n4170), .ZN(n4186) );
  NAND2_X1 U5513 ( .A1(n7551), .A2(pmp_addr_i[66]), .ZN(n4171) );
  OAI21_X1 U5514 ( .B1(n4173), .B2(n4172), .A(n4171), .ZN(n7560) );
  INV_X1 U5515 ( .A(n7560), .ZN(n4816) );
  NOR2_X1 U5516 ( .A1(n5899), .A2(n4816), .ZN(n4181) );
  AND2_X1 U5517 ( .A1(pmp_cfg_i[27]), .A2(pmp_addr_i[96]), .ZN(n4176) );
  NAND2_X1 U5518 ( .A1(pmp_cfg_i[28]), .A2(pmp_addr_i[97]), .ZN(n4175) );
  NAND2_X1 U5519 ( .A1(n7551), .A2(pmp_addr_i[65]), .ZN(n4174) );
  OAI21_X1 U5520 ( .B1(n4176), .B2(n4175), .A(n4174), .ZN(n7335) );
  INV_X1 U5521 ( .A(n7335), .ZN(n7606) );
  NOR2_X1 U5522 ( .A1(n4229), .A2(pmp_cfg_i[27]), .ZN(n7604) );
  NAND2_X1 U5523 ( .A1(n7604), .A2(pmp_addr_i[96]), .ZN(n4179) );
  NAND2_X1 U5524 ( .A1(n7551), .A2(pmp_addr_i[64]), .ZN(n4178) );
  NAND2_X1 U5525 ( .A1(n7606), .A2(n157), .ZN(n4180) );
  NAND2_X1 U5526 ( .A1(n12150), .A2(n4816), .ZN(n4791) );
  OAI21_X1 U5527 ( .B1(n4181), .B2(n4180), .A(n4791), .ZN(n4185) );
  NAND2_X1 U5528 ( .A1(n20), .A2(n4182), .ZN(n4794) );
  NAND2_X1 U5529 ( .A1(n5277), .A2(n7563), .ZN(n4740) );
  OAI21_X1 U5530 ( .B1(n4183), .B2(n4794), .A(n4740), .ZN(n4184) );
  AOI21_X1 U5531 ( .B1(n4186), .B2(n4185), .A(n4184), .ZN(n4212) );
  NAND3_X1 U5532 ( .A1(n4187), .A2(pmp_addr_i[101]), .A3(pmp_addr_i[102]), 
        .ZN(n4193) );
  OAI21_X1 U5533 ( .B1(n4193), .B2(n4194), .A(pmp_cfg_i[28]), .ZN(n4198) );
  NAND2_X1 U5534 ( .A1(n7551), .A2(pmp_addr_i[70]), .ZN(n4188) );
  OAI21_X1 U5535 ( .B1(n4198), .B2(n4780), .A(n4188), .ZN(n7348) );
  INV_X1 U5536 ( .A(n7348), .ZN(n4201) );
  NOR2_X1 U5537 ( .A1(n205), .A2(n4201), .ZN(n4202) );
  INV_X1 U5538 ( .A(pmp_addr_i[69]), .ZN(n5679) );
  NAND2_X1 U5539 ( .A1(n4189), .A2(pmp_addr_i[101]), .ZN(n4190) );
  OAI21_X1 U5540 ( .B1(n4274), .B2(n5679), .A(n4190), .ZN(n7349) );
  INV_X1 U5541 ( .A(n7349), .ZN(n7557) );
  NOR2_X1 U5542 ( .A1(n5268), .A2(n7557), .ZN(n4191) );
  NOR2_X1 U5543 ( .A1(n4202), .A2(n4191), .ZN(n4199) );
  NAND2_X1 U5544 ( .A1(pmp_addr_i[104]), .A2(pmp_addr_i[103]), .ZN(n4192) );
  OR2_X1 U5545 ( .A1(n4193), .A2(n4192), .ZN(n11730) );
  NOR2_X1 U5546 ( .A1(n11730), .A2(n4194), .ZN(n4217) );
  OR2_X1 U5547 ( .A1(n4217), .A2(n4229), .ZN(n4222) );
  INV_X1 U5548 ( .A(pmp_addr_i[104]), .ZN(n4196) );
  NAND2_X1 U5549 ( .A1(n7551), .A2(pmp_addr_i[72]), .ZN(n4195) );
  OAI21_X1 U5550 ( .B1(n4222), .B2(n4196), .A(n4195), .ZN(n7346) );
  INV_X1 U5551 ( .A(n7346), .ZN(n4205) );
  NOR2_X1 U5552 ( .A1(n213), .A2(n4205), .ZN(n4206) );
  NAND2_X1 U5553 ( .A1(n7551), .A2(pmp_addr_i[71]), .ZN(n4197) );
  OAI21_X1 U5554 ( .B1(n4198), .B2(n4782), .A(n4197), .ZN(n7345) );
  INV_X1 U5555 ( .A(n7345), .ZN(n4203) );
  NOR2_X1 U5556 ( .A1(n4204), .A2(n4203), .ZN(n4824) );
  NOR2_X1 U5557 ( .A1(n4206), .A2(n4824), .ZN(n4209) );
  NAND2_X1 U5558 ( .A1(n4199), .A2(n4209), .ZN(n4211) );
  OR2_X1 U5559 ( .A1(n4200), .A2(n7349), .ZN(n4766) );
  NAND2_X1 U5560 ( .A1(instr_addr_o_8_), .A2(n4201), .ZN(n4779) );
  OAI21_X1 U5561 ( .B1(n4202), .B2(n4766), .A(n4779), .ZN(n4208) );
  NAND2_X1 U5562 ( .A1(n4204), .A2(n4203), .ZN(n4749) );
  OAI21_X1 U5563 ( .B1(n4206), .B2(n4749), .A(n4785), .ZN(n4207) );
  AOI21_X1 U5564 ( .B1(n4209), .B2(n4208), .A(n4207), .ZN(n4210) );
  OAI21_X1 U5565 ( .B1(n4212), .B2(n4211), .A(n4210), .ZN(n4264) );
  NAND2_X1 U5566 ( .A1(pmp_addr_i[105]), .A2(pmp_addr_i[106]), .ZN(n4215) );
  NAND2_X1 U5567 ( .A1(pmp_addr_i[108]), .A2(pmp_addr_i[107]), .ZN(n4213) );
  NOR2_X1 U5568 ( .A1(n4215), .A2(n4213), .ZN(n4235) );
  AOI21_X1 U5569 ( .B1(n4217), .B2(n4235), .A(n4229), .ZN(n4231) );
  NAND2_X1 U5570 ( .A1(n4231), .A2(pmp_addr_i[108]), .ZN(n4214) );
  OAI21_X1 U5571 ( .B1(n4274), .B2(n2056), .A(n4214), .ZN(n7362) );
  INV_X1 U5572 ( .A(n7362), .ZN(n4807) );
  INV_X1 U5573 ( .A(n4215), .ZN(n4216) );
  AOI21_X1 U5574 ( .B1(n4217), .B2(n4216), .A(n4229), .ZN(n4223) );
  NAND2_X1 U5575 ( .A1(n4223), .A2(pmp_addr_i[107]), .ZN(n4218) );
  OAI21_X1 U5576 ( .B1(n4274), .B2(n4219), .A(n4218), .ZN(n7328) );
  NOR2_X1 U5577 ( .A1(n4061), .A2(n7564), .ZN(n4220) );
  NOR2_X1 U5578 ( .A1(n4245), .A2(n4220), .ZN(n4248) );
  NAND2_X1 U5579 ( .A1(n7551), .A2(pmp_addr_i[73]), .ZN(n4221) );
  OAI21_X1 U5580 ( .B1(n4222), .B2(n4771), .A(n4221), .ZN(n7325) );
  NOR2_X1 U5581 ( .A1(n5069), .A2(n7360), .ZN(n4226) );
  NAND2_X1 U5582 ( .A1(n4223), .A2(pmp_addr_i[106]), .ZN(n4224) );
  OAI21_X1 U5583 ( .B1(n4274), .B2(n4225), .A(n4224), .ZN(n7326) );
  INV_X1 U5584 ( .A(n7326), .ZN(n4242) );
  NOR2_X1 U5585 ( .A1(n4494), .A2(n4242), .ZN(n4243) );
  NOR2_X1 U5586 ( .A1(n4226), .A2(n4243), .ZN(n4227) );
  NAND2_X1 U5587 ( .A1(n4248), .A2(n4227), .ZN(n4241) );
  NAND2_X1 U5588 ( .A1(n4231), .A2(pmp_addr_i[109]), .ZN(n4228) );
  OAI21_X1 U5589 ( .B1(n4274), .B2(n2077), .A(n4228), .ZN(n7367) );
  INV_X1 U5590 ( .A(n7367), .ZN(n4810) );
  NOR2_X1 U5591 ( .A1(instr_addr_o_15_), .A2(n4810), .ZN(n4233) );
  NOR2_X1 U5592 ( .A1(n4229), .A2(pmp_addr_i[109]), .ZN(n4230) );
  OAI21_X1 U5593 ( .B1(n4231), .B2(n4230), .A(pmp_addr_i[110]), .ZN(n4232) );
  OAI21_X1 U5594 ( .B1(n4274), .B2(n2055), .A(n4232), .ZN(n7320) );
  NOR2_X1 U5595 ( .A1(n4233), .A2(n4250), .ZN(n4240) );
  INV_X1 U5596 ( .A(n4235), .ZN(n4236) );
  NOR2_X1 U5597 ( .A1(n11730), .A2(n4236), .ZN(n11701) );
  AND3_X1 U5598 ( .A1(pmp_addr_i[109]), .A2(pmp_addr_i[110]), .A3(
        pmp_addr_i[111]), .ZN(n4237) );
  NAND2_X1 U5599 ( .A1(pmp_cfg_i[27]), .A2(pmp_cfg_i[28]), .ZN(n4792) );
  AOI21_X1 U5600 ( .B1(n11701), .B2(n4237), .A(n4792), .ZN(n4761) );
  OR2_X1 U5601 ( .A1(n4761), .A2(n7604), .ZN(n4741) );
  NAND2_X1 U5602 ( .A1(n4741), .A2(pmp_addr_i[111]), .ZN(n4238) );
  OAI21_X1 U5603 ( .B1(n4274), .B2(n2081), .A(n4238), .ZN(n7322) );
  NAND2_X1 U5604 ( .A1(n4741), .A2(pmp_addr_i[112]), .ZN(n4239) );
  OAI21_X1 U5605 ( .B1(n4274), .B2(n2053), .A(n4239), .ZN(n7571) );
  INV_X1 U5606 ( .A(n7571), .ZN(n4252) );
  NOR2_X1 U5607 ( .A1(n337), .A2(n4255), .ZN(n4258) );
  NAND2_X1 U5608 ( .A1(n4240), .A2(n4258), .ZN(n4260) );
  NOR2_X1 U5609 ( .A1(n4241), .A2(n4260), .ZN(n4263) );
  NAND2_X1 U5610 ( .A1(n4494), .A2(n4242), .ZN(n4778) );
  OAI21_X1 U5611 ( .B1(n4243), .B2(n4765), .A(n4778), .ZN(n4247) );
  NAND2_X1 U5612 ( .A1(n5997), .A2(n7564), .ZN(n4748) );
  NAND2_X1 U5613 ( .A1(n206), .A2(n4807), .ZN(n4244) );
  OAI21_X1 U5614 ( .B1(n4245), .B2(n4748), .A(n4244), .ZN(n4246) );
  AOI21_X1 U5615 ( .B1(n4247), .B2(n4248), .A(n4246), .ZN(n4261) );
  NAND2_X1 U5616 ( .A1(n4498), .A2(n4810), .ZN(n4744) );
  NAND2_X1 U5617 ( .A1(n12266), .A2(n7556), .ZN(n4249) );
  OAI21_X1 U5618 ( .B1(n4250), .B2(n4744), .A(n4249), .ZN(n4257) );
  INV_X1 U5619 ( .A(n7322), .ZN(n4251) );
  OAI21_X1 U5620 ( .B1(n4255), .B2(n4254), .A(n4253), .ZN(n4256) );
  AOI21_X1 U5621 ( .B1(n4258), .B2(n4257), .A(n4256), .ZN(n4259) );
  OAI21_X1 U5622 ( .B1(n4261), .B2(n4260), .A(n4259), .ZN(n4262) );
  AOI21_X1 U5623 ( .B1(n4264), .B2(n4263), .A(n4262), .ZN(n4361) );
  NAND2_X1 U5624 ( .A1(n4741), .A2(pmp_addr_i[114]), .ZN(n4265) );
  OAI21_X1 U5625 ( .B1(n4274), .B2(n4266), .A(n4265), .ZN(n7583) );
  INV_X1 U5626 ( .A(n7583), .ZN(n4328) );
  NAND2_X1 U5627 ( .A1(n4741), .A2(pmp_addr_i[113]), .ZN(n4267) );
  OAI21_X1 U5628 ( .B1(n4274), .B2(n4268), .A(n4267), .ZN(n7572) );
  INV_X1 U5629 ( .A(n7572), .ZN(n4327) );
  NOR2_X1 U5630 ( .A1(n4907), .A2(n4327), .ZN(n4269) );
  NOR2_X1 U5631 ( .A1(n4331), .A2(n4269), .ZN(n4276) );
  NAND2_X1 U5632 ( .A1(n4741), .A2(pmp_addr_i[116]), .ZN(n4270) );
  OAI21_X1 U5633 ( .B1(n4274), .B2(n4271), .A(n4270), .ZN(n7585) );
  INV_X1 U5634 ( .A(n7585), .ZN(n4333) );
  NOR2_X1 U5635 ( .A1(n5181), .A2(n4333), .ZN(n4336) );
  NAND2_X1 U5636 ( .A1(n4741), .A2(pmp_addr_i[115]), .ZN(n4272) );
  OAI21_X1 U5637 ( .B1(n4274), .B2(n4273), .A(n4272), .ZN(n7584) );
  INV_X1 U5638 ( .A(n7584), .ZN(n4332) );
  NOR2_X1 U5639 ( .A1(n4533), .A2(n4332), .ZN(n4275) );
  NOR2_X1 U5640 ( .A1(n4336), .A2(n4275), .ZN(n4339) );
  NAND2_X1 U5641 ( .A1(n4276), .A2(n4339), .ZN(n4288) );
  NAND2_X1 U5642 ( .A1(n4741), .A2(pmp_addr_i[118]), .ZN(n4277) );
  OAI21_X1 U5643 ( .B1(n4274), .B2(n4278), .A(n4277), .ZN(n7591) );
  INV_X1 U5644 ( .A(n7591), .ZN(n4341) );
  NOR2_X1 U5645 ( .A1(instr_addr_o_24_), .A2(n4341), .ZN(n4344) );
  NAND2_X1 U5646 ( .A1(n4741), .A2(pmp_addr_i[117]), .ZN(n4279) );
  OAI21_X1 U5647 ( .B1(n4274), .B2(n4280), .A(n4279), .ZN(n7586) );
  INV_X1 U5648 ( .A(n7586), .ZN(n4340) );
  NOR2_X1 U5649 ( .A1(n4859), .A2(n4340), .ZN(n4281) );
  NOR2_X1 U5650 ( .A1(n4344), .A2(n4281), .ZN(n4287) );
  NAND2_X1 U5651 ( .A1(n4741), .A2(pmp_addr_i[120]), .ZN(n4282) );
  OAI21_X1 U5652 ( .B1(n4274), .B2(n4283), .A(n4282), .ZN(n7593) );
  INV_X1 U5653 ( .A(n7593), .ZN(n4346) );
  NOR2_X1 U5654 ( .A1(n4909), .A2(n4346), .ZN(n4349) );
  NAND2_X1 U5655 ( .A1(n4741), .A2(pmp_addr_i[119]), .ZN(n4284) );
  OAI21_X1 U5656 ( .B1(n4274), .B2(n4285), .A(n4284), .ZN(n7592) );
  INV_X1 U5657 ( .A(n7592), .ZN(n4345) );
  NOR2_X1 U5658 ( .A1(instr_addr_o_25_), .A2(n4345), .ZN(n4286) );
  NOR2_X1 U5659 ( .A1(n4349), .A2(n4286), .ZN(n4352) );
  NAND2_X1 U5660 ( .A1(n4287), .A2(n4352), .ZN(n4354) );
  NOR2_X1 U5661 ( .A1(n4288), .A2(n4354), .ZN(n4306) );
  NAND2_X1 U5662 ( .A1(n4741), .A2(pmp_addr_i[124]), .ZN(n4289) );
  OAI21_X1 U5663 ( .B1(n4274), .B2(n4290), .A(n4289), .ZN(n7578) );
  INV_X1 U5664 ( .A(n7578), .ZN(n4313) );
  NOR2_X1 U5665 ( .A1(n4560), .A2(n4313), .ZN(n4316) );
  NAND2_X1 U5666 ( .A1(n4741), .A2(pmp_addr_i[123]), .ZN(n4291) );
  OAI21_X1 U5667 ( .B1(n4274), .B2(n4292), .A(n4291), .ZN(n7603) );
  INV_X1 U5668 ( .A(n7603), .ZN(n4312) );
  NOR2_X1 U5669 ( .A1(n4900), .A2(n4312), .ZN(n4293) );
  NOR2_X1 U5670 ( .A1(n4316), .A2(n4293), .ZN(n4319) );
  NAND2_X1 U5671 ( .A1(n4741), .A2(pmp_addr_i[121]), .ZN(n4294) );
  OAI21_X1 U5672 ( .B1(n4274), .B2(n4295), .A(n4294), .ZN(n7594) );
  INV_X1 U5673 ( .A(n7594), .ZN(n4307) );
  NOR2_X1 U5674 ( .A1(n4556), .A2(n4307), .ZN(n4298) );
  NAND2_X1 U5675 ( .A1(n4741), .A2(pmp_addr_i[122]), .ZN(n4296) );
  OAI21_X1 U5676 ( .B1(n4274), .B2(n4297), .A(n4296), .ZN(n7577) );
  INV_X1 U5677 ( .A(n7577), .ZN(n4308) );
  NOR2_X1 U5678 ( .A1(n5368), .A2(n4308), .ZN(n4311) );
  NOR2_X1 U5679 ( .A1(n4298), .A2(n4311), .ZN(n4299) );
  NAND2_X1 U5680 ( .A1(n4319), .A2(n4299), .ZN(n4305) );
  NAND2_X1 U5681 ( .A1(n4741), .A2(pmp_addr_i[125]), .ZN(n11758) );
  OAI21_X1 U5682 ( .B1(n4274), .B2(n12071), .A(n11758), .ZN(n7614) );
  INV_X1 U5683 ( .A(n7614), .ZN(n4320) );
  NOR2_X1 U5684 ( .A1(n4866), .A2(n4320), .ZN(n4302) );
  INV_X1 U5685 ( .A(pmp_addr_i[94]), .ZN(n4301) );
  NOR2_X1 U5686 ( .A1(n4302), .A2(pmp_addr_i[94]), .ZN(n4304) );
  INV_X1 U5687 ( .A(pmp_addr_i[95]), .ZN(n4303) );
  NAND2_X1 U5688 ( .A1(n4304), .A2(n4303), .ZN(n4324) );
  NOR2_X1 U5689 ( .A1(n4305), .A2(n4324), .ZN(n4356) );
  NAND2_X1 U5690 ( .A1(n4306), .A2(n4356), .ZN(n4360) );
  NAND2_X1 U5691 ( .A1(n4556), .A2(n4307), .ZN(n4310) );
  NAND2_X1 U5692 ( .A1(instr_addr_o_28_), .A2(n4308), .ZN(n4309) );
  OAI21_X1 U5693 ( .B1(n4311), .B2(n4310), .A(n4309), .ZN(n4318) );
  NAND2_X1 U5694 ( .A1(n4900), .A2(n4312), .ZN(n4315) );
  NAND2_X1 U5695 ( .A1(n4560), .A2(n4313), .ZN(n4314) );
  OAI21_X1 U5696 ( .B1(n4316), .B2(n4315), .A(n4314), .ZN(n4317) );
  AOI21_X1 U5697 ( .B1(n4319), .B2(n4318), .A(n4317), .ZN(n4325) );
  NAND2_X1 U5698 ( .A1(instr_addr_o_31_), .A2(n4320), .ZN(n4321) );
  NOR2_X1 U5699 ( .A1(n4321), .A2(pmp_addr_i[94]), .ZN(n4322) );
  NAND2_X1 U5700 ( .A1(n4322), .A2(n4303), .ZN(n4323) );
  OAI21_X1 U5701 ( .B1(n4325), .B2(n4324), .A(n4323), .ZN(n4326) );
  NAND2_X1 U5702 ( .A1(n3793), .A2(n4327), .ZN(n4330) );
  NAND2_X1 U5703 ( .A1(n4802), .A2(n4328), .ZN(n4329) );
  OAI21_X1 U5704 ( .B1(n4331), .B2(n4330), .A(n4329), .ZN(n4338) );
  NAND2_X1 U5705 ( .A1(n4533), .A2(n4332), .ZN(n4335) );
  NAND2_X1 U5706 ( .A1(instr_addr_o_22_), .A2(n4333), .ZN(n4334) );
  OAI21_X1 U5707 ( .B1(n4336), .B2(n4335), .A(n4334), .ZN(n4337) );
  AOI21_X1 U5708 ( .B1(n4339), .B2(n4338), .A(n4337), .ZN(n4355) );
  NAND2_X1 U5709 ( .A1(n4859), .A2(n4340), .ZN(n4343) );
  NAND2_X1 U5710 ( .A1(instr_addr_o_24_), .A2(n4341), .ZN(n4342) );
  OAI21_X1 U5711 ( .B1(n4344), .B2(n4343), .A(n4342), .ZN(n4351) );
  NAND2_X1 U5712 ( .A1(n136), .A2(n4345), .ZN(n4348) );
  NAND2_X1 U5713 ( .A1(n4909), .A2(n4346), .ZN(n4347) );
  OAI21_X1 U5714 ( .B1(n4349), .B2(n4348), .A(n4347), .ZN(n4350) );
  AOI21_X1 U5715 ( .B1(n4352), .B2(n4351), .A(n4350), .ZN(n4353) );
  OAI21_X1 U5716 ( .B1(n4355), .B2(n4354), .A(n4353), .ZN(n4357) );
  NAND2_X1 U5717 ( .A1(n4357), .A2(n4356), .ZN(n4358) );
  OAI211_X1 U5718 ( .C1(n4361), .C2(n4360), .A(n4359), .B(n4358), .ZN(n4453)
         );
  NAND2_X1 U5719 ( .A1(n5047), .A2(n1193), .ZN(n4374) );
  OAI21_X1 U5720 ( .B1(n5048), .B2(pmp_addr_i[111]), .A(n4374), .ZN(n4376) );
  NAND2_X1 U5721 ( .A1(n4743), .A2(n4767), .ZN(n4372) );
  OAI21_X1 U5722 ( .B1(n6017), .B2(pmp_addr_i[109]), .A(n4372), .ZN(n4362) );
  NOR2_X1 U5723 ( .A1(n4376), .A2(n4362), .ZN(n4403) );
  INV_X1 U5724 ( .A(pmp_addr_i[106]), .ZN(n4363) );
  NAND2_X1 U5725 ( .A1(n5250), .A2(n4363), .ZN(n4394) );
  NOR2_X1 U5726 ( .A1(n4493), .A2(n4771), .ZN(n4364) );
  AOI22_X1 U5727 ( .A1(n4394), .A2(n4364), .B1(n5070), .B2(pmp_addr_i[106]), 
        .ZN(n4370) );
  NAND2_X1 U5728 ( .A1(n4788), .A2(n1208), .ZN(n4368) );
  INV_X1 U5729 ( .A(pmp_addr_i[107]), .ZN(n4366) );
  NAND2_X1 U5730 ( .A1(instr_addr_o_13_), .A2(n4366), .ZN(n4365) );
  NAND2_X1 U5731 ( .A1(n4368), .A2(n4365), .ZN(n4396) );
  NOR2_X1 U5732 ( .A1(n5997), .A2(n4366), .ZN(n4367) );
  AOI22_X1 U5733 ( .A1(n4368), .A2(n4367), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[108]), .ZN(n4369) );
  OAI21_X1 U5734 ( .B1(n4370), .B2(n4396), .A(n4369), .ZN(n4379) );
  NOR2_X1 U5735 ( .A1(n5057), .A2(n1200), .ZN(n4371) );
  AOI22_X1 U5736 ( .A1(n4372), .A2(n4371), .B1(n5058), .B2(pmp_addr_i[110]), 
        .ZN(n4377) );
  NOR2_X1 U5737 ( .A1(n5974), .A2(n1196), .ZN(n4373) );
  AOI22_X1 U5738 ( .A1(n4374), .A2(n4373), .B1(instr_addr_o_18__BAR), .B2(
        pmp_addr_i[112]), .ZN(n4375) );
  OAI21_X1 U5739 ( .B1(n4377), .B2(n4376), .A(n4375), .ZN(n4378) );
  AOI21_X1 U5740 ( .B1(n4403), .B2(n4379), .A(n4378), .ZN(n4416) );
  NOR2_X1 U5741 ( .A1(n12152), .A2(n4763), .ZN(n4387) );
  NOR2_X1 U5742 ( .A1(pmp_addr_i[97]), .A2(pmp_addr_i[96]), .ZN(n4380) );
  OAI22_X1 U5743 ( .A1(instr_addr_o_5_), .A2(n4762), .B1(n4380), .B2(n4172), 
        .ZN(n4384) );
  INV_X1 U5744 ( .A(n4380), .ZN(n4381) );
  NOR2_X1 U5745 ( .A1(n4381), .A2(pmp_addr_i[98]), .ZN(n4382) );
  NOR2_X1 U5746 ( .A1(n5291), .A2(n4382), .ZN(n4383) );
  NOR3_X1 U5747 ( .A1(n4387), .A2(n4384), .A3(n4383), .ZN(n4393) );
  NAND2_X1 U5748 ( .A1(n5293), .A2(n4762), .ZN(n4386) );
  AOI22_X1 U5749 ( .A1(instr_addr_o_6_), .A2(n4763), .B1(n5740), .B2(n4776), 
        .ZN(n4385) );
  NAND2_X1 U5750 ( .A1(n5269), .A2(n4780), .ZN(n4390) );
  OAI211_X1 U5751 ( .C1(n4387), .C2(n4386), .A(n4385), .B(n4390), .ZN(n4392)
         );
  NAND2_X1 U5752 ( .A1(n5262), .A2(n4196), .ZN(n4398) );
  NOR2_X1 U5753 ( .A1(n12267), .A2(n4776), .ZN(n4389) );
  AOI22_X1 U5754 ( .A1(n4390), .A2(n4389), .B1(n4606), .B2(pmp_addr_i[102]), 
        .ZN(n4391) );
  OAI211_X1 U5755 ( .C1(n4393), .C2(n4392), .A(n4400), .B(n4391), .ZN(n4404)
         );
  OAI21_X1 U5756 ( .B1(n5052), .B2(pmp_addr_i[105]), .A(n4394), .ZN(n4395) );
  NOR2_X1 U5757 ( .A1(n4396), .A2(n4395), .ZN(n4402) );
  NAND2_X1 U5758 ( .A1(instr_addr_o_9_), .A2(n4782), .ZN(n4397) );
  NAND2_X1 U5759 ( .A1(n4398), .A2(n4397), .ZN(n4399) );
  NAND2_X1 U5760 ( .A1(n4400), .A2(n4399), .ZN(n4401) );
  NAND4_X1 U5761 ( .A1(n4404), .A2(n4403), .A3(n4402), .A4(n4401), .ZN(n4415)
         );
  NAND2_X1 U5762 ( .A1(n210), .A2(n1184), .ZN(n4431) );
  NAND2_X1 U5763 ( .A1(n136), .A2(n1182), .ZN(n4405) );
  NAND2_X1 U5764 ( .A1(n4431), .A2(n4405), .ZN(n4433) );
  NOR2_X1 U5765 ( .A1(n4418), .A2(n4433), .ZN(n4413) );
  INV_X1 U5766 ( .A(pmp_addr_i[125]), .ZN(n4407) );
  NAND2_X1 U5767 ( .A1(n5187), .A2(n1175), .ZN(n4419) );
  OAI211_X1 U5768 ( .C1(n5313), .C2(pmp_addr_i[113]), .A(n4442), .B(n4419), 
        .ZN(n4408) );
  NOR2_X1 U5769 ( .A1(n4437), .A2(n4408), .ZN(n4412) );
  NAND2_X1 U5770 ( .A1(n5191), .A2(n1167), .ZN(n4409) );
  NAND2_X1 U5771 ( .A1(n5181), .A2(n1169), .ZN(n4421) );
  NAND2_X1 U5772 ( .A1(n4409), .A2(n4421), .ZN(n4424) );
  NAND2_X1 U5773 ( .A1(instr_addr_o_24_), .A2(n1188), .ZN(n4428) );
  NAND2_X1 U5774 ( .A1(instr_addr_o_23_), .A2(n1180), .ZN(n4410) );
  AND2_X1 U5775 ( .A1(n4428), .A2(n4410), .ZN(n4426) );
  NAND4_X1 U5776 ( .A1(n4413), .A2(n4412), .A3(n4411), .A4(n4426), .ZN(n4414)
         );
  AOI21_X1 U5777 ( .B1(n4416), .B2(n4415), .A(n4414), .ZN(n4452) );
  INV_X1 U5778 ( .A(n4442), .ZN(n4417) );
  INV_X1 U5779 ( .A(n4433), .ZN(n4427) );
  AOI22_X1 U5780 ( .A1(n4420), .A2(n4419), .B1(n2569), .B2(pmp_addr_i[114]), 
        .ZN(n4425) );
  NOR2_X1 U5781 ( .A1(n5842), .A2(n1167), .ZN(n4422) );
  AOI22_X1 U5782 ( .A1(n4422), .A2(n4421), .B1(n5192), .B2(pmp_addr_i[116]), 
        .ZN(n4423) );
  NOR2_X1 U5783 ( .A1(n4859), .A2(n1180), .ZN(n4429) );
  AOI22_X1 U5784 ( .A1(n4429), .A2(n4428), .B1(pmp_addr_i[118]), .B2(n1269), 
        .ZN(n4434) );
  NOR2_X1 U5785 ( .A1(n4644), .A2(n1182), .ZN(n4430) );
  AOI22_X1 U5786 ( .A1(n4431), .A2(n4430), .B1(n3806), .B2(pmp_addr_i[120]), 
        .ZN(n4432) );
  OAI21_X1 U5787 ( .B1(n4434), .B2(n4433), .A(n4432), .ZN(n4435) );
  NOR2_X1 U5788 ( .A1(n4437), .A2(n4417), .ZN(n4447) );
  NAND2_X1 U5789 ( .A1(n4438), .A2(pmp_addr_i[122]), .ZN(n4439) );
  NAND2_X1 U5790 ( .A1(n4440), .A2(n4439), .ZN(n4446) );
  NAND2_X1 U5791 ( .A1(n4660), .A2(pmp_addr_i[125]), .ZN(n4443) );
  AOI21_X1 U5792 ( .B1(n4447), .B2(n4446), .A(n4445), .ZN(n4448) );
  NAND3_X1 U5793 ( .A1(n4450), .A2(n4449), .A3(n4448), .ZN(n4451) );
  NOR2_X1 U5794 ( .A1(n4560), .A2(n9896), .ZN(n4563) );
  NOR2_X1 U5795 ( .A1(n4900), .A2(n9895), .ZN(n4454) );
  NOR2_X1 U5796 ( .A1(n4563), .A2(n4454), .ZN(n4566) );
  NOR2_X1 U5797 ( .A1(n4556), .A2(n9887), .ZN(n4455) );
  NOR2_X1 U5798 ( .A1(n5368), .A2(n9888), .ZN(n4559) );
  NOR2_X1 U5799 ( .A1(n4455), .A2(n4559), .ZN(n4456) );
  NAND2_X1 U5800 ( .A1(n4566), .A2(n4456), .ZN(n4461) );
  INV_X1 U5801 ( .A(n9964), .ZN(n4567) );
  NOR2_X1 U5802 ( .A1(instr_addr_o_31_), .A2(n4567), .ZN(n4458) );
  INV_X1 U5803 ( .A(pmp_addr_i[414]), .ZN(n4457) );
  NOR2_X1 U5804 ( .A1(n4458), .A2(pmp_addr_i[414]), .ZN(n4460) );
  INV_X1 U5805 ( .A(pmp_addr_i[415]), .ZN(n4459) );
  NAND2_X1 U5806 ( .A1(n4460), .A2(n4459), .ZN(n4571) );
  NOR2_X1 U5807 ( .A1(n4461), .A2(n4571), .ZN(n4554) );
  INV_X1 U5808 ( .A(n9936), .ZN(n4529) );
  NOR2_X1 U5809 ( .A1(n4907), .A2(n9847), .ZN(n4462) );
  NOR2_X1 U5810 ( .A1(n4532), .A2(n4462), .ZN(n4464) );
  NOR2_X1 U5811 ( .A1(n5181), .A2(n9855), .ZN(n4536) );
  NOR2_X1 U5812 ( .A1(n4533), .A2(n9854), .ZN(n4463) );
  NOR2_X1 U5813 ( .A1(n4536), .A2(n4463), .ZN(n4539) );
  NAND2_X1 U5814 ( .A1(n4464), .A2(n4539), .ZN(n4468) );
  NOR2_X1 U5815 ( .A1(instr_addr_o_24_), .A2(n9860), .ZN(n4543) );
  NOR2_X1 U5816 ( .A1(n4859), .A2(n9859), .ZN(n4465) );
  NOR2_X1 U5817 ( .A1(n4543), .A2(n4465), .ZN(n4467) );
  NOR2_X1 U5818 ( .A1(n4909), .A2(n9882), .ZN(n4547) );
  NOR2_X1 U5819 ( .A1(n136), .A2(n9881), .ZN(n4466) );
  NOR2_X1 U5820 ( .A1(n4547), .A2(n4466), .ZN(n4550) );
  NAND2_X1 U5821 ( .A1(n4467), .A2(n4550), .ZN(n4552) );
  NOR2_X1 U5822 ( .A1(n4468), .A2(n4552), .ZN(n4469) );
  NAND2_X1 U5823 ( .A1(n4554), .A2(n4469), .ZN(n4577) );
  AND2_X1 U5824 ( .A1(n5023), .A2(n9790), .ZN(n4475) );
  NOR2_X1 U5825 ( .A1(n5291), .A2(n9974), .ZN(n4472) );
  INV_X1 U5826 ( .A(n9784), .ZN(n9967) );
  INV_X1 U5827 ( .A(n9783), .ZN(n9973) );
  NAND2_X1 U5828 ( .A1(n9967), .A2(n9973), .ZN(n4471) );
  NAND2_X1 U5829 ( .A1(n5291), .A2(n9974), .ZN(n4470) );
  NAND2_X1 U5830 ( .A1(n20), .A2(n9971), .ZN(n4474) );
  NOR2_X1 U5831 ( .A1(n5342), .A2(n9979), .ZN(n4482) );
  NOR2_X1 U5832 ( .A1(n5268), .A2(n4476), .ZN(n4477) );
  NOR2_X1 U5833 ( .A1(n4482), .A2(n4477), .ZN(n4479) );
  NOR2_X1 U5834 ( .A1(n214), .A2(n9966), .ZN(n4485) );
  NOR2_X1 U5835 ( .A1(n4485), .A2(n4478), .ZN(n4488) );
  NAND2_X1 U5836 ( .A1(n4479), .A2(n4488), .ZN(n4490) );
  NAND2_X1 U5837 ( .A1(n5342), .A2(n9979), .ZN(n4480) );
  OAI21_X1 U5838 ( .B1(n4482), .B2(n4481), .A(n4480), .ZN(n4487) );
  NAND2_X1 U5839 ( .A1(instr_addr_o_10_), .A2(n9966), .ZN(n4483) );
  OAI21_X1 U5840 ( .B1(n4485), .B2(n4484), .A(n4483), .ZN(n4486) );
  AOI21_X1 U5841 ( .B1(n4488), .B2(n4487), .A(n4486), .ZN(n4489) );
  OAI21_X1 U5842 ( .B1(n4491), .B2(n4490), .A(n4489), .ZN(n4528) );
  NOR2_X1 U5843 ( .A1(n4061), .A2(n9982), .ZN(n4492) );
  NOR2_X1 U5844 ( .A1(n4508), .A2(n4492), .ZN(n4511) );
  NOR2_X1 U5845 ( .A1(n3934), .A2(n9965), .ZN(n4495) );
  NOR2_X1 U5846 ( .A1(n4494), .A2(n9983), .ZN(n4505) );
  NOR2_X1 U5847 ( .A1(n4495), .A2(n12214), .ZN(n4496) );
  NAND2_X1 U5848 ( .A1(n4511), .A2(n4496), .ZN(n4502) );
  NOR2_X1 U5849 ( .A1(n4498), .A2(n4497), .ZN(n4499) );
  NOR2_X1 U5850 ( .A1(n4743), .A2(n9986), .ZN(n4515) );
  NOR2_X1 U5851 ( .A1(n4499), .A2(n4515), .ZN(n4501) );
  NOR2_X1 U5852 ( .A1(n4500), .A2(n4519), .ZN(n4522) );
  NAND2_X1 U5853 ( .A1(n4501), .A2(n4522), .ZN(n4524) );
  NOR2_X1 U5854 ( .A1(n4502), .A2(n4524), .ZN(n4527) );
  OAI21_X1 U5855 ( .B1(n4505), .B2(n4504), .A(n4503), .ZN(n4510) );
  OAI21_X1 U5856 ( .B1(n4508), .B2(n4507), .A(n4506), .ZN(n4509) );
  AOI21_X1 U5857 ( .B1(n4511), .B2(n4510), .A(n4509), .ZN(n4525) );
  NAND2_X1 U5858 ( .A1(n12266), .A2(n9986), .ZN(n4513) );
  OAI21_X1 U5859 ( .B1(n4515), .B2(n4514), .A(n4513), .ZN(n4521) );
  OAI21_X1 U5860 ( .B1(n4519), .B2(n4518), .A(n4517), .ZN(n4520) );
  AOI21_X1 U5861 ( .B1(n4521), .B2(n4522), .A(n4520), .ZN(n4523) );
  OAI21_X1 U5862 ( .B1(n4525), .B2(n4524), .A(n4523), .ZN(n4526) );
  AOI21_X1 U5863 ( .B1(n4528), .B2(n4527), .A(n4526), .ZN(n4576) );
  NAND2_X1 U5864 ( .A1(n3793), .A2(n9847), .ZN(n4531) );
  NAND2_X1 U5865 ( .A1(n6027), .A2(n4529), .ZN(n4530) );
  OAI21_X1 U5866 ( .B1(n4532), .B2(n4531), .A(n4530), .ZN(n4538) );
  NAND2_X1 U5867 ( .A1(n4533), .A2(n9854), .ZN(n4535) );
  NAND2_X1 U5868 ( .A1(n4836), .A2(n9855), .ZN(n4534) );
  OAI21_X1 U5869 ( .B1(n4536), .B2(n4535), .A(n4534), .ZN(n4537) );
  AOI21_X1 U5870 ( .B1(n4539), .B2(n4538), .A(n4537), .ZN(n4553) );
  NAND2_X1 U5871 ( .A1(n4859), .A2(n9859), .ZN(n4542) );
  NAND2_X1 U5872 ( .A1(instr_addr_o_24_), .A2(n9860), .ZN(n4541) );
  OAI21_X1 U5873 ( .B1(n4543), .B2(n4542), .A(n4541), .ZN(n4549) );
  NAND2_X1 U5874 ( .A1(n136), .A2(n9881), .ZN(n4546) );
  NAND2_X1 U5875 ( .A1(n4909), .A2(n9882), .ZN(n4545) );
  OAI21_X1 U5876 ( .B1(n4547), .B2(n4546), .A(n4545), .ZN(n4548) );
  AOI21_X1 U5877 ( .B1(n4550), .B2(n4549), .A(n4548), .ZN(n4551) );
  OAI21_X1 U5878 ( .B1(n4553), .B2(n4552), .A(n4551), .ZN(n4555) );
  NAND2_X1 U5879 ( .A1(n4555), .A2(n4554), .ZN(n4575) );
  NAND2_X1 U5880 ( .A1(n4556), .A2(n9887), .ZN(n4558) );
  NAND2_X1 U5881 ( .A1(instr_addr_o_28_), .A2(n9888), .ZN(n4557) );
  OAI21_X1 U5882 ( .B1(n4559), .B2(n4558), .A(n4557), .ZN(n4565) );
  NAND2_X1 U5883 ( .A1(n4900), .A2(n9895), .ZN(n4562) );
  NAND2_X1 U5884 ( .A1(n4560), .A2(n9896), .ZN(n4561) );
  OAI21_X1 U5885 ( .B1(n4563), .B2(n4562), .A(n4561), .ZN(n4564) );
  AOI21_X1 U5886 ( .B1(n4566), .B2(n4565), .A(n4564), .ZN(n4572) );
  NAND2_X1 U5887 ( .A1(n6018), .A2(n4567), .ZN(n4568) );
  NOR2_X1 U5888 ( .A1(n4568), .A2(pmp_addr_i[414]), .ZN(n4569) );
  NAND2_X1 U5889 ( .A1(n4569), .A2(n4459), .ZN(n4570) );
  OAI21_X1 U5890 ( .B1(n4572), .B2(n4571), .A(n4570), .ZN(n4573) );
  INV_X1 U5891 ( .A(n4573), .ZN(n4574) );
  OAI211_X1 U5892 ( .C1(n4576), .C2(n4577), .A(n4575), .B(n4574), .ZN(n4668)
         );
  OAI21_X1 U5893 ( .B1(n5048), .B2(pmp_addr_i[431]), .A(n4590), .ZN(n4592) );
  NAND2_X1 U5894 ( .A1(n4743), .A2(n3507), .ZN(n4588) );
  OAI21_X1 U5895 ( .B1(n4578), .B2(pmp_addr_i[429]), .A(n4588), .ZN(n4579) );
  NOR2_X1 U5896 ( .A1(n4592), .A2(n4579), .ZN(n4619) );
  NAND2_X1 U5897 ( .A1(n5250), .A2(n3538), .ZN(n4612) );
  NOR2_X1 U5898 ( .A1(n4493), .A2(n3499), .ZN(n4580) );
  AOI22_X1 U5899 ( .A1(n4612), .A2(n4580), .B1(n5070), .B2(pmp_addr_i[426]), 
        .ZN(n4586) );
  NAND2_X1 U5900 ( .A1(n4788), .A2(n3501), .ZN(n4584) );
  INV_X1 U5901 ( .A(pmp_addr_i[427]), .ZN(n4582) );
  NAND2_X1 U5902 ( .A1(instr_addr_o_13_), .A2(n4582), .ZN(n4581) );
  NAND2_X1 U5903 ( .A1(n4584), .A2(n4581), .ZN(n4614) );
  NOR2_X1 U5904 ( .A1(n5997), .A2(n4582), .ZN(n4583) );
  AOI22_X1 U5905 ( .A1(n4584), .A2(n4583), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[428]), .ZN(n4585) );
  NOR2_X1 U5906 ( .A1(n4498), .A2(n3533), .ZN(n4587) );
  AOI22_X1 U5907 ( .A1(n4588), .A2(n4587), .B1(n5058), .B2(pmp_addr_i[430]), 
        .ZN(n4593) );
  AND2_X1 U5908 ( .A1(n4234), .A2(pmp_addr_i[431]), .ZN(n4589) );
  AOI22_X1 U5909 ( .A1(n4590), .A2(n4589), .B1(instr_addr_o_18__BAR), .B2(
        pmp_addr_i[432]), .ZN(n4591) );
  NOR2_X1 U5910 ( .A1(n5277), .A2(n2408), .ZN(n4601) );
  NAND2_X1 U5911 ( .A1(instr_addr_o_5_), .A2(n3514), .ZN(n4595) );
  INV_X1 U5912 ( .A(pmp_addr_i[421]), .ZN(n4604) );
  AOI22_X1 U5913 ( .A1(instr_addr_o_6_), .A2(n2408), .B1(n5740), .B2(n4604), 
        .ZN(n4594) );
  NAND2_X1 U5914 ( .A1(n5269), .A2(n3505), .ZN(n4608) );
  OAI211_X1 U5915 ( .C1(n4601), .C2(n4595), .A(n4594), .B(n4608), .ZN(n4611)
         );
  NOR2_X1 U5916 ( .A1(pmp_addr_i[417]), .A2(pmp_addr_i[416]), .ZN(n4597) );
  OAI22_X1 U5917 ( .A1(n20), .A2(n3514), .B1(n4597), .B2(n3497), .ZN(n4600) );
  AND2_X1 U5918 ( .A1(n4597), .A2(n3497), .ZN(n4598) );
  NOR2_X1 U5919 ( .A1(n5291), .A2(n4598), .ZN(n4599) );
  NOR3_X1 U5920 ( .A1(n4601), .A2(n4600), .A3(n4599), .ZN(n4610) );
  NOR2_X1 U5921 ( .A1(n153), .A2(n3549), .ZN(n4603) );
  NAND2_X1 U5922 ( .A1(n5262), .A2(n3522), .ZN(n4616) );
  NOR2_X1 U5924 ( .A1(n12267), .A2(n4604), .ZN(n4607) );
  AOI22_X1 U5925 ( .A1(n4608), .A2(n4607), .B1(n4606), .B2(pmp_addr_i[422]), 
        .ZN(n4609) );
  OAI21_X1 U5926 ( .B1(n5052), .B2(pmp_addr_i[425]), .A(n4612), .ZN(n4613) );
  NOR2_X1 U5927 ( .A1(n4614), .A2(n4613), .ZN(n4620) );
  NAND2_X1 U5928 ( .A1(instr_addr_o_9_), .A2(n3549), .ZN(n4615) );
  NAND2_X1 U5929 ( .A1(n210), .A2(n2481), .ZN(n4646) );
  NAND2_X1 U5930 ( .A1(n12226), .A2(n2484), .ZN(n4621) );
  NOR2_X1 U5931 ( .A1(n4640), .A2(n4648), .ZN(n4629) );
  NAND2_X1 U5932 ( .A1(n12263), .A2(n2503), .ZN(n4657) );
  OAI21_X1 U5933 ( .B1(n4623), .B2(pmp_addr_i[443]), .A(n4657), .ZN(n4651) );
  NAND2_X1 U5934 ( .A1(n4802), .A2(n2498), .ZN(n4632) );
  OAI211_X1 U5935 ( .C1(n12208), .C2(pmp_addr_i[433]), .A(n4659), .B(n4632), 
        .ZN(n4624) );
  NOR2_X1 U5936 ( .A1(n4651), .A2(n4624), .ZN(n4628) );
  NAND2_X1 U5937 ( .A1(n5191), .A2(n2495), .ZN(n4625) );
  NAND2_X1 U5938 ( .A1(n5181), .A2(n2493), .ZN(n4634) );
  NAND2_X1 U5939 ( .A1(n4625), .A2(n4634), .ZN(n4637) );
  NAND2_X1 U5940 ( .A1(instr_addr_o_24_), .A2(n2489), .ZN(n4643) );
  NAND2_X1 U5941 ( .A1(instr_addr_o_23_), .A2(n2487), .ZN(n4626) );
  AND2_X1 U5942 ( .A1(n4643), .A2(n4626), .ZN(n4641) );
  NAND4_X1 U5943 ( .A1(n4629), .A2(n4628), .A3(n4627), .A4(n4641), .ZN(n4630)
         );
  AOI22_X1 U5944 ( .A1(n4633), .A2(n4632), .B1(n4631), .B2(pmp_addr_i[434]), 
        .ZN(n4638) );
  NOR2_X1 U5945 ( .A1(n5842), .A2(n2495), .ZN(n4635) );
  AOI22_X1 U5946 ( .A1(n4635), .A2(n4634), .B1(n999), .B2(pmp_addr_i[436]), 
        .ZN(n4636) );
  INV_X1 U5947 ( .A(n4659), .ZN(n4639) );
  AOI22_X1 U5948 ( .A1(n4643), .A2(n4642), .B1(n2580), .B2(pmp_addr_i[438]), 
        .ZN(n4649) );
  NOR2_X1 U5949 ( .A1(n4644), .A2(n2484), .ZN(n4645) );
  AOI22_X1 U5950 ( .A1(n4646), .A2(n4645), .B1(n1273), .B2(pmp_addr_i[440]), 
        .ZN(n4647) );
  OAI21_X1 U5951 ( .B1(n4649), .B2(n4648), .A(n4647), .ZN(n4650) );
  NOR2_X1 U5952 ( .A1(n4651), .A2(n4639), .ZN(n4666) );
  NAND3_X1 U5953 ( .A1(n4653), .A2(pmp_addr_i[441]), .A3(n4652), .ZN(n4655) );
  NAND2_X1 U5954 ( .A1(n5111), .A2(pmp_addr_i[442]), .ZN(n4654) );
  NAND2_X1 U5955 ( .A1(n4655), .A2(n4654), .ZN(n4665) );
  NAND4_X1 U5956 ( .A1(n4657), .A2(n4659), .A3(pmp_addr_i[443]), .A4(n4656), 
        .ZN(n4663) );
  NAND3_X1 U5957 ( .A1(n4659), .A2(pmp_addr_i[444]), .A3(n4658), .ZN(n4662) );
  NAND2_X1 U5958 ( .A1(n4660), .A2(pmp_addr_i[445]), .ZN(n4661) );
  NAND4_X1 U5959 ( .A1(n4663), .A2(n9764), .A3(n4662), .A4(n4661), .ZN(n4664)
         );
  NAND3_X1 U5960 ( .A1(n5269), .A2(n3909), .A3(n11779), .ZN(n4670) );
  NAND3_X1 U5961 ( .A1(n5040), .A2(n6654), .A3(n11769), .ZN(n4669) );
  OAI211_X1 U5962 ( .C1(n4703), .C2(n11790), .A(n4670), .B(n4669), .ZN(n4680)
         );
  INV_X1 U5963 ( .A(pmp_addr_i[487]), .ZN(n11761) );
  NOR2_X1 U5964 ( .A1(n6525), .A2(n4671), .ZN(n4672) );
  NAND2_X1 U5965 ( .A1(instr_addr_o_10_), .A2(n4672), .ZN(n4678) );
  NAND3_X1 U5966 ( .A1(n12150), .A2(n6674), .A3(n3877), .ZN(n4677) );
  INV_X1 U5967 ( .A(n4673), .ZN(n11784) );
  NAND3_X1 U5968 ( .A1(instr_addr_o_5_), .A2(n3887), .A3(n11784), .ZN(n4676)
         );
  OR2_X1 U5969 ( .A1(n4674), .A2(n6624), .ZN(n6695) );
  NAND2_X1 U5970 ( .A1(n6695), .A2(pmp_cfg_i[122]), .ZN(n4690) );
  NAND2_X1 U5971 ( .A1(pmp_cfg_i[124]), .A2(pmp_cfg_i[123]), .ZN(n11796) );
  NOR2_X1 U5972 ( .A1(n4690), .A2(n11796), .ZN(n4675) );
  AND2_X1 U5973 ( .A1(n6002), .A2(n3955), .ZN(n4696) );
  INV_X1 U5974 ( .A(n4681), .ZN(n11781) );
  AND2_X1 U5975 ( .A1(n5251), .A2(n4733), .ZN(n4700) );
  AOI22_X1 U5976 ( .A1(n4696), .A2(n11781), .B1(n4700), .B2(n11762), .ZN(n4683) );
  AND2_X1 U5977 ( .A1(n12266), .A2(n3965), .ZN(n4701) );
  INV_X1 U5978 ( .A(n6528), .ZN(n6683) );
  AND2_X1 U5979 ( .A1(n5245), .A2(n6683), .ZN(n4702) );
  NAND2_X1 U5980 ( .A1(n4681), .A2(pmp_addr_i[489]), .ZN(n11802) );
  AOI22_X1 U5981 ( .A1(n4701), .A2(n11807), .B1(n4702), .B2(n11802), .ZN(n4682) );
  INV_X1 U5982 ( .A(n4684), .ZN(n11805) );
  NOR2_X1 U5983 ( .A1(n11802), .A2(n4685), .ZN(n11789) );
  OAI22_X1 U5984 ( .A1(n11805), .A2(n4694), .B1(n4698), .B2(n11789), .ZN(n4688) );
  INV_X1 U5985 ( .A(n11785), .ZN(n4686) );
  NOR2_X1 U5986 ( .A1(n11785), .A2(n4083), .ZN(n11765) );
  OAI22_X1 U5987 ( .A1(n4686), .A2(n4697), .B1(n4699), .B2(n11765), .ZN(n4687)
         );
  AOI22_X1 U5988 ( .A1(n155), .A2(n6654), .B1(n205), .B2(n3909), .ZN(n4695) );
  AOI22_X1 U5989 ( .A1(n12202), .A2(n3912), .B1(n5899), .B2(n6674), .ZN(n4693)
         );
  OR2_X1 U5990 ( .A1(n4690), .A2(pmp_cfg_i[123]), .ZN(n4691) );
  AOI21_X1 U5991 ( .B1(n6015), .B2(n3887), .A(n4691), .ZN(n4692) );
  NAND4_X1 U5992 ( .A1(n4695), .A2(n4694), .A3(n4693), .A4(n4692), .ZN(n4706)
         );
  NAND4_X1 U5993 ( .A1(n4699), .A2(n4698), .A3(n4697), .A4(n3957), .ZN(n4705)
         );
  NOR3_X1 U5994 ( .A1(n4706), .A2(n4705), .A3(n4704), .ZN(n4739) );
  OAI211_X1 U5995 ( .C1(n5293), .C2(n3887), .A(n6677), .B(n323), .ZN(n4707) );
  NOR2_X1 U5996 ( .A1(n4708), .A2(n4707), .ZN(n4712) );
  XNOR2_X1 U5997 ( .A(n4908), .B(n6648), .ZN(n4711) );
  XNOR2_X1 U5998 ( .A(n4907), .B(n6644), .ZN(n4710) );
  XNOR2_X1 U5999 ( .A(n6018), .B(n6671), .ZN(n4709) );
  NAND4_X1 U6000 ( .A1(n4712), .A2(n4711), .A3(n4710), .A4(n4709), .ZN(n4718)
         );
  XNOR2_X1 U6001 ( .A(n5985), .B(n6635), .ZN(n4716) );
  XNOR2_X1 U6002 ( .A(n5550), .B(n6664), .ZN(n4715) );
  XNOR2_X1 U6003 ( .A(instr_addr_o_25_), .B(n6634), .ZN(n4714) );
  XNOR2_X1 U6004 ( .A(instr_addr_o_21_), .B(n6626), .ZN(n4713) );
  NAND4_X1 U6005 ( .A1(n4716), .A2(n4715), .A3(n4714), .A4(n4713), .ZN(n4717)
         );
  NOR2_X1 U6006 ( .A1(n4718), .A2(n4717), .ZN(n4738) );
  OAI22_X1 U6007 ( .A1(n5245), .A2(n6683), .B1(n5974), .B2(n4719), .ZN(n4721)
         );
  OAI22_X1 U6008 ( .A1(n12202), .A2(n3912), .B1(n5976), .B2(n6674), .ZN(n4720)
         );
  NOR2_X1 U6009 ( .A1(n4721), .A2(n4720), .ZN(n4725) );
  XNOR2_X1 U6010 ( .A(n4753), .B(n6637), .ZN(n4724) );
  XNOR2_X1 U6011 ( .A(instr_addr_o_27_), .B(n6663), .ZN(n4723) );
  XNOR2_X1 U6012 ( .A(n4901), .B(n6636), .ZN(n4722) );
  NAND4_X1 U6013 ( .A1(n4725), .A2(n4724), .A3(n4723), .A4(n4722), .ZN(n4737)
         );
  XNOR2_X1 U6014 ( .A(n4859), .B(n6628), .ZN(n4729) );
  XNOR2_X1 U6015 ( .A(n4836), .B(n6627), .ZN(n4728) );
  XNOR2_X1 U6016 ( .A(n4835), .B(n6629), .ZN(n4727) );
  XNOR2_X1 U6017 ( .A(n6027), .B(n6645), .ZN(n4726) );
  INV_X1 U6018 ( .A(n6533), .ZN(n4730) );
  OAI22_X1 U6019 ( .A1(n5997), .A2(n3959), .B1(n12179), .B2(n4730), .ZN(n4732)
         );
  OAI22_X1 U6020 ( .A1(instr_addr_o_6_), .A2(n3888), .B1(n12267), .B2(n3908), 
        .ZN(n4731) );
  NOR2_X1 U6021 ( .A1(n4732), .A2(n4731), .ZN(n4736) );
  OAI22_X1 U6022 ( .A1(n6002), .A2(n3955), .B1(n5251), .B2(n4733), .ZN(n4735)
         );
  OAI22_X1 U6023 ( .A1(n6005), .A2(n3909), .B1(n5229), .B2(n3965), .ZN(n4734)
         );
  AND2_X1 U6024 ( .A1(n4740), .A2(n4794), .ZN(n4747) );
  OR2_X1 U6025 ( .A1(n4741), .A2(n7551), .ZN(n7619) );
  AND2_X1 U6026 ( .A1(n7619), .A2(pmp_cfg_i[26]), .ZN(n4768) );
  NAND2_X1 U6027 ( .A1(n4768), .A2(n7604), .ZN(n4742) );
  AOI21_X1 U6028 ( .B1(n12156), .B2(n4251), .A(n4742), .ZN(n4746) );
  INV_X1 U6029 ( .A(n7320), .ZN(n7556) );
  AOI22_X1 U6030 ( .A1(n12181), .A2(n4807), .B1(n12266), .B2(n7556), .ZN(n4745) );
  NAND4_X1 U6031 ( .A1(n4747), .A2(n4746), .A3(n4745), .A4(n4744), .ZN(n4752)
         );
  NAND4_X1 U6032 ( .A1(n4766), .A2(n4765), .A3(n4779), .A4(n4778), .ZN(n4751)
         );
  NAND4_X1 U6033 ( .A1(n4749), .A2(n4748), .A3(n4785), .A4(n4791), .ZN(n4750)
         );
  NOR3_X1 U6034 ( .A1(n4752), .A2(n4751), .A3(n4750), .ZN(n4758) );
  XNOR2_X1 U6035 ( .A(n4753), .B(n7578), .ZN(n4757) );
  XNOR2_X1 U6036 ( .A(n138), .B(n7577), .ZN(n4756) );
  XNOR2_X1 U6037 ( .A(n4900), .B(n7603), .ZN(n4755) );
  XNOR2_X1 U6038 ( .A(n5154), .B(n7614), .ZN(n4754) );
  AND4_X1 U6039 ( .A1(n4755), .A2(n4756), .A3(n4757), .A4(n4754), .ZN(n4800)
         );
  INV_X1 U6041 ( .A(n4759), .ZN(n4760) );
  NAND2_X1 U6042 ( .A1(n4761), .A2(n4760), .ZN(n11728) );
  OR2_X1 U6043 ( .A1(n11728), .A2(n4762), .ZN(n11736) );
  NOR2_X1 U6044 ( .A1(n11736), .A2(n4763), .ZN(n11749) );
  INV_X1 U6045 ( .A(n11730), .ZN(n4764) );
  OAI22_X1 U6046 ( .A1(n11749), .A2(n4766), .B1(n4765), .B2(n4764), .ZN(n4775)
         );
  NAND2_X1 U6047 ( .A1(n11701), .A2(pmp_addr_i[109]), .ZN(n11708) );
  NOR2_X1 U6048 ( .A1(n11708), .A2(n4767), .ZN(n11707) );
  NOR2_X1 U6049 ( .A1(n7322), .A2(n11707), .ZN(n4770) );
  INV_X1 U6050 ( .A(n4768), .ZN(n4769) );
  AOI21_X1 U6051 ( .B1(n12265), .B2(n4770), .A(n4769), .ZN(n4773) );
  INV_X1 U6052 ( .A(n7328), .ZN(n7564) );
  NOR2_X1 U6053 ( .A1(n11730), .A2(n4771), .ZN(n11713) );
  NAND2_X1 U6054 ( .A1(n11713), .A2(pmp_addr_i[106]), .ZN(n11710) );
  NAND3_X1 U6055 ( .A1(instr_addr_o_13_), .A2(n7564), .A3(n11710), .ZN(n4772)
         );
  OAI211_X1 U6056 ( .C1(n4744), .C2(n11701), .A(n4773), .B(n4772), .ZN(n4774)
         );
  NOR2_X1 U6057 ( .A1(n4775), .A2(n4774), .ZN(n4799) );
  INV_X1 U6058 ( .A(n11749), .ZN(n4777) );
  NOR2_X1 U6059 ( .A1(n4777), .A2(n4776), .ZN(n11722) );
  INV_X1 U6060 ( .A(n11722), .ZN(n4781) );
  OR2_X1 U6061 ( .A1(n4781), .A2(n4780), .ZN(n11751) );
  NOR2_X1 U6062 ( .A1(n11751), .A2(n4782), .ZN(n11746) );
  NAND3_X1 U6063 ( .A1(n5040), .A2(n4203), .A3(n11751), .ZN(n4784) );
  NAND3_X1 U6064 ( .A1(instr_addr_o_6_), .A2(n7563), .A3(n11736), .ZN(n4783)
         );
  OAI211_X1 U6065 ( .C1(n4785), .C2(n11746), .A(n4784), .B(n4783), .ZN(n4786)
         );
  INV_X1 U6066 ( .A(n4787), .ZN(n11727) );
  OR2_X1 U6067 ( .A1(n11710), .A2(n4366), .ZN(n11704) );
  NAND3_X1 U6068 ( .A1(n206), .A2(n4807), .A3(n11704), .ZN(n4790) );
  NAND3_X1 U6069 ( .A1(n5229), .A2(n7556), .A3(n11708), .ZN(n4789) );
  OAI211_X1 U6070 ( .C1(n4791), .C2(n11727), .A(n4790), .B(n4789), .ZN(n4796)
         );
  INV_X1 U6071 ( .A(n4792), .ZN(n11733) );
  INV_X1 U6072 ( .A(n11728), .ZN(n4793) );
  AOI21_X1 U6073 ( .B1(n4794), .B2(n11733), .A(n4793), .ZN(n4795) );
  NOR2_X1 U6074 ( .A1(n4796), .A2(n4795), .ZN(n4797) );
  XNOR2_X1 U6075 ( .A(n4859), .B(n7586), .ZN(n4806) );
  XNOR2_X1 U6076 ( .A(n12157), .B(n7585), .ZN(n4805) );
  XNOR2_X1 U6077 ( .A(instr_addr_o_20_), .B(n7583), .ZN(n4804) );
  XNOR2_X1 U6078 ( .A(n4835), .B(n7591), .ZN(n4803) );
  AND4_X1 U6079 ( .A1(n4806), .A2(n4805), .A3(n4804), .A4(n4803), .ZN(n4815)
         );
  OAI22_X1 U6080 ( .A1(n5069), .A2(n7360), .B1(n12180), .B2(n4807), .ZN(n4809)
         );
  OAI22_X1 U6081 ( .A1(n6005), .A2(n4201), .B1(n12266), .B2(n7556), .ZN(n4808)
         );
  NOR2_X1 U6082 ( .A1(n4809), .A2(n4808), .ZN(n4814) );
  OAI22_X1 U6083 ( .A1(n5997), .A2(n7564), .B1(n12179), .B2(n4810), .ZN(n4812)
         );
  OAI22_X1 U6084 ( .A1(instr_addr_o_6_), .A2(n7563), .B1(n4605), .B2(n7557), 
        .ZN(n4811) );
  NOR2_X1 U6085 ( .A1(n4812), .A2(n4811), .ZN(n4813) );
  NAND3_X1 U6086 ( .A1(n4815), .A2(n4814), .A3(n4813), .ZN(n4831) );
  OAI22_X1 U6087 ( .A1(n5245), .A2(n4242), .B1(n4069), .B2(n4251), .ZN(n4818)
         );
  OAI22_X1 U6088 ( .A1(n12202), .A2(n4205), .B1(n5976), .B2(n4816), .ZN(n4817)
         );
  NOR2_X1 U6089 ( .A1(n4818), .A2(n4817), .ZN(n4822) );
  XNOR2_X1 U6090 ( .A(instr_addr_o_25_), .B(n7592), .ZN(n4821) );
  XNOR2_X1 U6091 ( .A(n5985), .B(n7593), .ZN(n4820) );
  XNOR2_X1 U6092 ( .A(instr_addr_o_27_), .B(n7594), .ZN(n4819) );
  NAND4_X1 U6093 ( .A1(n4822), .A2(n4821), .A3(n4820), .A4(n4819), .ZN(n4830)
         );
  OAI211_X1 U6094 ( .C1(n5293), .C2(n4182), .A(n7606), .B(n157), .ZN(n4823) );
  NOR2_X1 U6095 ( .A1(n4824), .A2(n4823), .ZN(n4828) );
  XNOR2_X1 U6096 ( .A(n4908), .B(n7571), .ZN(n4827) );
  XNOR2_X1 U6097 ( .A(n4907), .B(n7572), .ZN(n4826) );
  XNOR2_X1 U6098 ( .A(instr_addr_o_21_), .B(n7584), .ZN(n4825) );
  NAND4_X1 U6099 ( .A1(n4828), .A2(n4827), .A3(n4826), .A4(n4825), .ZN(n4829)
         );
  NOR3_X1 U6100 ( .A1(n4831), .A2(n4830), .A3(n4829), .ZN(n4832) );
  INV_X1 U6101 ( .A(n4833), .ZN(n4834) );
  NAND2_X1 U6102 ( .A1(n4834), .A2(n11533), .ZN(n4840) );
  XNOR2_X1 U6103 ( .A(n4802), .B(n10636), .ZN(n4839) );
  XNOR2_X1 U6104 ( .A(n4835), .B(n10628), .ZN(n4838) );
  XNOR2_X1 U6105 ( .A(n12213), .B(n10637), .ZN(n4837) );
  NAND4_X1 U6106 ( .A1(n4840), .A2(n4839), .A3(n4838), .A4(n4837), .ZN(n4856)
         );
  INV_X1 U6107 ( .A(n4841), .ZN(n4847) );
  NAND2_X1 U6108 ( .A1(n11530), .A2(pmp_addr_i[200]), .ZN(n11553) );
  NAND3_X1 U6109 ( .A1(instr_addr_o_11_), .A2(n10498), .A3(n11553), .ZN(n4846)
         );
  INV_X1 U6110 ( .A(n4842), .ZN(n11535) );
  NAND3_X1 U6111 ( .A1(instr_addr_o_6_), .A2(n10654), .A3(n11535), .ZN(n4845)
         );
  NAND3_X1 U6112 ( .A1(n5740), .A2(n4843), .A3(n11543), .ZN(n4844) );
  NAND4_X1 U6113 ( .A1(n4847), .A2(n4846), .A3(n4845), .A4(n4844), .ZN(n4855)
         );
  NAND3_X1 U6114 ( .A1(n154), .A2(n4848), .A3(n11526), .ZN(n4852) );
  NAND3_X1 U6115 ( .A1(instr_addr_o_15_), .A2(n10658), .A3(n11522), .ZN(n4851)
         );
  NAND3_X1 U6116 ( .A1(instr_addr_o_13_), .A2(n4849), .A3(n11570), .ZN(n4850)
         );
  NAND4_X1 U6117 ( .A1(n4853), .A2(n4852), .A3(n4851), .A4(n4850), .ZN(n4854)
         );
  NOR3_X1 U6118 ( .A1(n4856), .A2(n4855), .A3(n4854), .ZN(n4919) );
  XNOR2_X1 U6119 ( .A(n5062), .B(n4857), .ZN(n4858) );
  NAND2_X1 U6120 ( .A1(n4858), .A2(n11564), .ZN(n4864) );
  XNOR2_X1 U6121 ( .A(n6025), .B(n10639), .ZN(n4863) );
  INV_X1 U6122 ( .A(n4860), .ZN(n4862) );
  NAND4_X1 U6123 ( .A1(n4864), .A2(n4863), .A3(n4862), .A4(n4861), .ZN(n4878)
         );
  INV_X1 U6124 ( .A(n4865), .ZN(n4868) );
  XNOR2_X1 U6125 ( .A(n4866), .B(n10661), .ZN(n4867) );
  NAND3_X1 U6126 ( .A1(n4869), .A2(n4868), .A3(n4867), .ZN(n4877) );
  INV_X1 U6127 ( .A(n4870), .ZN(n4875) );
  INV_X1 U6128 ( .A(n4871), .ZN(n4874) );
  INV_X1 U6129 ( .A(n4872), .ZN(n4873) );
  NAND4_X1 U6130 ( .A1(n4875), .A2(n4874), .A3(n320), .A4(n4873), .ZN(n4876)
         );
  NOR3_X1 U6131 ( .A1(n4878), .A2(n4877), .A3(n4876), .ZN(n4918) );
  XNOR2_X1 U6132 ( .A(n5162), .B(n10615), .ZN(n4882) );
  NOR2_X1 U6133 ( .A1(n10506), .A2(n11521), .ZN(n4880) );
  NOR2_X1 U6134 ( .A1(n10502), .A2(n11530), .ZN(n4879) );
  AOI22_X1 U6135 ( .A1(instr_addr_o_12_), .A2(n4880), .B1(n5262), .B2(n4879), 
        .ZN(n4881) );
  NAND2_X1 U6136 ( .A1(n4882), .A2(n4881), .ZN(n4890) );
  NOR2_X1 U6137 ( .A1(n10519), .A2(n11561), .ZN(n4885) );
  INV_X1 U6138 ( .A(n4883), .ZN(n4884) );
  NOR2_X1 U6139 ( .A1(n11568), .A2(n4884), .ZN(n11567) );
  AOI22_X1 U6140 ( .A1(n12180), .A2(n4885), .B1(n12203), .B2(n11567), .ZN(
        n4888) );
  XNOR2_X1 U6141 ( .A(n137), .B(n10613), .ZN(n4887) );
  NAND3_X1 U6142 ( .A1(n4888), .A2(n4887), .A3(n4886), .ZN(n4889) );
  NAND3_X1 U6143 ( .A1(n12150), .A2(n10650), .A3(n651), .ZN(n4898) );
  INV_X1 U6144 ( .A(n4891), .ZN(n11545) );
  NOR2_X1 U6145 ( .A1(n10485), .A2(n11545), .ZN(n4896) );
  NAND2_X1 U6146 ( .A1(n4893), .A2(n4892), .ZN(n10670) );
  NAND4_X1 U6147 ( .A1(n10670), .A2(pmp_cfg_i[52]), .A3(n4894), .A4(
        pmp_cfg_i[50]), .ZN(n4895) );
  AOI21_X1 U6148 ( .B1(n6015), .B2(n4896), .A(n4895), .ZN(n4897) );
  OAI211_X1 U6149 ( .C1(n12150), .C2(n10650), .A(n4898), .B(n4897), .ZN(n4899)
         );
  INV_X1 U6150 ( .A(n4899), .ZN(n4905) );
  XNOR2_X1 U6151 ( .A(n4900), .B(n10648), .ZN(n4904) );
  XNOR2_X1 U6152 ( .A(n5980), .B(n10623), .ZN(n4903) );
  XNOR2_X1 U6153 ( .A(n4901), .B(n10634), .ZN(n4902) );
  NAND4_X1 U6154 ( .A1(n4905), .A2(n4904), .A3(n4903), .A4(n4902), .ZN(n4915)
         );
  XNOR2_X1 U6155 ( .A(instr_addr_o_21_), .B(n10611), .ZN(n4913) );
  XNOR2_X1 U6156 ( .A(n4907), .B(n10626), .ZN(n4912) );
  XNOR2_X1 U6157 ( .A(n4908), .B(n10625), .ZN(n4911) );
  XNOR2_X1 U6158 ( .A(n5985), .B(n10605), .ZN(n4910) );
  NAND4_X1 U6159 ( .A1(n4913), .A2(n4912), .A3(n4911), .A4(n4910), .ZN(n4914)
         );
  NOR2_X1 U6160 ( .A1(n4915), .A2(n4914), .ZN(n4916) );
  NAND4_X1 U6161 ( .A1(n4919), .A2(n4918), .A3(n4917), .A4(n4916), .ZN(n5016)
         );
  INV_X1 U6162 ( .A(n4920), .ZN(n4927) );
  INV_X1 U6163 ( .A(n4921), .ZN(n4926) );
  NOR2_X1 U6164 ( .A1(n8235), .A2(pmp_addr_i[39]), .ZN(n4922) );
  NAND2_X1 U6165 ( .A1(n5270), .A2(n4922), .ZN(n4924) );
  INV_X1 U6166 ( .A(n11479), .ZN(n4923) );
  NAND4_X1 U6167 ( .A1(n4924), .A2(pmp_addr_i[37]), .A3(pmp_addr_i[38]), .A4(
        n4923), .ZN(n4925) );
  OAI21_X1 U6168 ( .B1(n4927), .B2(n4926), .A(n4925), .ZN(n4931) );
  NOR2_X1 U6169 ( .A1(n4929), .A2(n4928), .ZN(n4930) );
  OAI211_X1 U6170 ( .C1(n11476), .C2(n4932), .A(n4931), .B(n4930), .ZN(n4947)
         );
  OR2_X1 U6171 ( .A1(n11512), .A2(n4933), .ZN(n11502) );
  NOR2_X1 U6172 ( .A1(n11502), .A2(n4934), .ZN(n11492) );
  XNOR2_X1 U6173 ( .A(n6025), .B(n8351), .ZN(n4935) );
  OAI21_X1 U6174 ( .B1(n4936), .B2(n11492), .A(n4935), .ZN(n4946) );
  OR2_X1 U6175 ( .A1(n11493), .A2(n4937), .ZN(n4938) );
  NOR2_X1 U6176 ( .A1(n11512), .A2(n4938), .ZN(n11508) );
  INV_X1 U6177 ( .A(n4939), .ZN(n4944) );
  INV_X1 U6178 ( .A(n4940), .ZN(n4943) );
  INV_X1 U6179 ( .A(n4941), .ZN(n4942) );
  OAI211_X1 U6180 ( .C1(n11508), .C2(n4944), .A(n4943), .B(n4942), .ZN(n4945)
         );
  NOR2_X1 U6181 ( .A1(n4949), .A2(n4948), .ZN(n4953) );
  XNOR2_X1 U6182 ( .A(instr_addr_o_21_), .B(n8367), .ZN(n4952) );
  XNOR2_X1 U6183 ( .A(n5985), .B(n8359), .ZN(n4951) );
  XNOR2_X1 U6184 ( .A(n6020), .B(n8348), .ZN(n4950) );
  NAND4_X1 U6185 ( .A1(n4953), .A2(n4952), .A3(n4951), .A4(n4950), .ZN(n4964)
         );
  INV_X1 U6186 ( .A(n11502), .ZN(n4954) );
  AOI21_X1 U6187 ( .B1(n4956), .B2(n4955), .A(n4954), .ZN(n4963) );
  INV_X1 U6188 ( .A(n4957), .ZN(n4961) );
  INV_X1 U6189 ( .A(n4958), .ZN(n4960) );
  XNOR2_X1 U6190 ( .A(instr_addr_o_31_), .B(n8276), .ZN(n4959) );
  NAND3_X1 U6191 ( .A1(n4961), .A2(n4960), .A3(n4959), .ZN(n4962) );
  NOR3_X1 U6192 ( .A1(n4964), .A2(n4963), .A3(n4962), .ZN(n5013) );
  NOR2_X1 U6193 ( .A1(n4966), .A2(n4965), .ZN(n4975) );
  INV_X1 U6194 ( .A(n4967), .ZN(n4968) );
  NOR2_X1 U6195 ( .A1(n8204), .A2(n4968), .ZN(n4969) );
  AND2_X1 U6196 ( .A1(n12179), .A2(n4969), .ZN(n4971) );
  NOR2_X1 U6197 ( .A1(n4971), .A2(n4970), .ZN(n4974) );
  XNOR2_X1 U6198 ( .A(n4802), .B(n8349), .ZN(n4973) );
  XNOR2_X1 U6199 ( .A(n6028), .B(n8368), .ZN(n4972) );
  NAND4_X1 U6200 ( .A1(n4975), .A2(n4974), .A3(n4973), .A4(n4972), .ZN(n4987)
         );
  INV_X1 U6201 ( .A(n4976), .ZN(n4978) );
  OAI211_X1 U6202 ( .C1(n11473), .C2(n4979), .A(n4978), .B(n4977), .ZN(n4986)
         );
  INV_X1 U6203 ( .A(n4980), .ZN(n4984) );
  INV_X1 U6204 ( .A(n11508), .ZN(n4982) );
  NOR2_X1 U6205 ( .A1(n4982), .A2(n4981), .ZN(n11465) );
  XNOR2_X1 U6206 ( .A(instr_addr_o_22_), .B(n8350), .ZN(n4983) );
  OAI21_X1 U6207 ( .B1(n4984), .B2(n11465), .A(n4983), .ZN(n4985) );
  INV_X1 U6208 ( .A(n11487), .ZN(n4992) );
  NAND3_X1 U6209 ( .A1(n205), .A2(n8339), .A3(n11512), .ZN(n4991) );
  NAND3_X1 U6210 ( .A1(n12267), .A2(n4989), .A3(n11479), .ZN(n4990) );
  OAI211_X1 U6211 ( .C1(n4993), .C2(n4992), .A(n4991), .B(n4990), .ZN(n4994)
         );
  INV_X1 U6212 ( .A(n4994), .ZN(n5007) );
  INV_X1 U6213 ( .A(n4995), .ZN(n11484) );
  NOR2_X1 U6214 ( .A1(n8219), .A2(n11484), .ZN(n4999) );
  NAND2_X1 U6215 ( .A1(n4996), .A2(n160), .ZN(n8391) );
  NAND4_X1 U6216 ( .A1(n8391), .A2(pmp_cfg_i[12]), .A3(n4997), .A4(
        pmp_cfg_i[10]), .ZN(n4998) );
  AOI21_X1 U6217 ( .B1(n5976), .B2(n4999), .A(n4998), .ZN(n5002) );
  OAI211_X1 U6218 ( .C1(n12150), .C2(n8334), .A(n5002), .B(n5001), .ZN(n5003)
         );
  INV_X1 U6219 ( .A(n5003), .ZN(n5006) );
  XNOR2_X1 U6220 ( .A(n137), .B(n8358), .ZN(n5005) );
  XNOR2_X1 U6221 ( .A(instr_addr_o_28_), .B(n8360), .ZN(n5004) );
  XNOR2_X1 U6222 ( .A(n4908), .B(n8366), .ZN(n5011) );
  XNOR2_X1 U6223 ( .A(n4556), .B(n8369), .ZN(n5010) );
  XNOR2_X1 U6224 ( .A(n5980), .B(n8361), .ZN(n5009) );
  XNOR2_X1 U6225 ( .A(n5550), .B(n8330), .ZN(n5008) );
  NAND4_X1 U6226 ( .A1(n5011), .A2(n5010), .A3(n5009), .A4(n5008), .ZN(n5012)
         );
  AND4_X1 U6227 ( .A1(n5017), .A2(n5018), .A3(n5016), .A4(n5015), .ZN(n5019)
         );
  NAND4_X1 U6228 ( .A1(n5022), .A2(n5021), .A3(n5020), .A4(n5019), .ZN(n12133)
         );
  NOR2_X1 U6229 ( .A1(n5280), .A2(n5859), .ZN(n5024) );
  OR2_X1 U6230 ( .A1(pmp_addr_i[161]), .A2(pmp_addr_i[160]), .ZN(n5025) );
  NOR2_X1 U6231 ( .A1(n5025), .A2(pmp_addr_i[162]), .ZN(n5028) );
  INV_X1 U6232 ( .A(n5025), .ZN(n5027) );
  INV_X1 U6233 ( .A(pmp_addr_i[162]), .ZN(n5026) );
  OAI22_X1 U6234 ( .A1(n5899), .A2(n5028), .B1(n5027), .B2(n5026), .ZN(n5029)
         );
  OAI211_X1 U6235 ( .C1(pmp_addr_i[163]), .C2(n3839), .A(n5030), .B(n5029), 
        .ZN(n5034) );
  INV_X1 U6237 ( .A(pmp_addr_i[166]), .ZN(n5036) );
  NAND2_X1 U6238 ( .A1(n5269), .A2(n5036), .ZN(n5037) );
  NAND2_X1 U6239 ( .A1(n5262), .A2(n5867), .ZN(n5042) );
  NAND2_X1 U6240 ( .A1(n5740), .A2(n5866), .ZN(n5032) );
  NAND4_X1 U6241 ( .A1(n5038), .A2(n5037), .A3(n5042), .A4(n5032), .ZN(n5033)
         );
  AOI21_X1 U6242 ( .B1(n5035), .B2(n5034), .A(n5033), .ZN(n5055) );
  OAI22_X1 U6243 ( .A1(n5740), .A2(n5866), .B1(n205), .B2(n5036), .ZN(n5039)
         );
  NAND4_X1 U6244 ( .A1(n5039), .A2(n5038), .A3(n5042), .A4(n5037), .ZN(n5045)
         );
  NOR2_X1 U6245 ( .A1(n5040), .A2(n5258), .ZN(n5043) );
  AOI22_X1 U6246 ( .A1(n5043), .A2(n5042), .B1(n4602), .B2(pmp_addr_i[168]), 
        .ZN(n5044) );
  INV_X1 U6247 ( .A(pmp_addr_i[176]), .ZN(n5046) );
  NAND2_X1 U6248 ( .A1(gte_x_382_A_16_), .A2(n5046), .ZN(n5064) );
  OAI21_X1 U6249 ( .B1(n5048), .B2(pmp_addr_i[175]), .A(n5064), .ZN(n5066) );
  INV_X1 U6250 ( .A(pmp_addr_i[174]), .ZN(n5049) );
  NAND2_X1 U6251 ( .A1(n12266), .A2(n5049), .ZN(n5060) );
  OAI21_X1 U6252 ( .B1(n6017), .B2(pmp_addr_i[173]), .A(n5060), .ZN(n5050) );
  NOR2_X1 U6253 ( .A1(n5066), .A2(n5050), .ZN(n5079) );
  NAND2_X1 U6254 ( .A1(n4788), .A2(n5235), .ZN(n5074) );
  NAND2_X1 U6255 ( .A1(instr_addr_o_13_), .A2(n5239), .ZN(n5051) );
  NAND2_X1 U6256 ( .A1(n5074), .A2(n5051), .ZN(n5076) );
  NAND2_X1 U6257 ( .A1(n5245), .A2(n5243), .ZN(n5072) );
  OAI21_X1 U6258 ( .B1(n5052), .B2(pmp_addr_i[169]), .A(n5072), .ZN(n5053) );
  NOR2_X1 U6259 ( .A1(n5076), .A2(n5053), .ZN(n5054) );
  INV_X1 U6260 ( .A(pmp_addr_i[173]), .ZN(n5056) );
  NOR2_X1 U6261 ( .A1(n4498), .A2(n5056), .ZN(n5059) );
  AOI22_X1 U6262 ( .A1(n5060), .A2(n5059), .B1(n5058), .B2(pmp_addr_i[174]), 
        .ZN(n5067) );
  INV_X1 U6263 ( .A(pmp_addr_i[175]), .ZN(n5061) );
  NOR2_X1 U6264 ( .A1(n5062), .A2(n5061), .ZN(n5063) );
  AOI22_X1 U6265 ( .A1(n5064), .A2(n5063), .B1(n2082), .B2(pmp_addr_i[176]), 
        .ZN(n5065) );
  OAI21_X1 U6266 ( .B1(n5067), .B2(n5066), .A(n5065), .ZN(n5068) );
  INV_X1 U6267 ( .A(n5068), .ZN(n5081) );
  NOR2_X1 U6268 ( .A1(n3934), .A2(n5868), .ZN(n5071) );
  AOI22_X1 U6269 ( .A1(n5072), .A2(n5071), .B1(n5070), .B2(pmp_addr_i[170]), 
        .ZN(n5077) );
  NOR2_X1 U6270 ( .A1(n5997), .A2(n5239), .ZN(n5073) );
  AOI22_X1 U6271 ( .A1(n5074), .A2(n5073), .B1(instr_addr_o_14__BAR), .B2(
        pmp_addr_i[172]), .ZN(n5075) );
  OAI21_X1 U6272 ( .B1(n5077), .B2(n5076), .A(n5075), .ZN(n5078) );
  NAND2_X1 U6273 ( .A1(n5078), .A2(n5079), .ZN(n5080) );
  INV_X1 U6274 ( .A(pmp_addr_i[184]), .ZN(n5083) );
  NAND2_X1 U6275 ( .A1(n210), .A2(n5083), .ZN(n5131) );
  INV_X1 U6276 ( .A(pmp_addr_i[183]), .ZN(n5129) );
  NAND2_X1 U6277 ( .A1(n136), .A2(n5129), .ZN(n5084) );
  AND2_X1 U6278 ( .A1(n5131), .A2(n5084), .ZN(n5125) );
  INV_X1 U6279 ( .A(pmp_addr_i[182]), .ZN(n5085) );
  NAND2_X1 U6280 ( .A1(n6028), .A2(n5085), .ZN(n5128) );
  OAI211_X1 U6281 ( .C1(pmp_addr_i[181]), .C2(n5086), .A(n5125), .B(n5128), 
        .ZN(n5097) );
  INV_X1 U6282 ( .A(pmp_addr_i[180]), .ZN(n5087) );
  NAND2_X1 U6283 ( .A1(n12157), .A2(n5087), .ZN(n5105) );
  INV_X1 U6284 ( .A(pmp_addr_i[179]), .ZN(n5104) );
  NAND2_X1 U6285 ( .A1(n5191), .A2(n5104), .ZN(n5088) );
  AND2_X1 U6286 ( .A1(n5105), .A2(n5088), .ZN(n5103) );
  INV_X1 U6287 ( .A(pmp_addr_i[178]), .ZN(n5089) );
  NAND2_X1 U6288 ( .A1(instr_addr_o_20_), .A2(n5089), .ZN(n5101) );
  OAI211_X1 U6289 ( .C1(pmp_addr_i[177]), .C2(n12208), .A(n5103), .B(n5101), 
        .ZN(n5091) );
  NOR2_X1 U6290 ( .A1(n5097), .A2(n5091), .ZN(n5096) );
  INV_X1 U6291 ( .A(pmp_addr_i[188]), .ZN(n5092) );
  NAND2_X1 U6292 ( .A1(n12161), .A2(n5092), .ZN(n5117) );
  OAI21_X1 U6293 ( .B1(n4656), .B2(pmp_addr_i[187]), .A(n5117), .ZN(n5119) );
  INV_X1 U6294 ( .A(pmp_addr_i[186]), .ZN(n5093) );
  NAND2_X1 U6295 ( .A1(n6018), .A2(n12073), .ZN(n5122) );
  NOR2_X1 U6296 ( .A1(n5119), .A2(n5095), .ZN(n5139) );
  INV_X1 U6297 ( .A(n5097), .ZN(n5098) );
  INV_X1 U6298 ( .A(pmp_addr_i[177]), .ZN(n5099) );
  NOR2_X1 U6299 ( .A1(n5100), .A2(n5099), .ZN(n5102) );
  AOI22_X1 U6300 ( .A1(n5102), .A2(n5101), .B1(n4631), .B2(pmp_addr_i[178]), 
        .ZN(n5109) );
  INV_X1 U6301 ( .A(n5103), .ZN(n5108) );
  NOR2_X1 U6302 ( .A1(instr_addr_o_21_), .A2(n5104), .ZN(n5106) );
  AOI22_X1 U6303 ( .A1(n5106), .A2(n5105), .B1(n999), .B2(pmp_addr_i[180]), 
        .ZN(n5107) );
  OAI21_X1 U6304 ( .B1(n5109), .B2(n5108), .A(n5107), .ZN(n5123) );
  INV_X1 U6305 ( .A(pmp_addr_i[185]), .ZN(n5110) );
  NOR2_X1 U6306 ( .A1(n5162), .A2(n5110), .ZN(n5112) );
  AOI22_X1 U6307 ( .A1(n5113), .A2(n5112), .B1(n5111), .B2(pmp_addr_i[186]), 
        .ZN(n5120) );
  INV_X1 U6308 ( .A(pmp_addr_i[187]), .ZN(n5114) );
  NOR2_X1 U6309 ( .A1(n5149), .A2(n5114), .ZN(n5116) );
  AOI22_X1 U6310 ( .A1(n5117), .A2(n5116), .B1(n5115), .B2(pmp_addr_i[188]), 
        .ZN(n5118) );
  OAI21_X1 U6311 ( .B1(n5120), .B2(n5119), .A(n5118), .ZN(n5121) );
  AOI22_X1 U6312 ( .A1(n5124), .A2(n5123), .B1(n5122), .B2(n5121), .ZN(n5141)
         );
  INV_X1 U6313 ( .A(n5125), .ZN(n5134) );
  INV_X1 U6314 ( .A(pmp_addr_i[181]), .ZN(n5126) );
  NOR2_X1 U6315 ( .A1(n5208), .A2(n5126), .ZN(n5127) );
  AOI22_X1 U6316 ( .A1(n5128), .A2(n5127), .B1(n2580), .B2(pmp_addr_i[182]), 
        .ZN(n5133) );
  NOR2_X1 U6317 ( .A1(n12226), .A2(n5129), .ZN(n5130) );
  AOI22_X1 U6318 ( .A1(n5131), .A2(n5130), .B1(n1273), .B2(pmp_addr_i[184]), 
        .ZN(n5132) );
  OAI21_X1 U6319 ( .B1(n5134), .B2(n5133), .A(n5132), .ZN(n5138) );
  OAI21_X1 U6320 ( .B1(n5136), .B2(n12073), .A(n5135), .ZN(n5137) );
  INV_X1 U6321 ( .A(pmp_addr_i[155]), .ZN(n5148) );
  INV_X1 U6322 ( .A(pmp_cfg_i[43]), .ZN(n5283) );
  INV_X1 U6323 ( .A(n161), .ZN(n5276) );
  INV_X1 U6324 ( .A(pmp_cfg_i[44]), .ZN(n5255) );
  NAND4_X1 U6325 ( .A1(pmp_addr_i[166]), .A2(pmp_addr_i[165]), .A3(
        pmp_addr_i[168]), .A4(pmp_addr_i[167]), .ZN(n5144) );
  NAND2_X1 U6326 ( .A1(pmp_addr_i[170]), .A2(pmp_addr_i[169]), .ZN(n5143) );
  NOR2_X1 U6327 ( .A1(n5144), .A2(n5143), .ZN(n5237) );
  AND2_X1 U6328 ( .A1(pmp_addr_i[171]), .A2(pmp_addr_i[172]), .ZN(n5861) );
  NAND2_X1 U6329 ( .A1(n5237), .A2(n5861), .ZN(n5227) );
  NAND2_X1 U6330 ( .A1(pmp_addr_i[164]), .A2(pmp_addr_i[163]), .ZN(n5222) );
  NOR2_X1 U6331 ( .A1(n5222), .A2(n5056), .ZN(n5145) );
  AND3_X1 U6332 ( .A1(pmp_addr_i[160]), .A2(pmp_addr_i[161]), .A3(
        pmp_addr_i[162]), .ZN(n5857) );
  NAND4_X1 U6333 ( .A1(n5145), .A2(n5857), .A3(pmp_addr_i[174]), .A4(
        pmp_addr_i[175]), .ZN(n5146) );
  AND2_X1 U6334 ( .A1(pmp_cfg_i[43]), .A2(pmp_cfg_i[44]), .ZN(n5880) );
  OAI21_X1 U6335 ( .B1(n5227), .B2(n5146), .A(n5880), .ZN(n11381) );
  OAI21_X1 U6336 ( .B1(pmp_cfg_i[43]), .B2(n5255), .A(n11381), .ZN(n5914) );
  NAND2_X1 U6337 ( .A1(n215), .A2(pmp_addr_i[187]), .ZN(n5147) );
  OAI21_X1 U6338 ( .B1(n5148), .B2(n5276), .A(n5147), .ZN(n11012) );
  INV_X1 U6339 ( .A(n11012), .ZN(n5155) );
  AND2_X1 U6340 ( .A1(n5149), .A2(n5155), .ZN(n5153) );
  NAND2_X1 U6341 ( .A1(n5914), .A2(pmp_addr_i[188]), .ZN(n5150) );
  OAI21_X1 U6342 ( .B1(n5276), .B2(n1349), .A(n5150), .ZN(n10974) );
  INV_X1 U6343 ( .A(n10974), .ZN(n5151) );
  NOR2_X1 U6344 ( .A1(n12263), .A2(n5151), .ZN(n5157) );
  INV_X1 U6345 ( .A(n5157), .ZN(n5152) );
  AOI22_X1 U6346 ( .A1(n5153), .A2(n5152), .B1(n12199), .B2(n5151), .ZN(n5170)
         );
  NAND2_X1 U6347 ( .A1(n215), .A2(pmp_addr_i[189]), .ZN(n11461) );
  OAI21_X1 U6348 ( .B1(n5276), .B2(n1373), .A(n11461), .ZN(n11007) );
  INV_X1 U6349 ( .A(n11007), .ZN(n5166) );
  OAI21_X1 U6350 ( .B1(n5154), .B2(n5166), .A(n9451), .ZN(n5169) );
  NOR2_X1 U6351 ( .A1(instr_addr_o_29_), .A2(n5155), .ZN(n5156) );
  NOR2_X1 U6352 ( .A1(n5157), .A2(n5156), .ZN(n5175) );
  INV_X1 U6353 ( .A(n5169), .ZN(n5174) );
  NAND2_X1 U6354 ( .A1(n5914), .A2(pmp_addr_i[186]), .ZN(n5158) );
  OAI21_X1 U6355 ( .B1(n1350), .B2(n5276), .A(n5158), .ZN(n10973) );
  INV_X1 U6356 ( .A(n10973), .ZN(n5159) );
  NOR2_X1 U6357 ( .A1(n5368), .A2(n5159), .ZN(n5171) );
  NAND2_X1 U6358 ( .A1(n215), .A2(pmp_addr_i[185]), .ZN(n5160) );
  OAI21_X1 U6359 ( .B1(n1389), .B2(n5276), .A(n5160), .ZN(n10990) );
  INV_X1 U6360 ( .A(n10990), .ZN(n5161) );
  NAND2_X1 U6361 ( .A1(n5162), .A2(n5161), .ZN(n5164) );
  OAI22_X1 U6362 ( .A1(n5171), .A2(n5164), .B1(n5163), .B2(n10973), .ZN(n5165)
         );
  NAND3_X1 U6363 ( .A1(n5175), .A2(n5174), .A3(n5165), .ZN(n5168) );
  NAND3_X1 U6364 ( .A1(n147), .A2(n5166), .A3(n9451), .ZN(n5167) );
  OAI211_X1 U6365 ( .C1(n5170), .C2(n5169), .A(n5168), .B(n5167), .ZN(n5321)
         );
  INV_X1 U6366 ( .A(n5321), .ZN(n5178) );
  INV_X1 U6367 ( .A(n5171), .ZN(n5173) );
  NAND2_X1 U6368 ( .A1(n4147), .A2(n10990), .ZN(n5172) );
  NAND4_X1 U6369 ( .A1(n5175), .A2(n5174), .A3(n5173), .A4(n5172), .ZN(n5177)
         );
  NAND2_X1 U6370 ( .A1(n161), .A2(pmp_cfg_i[42]), .ZN(n5176) );
  AOI21_X1 U6371 ( .B1(n5178), .B2(n5177), .A(n5176), .ZN(n5323) );
  NAND2_X1 U6372 ( .A1(n215), .A2(pmp_addr_i[180]), .ZN(n5179) );
  OAI21_X1 U6373 ( .B1(n5276), .B2(n1355), .A(n5179), .ZN(n10981) );
  INV_X1 U6374 ( .A(n10981), .ZN(n5180) );
  NOR2_X1 U6375 ( .A1(n5181), .A2(n5180), .ZN(n5194) );
  NAND2_X1 U6376 ( .A1(n215), .A2(pmp_addr_i[179]), .ZN(n5182) );
  OAI21_X1 U6377 ( .B1(n1383), .B2(n5276), .A(n5182), .ZN(n10980) );
  INV_X1 U6378 ( .A(n10980), .ZN(n5190) );
  NOR2_X1 U6379 ( .A1(n5183), .A2(n5190), .ZN(n5184) );
  NOR2_X1 U6380 ( .A1(n5194), .A2(n5184), .ZN(n5316) );
  NAND2_X1 U6381 ( .A1(n215), .A2(pmp_addr_i[178]), .ZN(n5185) );
  OAI21_X1 U6382 ( .B1(n1357), .B2(n5276), .A(n5185), .ZN(n10979) );
  INV_X1 U6383 ( .A(n10979), .ZN(n5186) );
  NOR2_X1 U6384 ( .A1(n5187), .A2(n5186), .ZN(n5312) );
  NAND2_X1 U6385 ( .A1(n215), .A2(pmp_addr_i[177]), .ZN(n5188) );
  OAI21_X1 U6386 ( .B1(n5276), .B2(n1380), .A(n5188), .ZN(n10968) );
  NAND2_X1 U6387 ( .A1(n3793), .A2(n10885), .ZN(n5189) );
  OAI22_X1 U6388 ( .A1(n5312), .A2(n5189), .B1(n4631), .B2(n10979), .ZN(n5196)
         );
  NAND2_X1 U6389 ( .A1(n5191), .A2(n5190), .ZN(n5193) );
  OAI22_X1 U6390 ( .A1(n5194), .A2(n5193), .B1(n5192), .B2(n10981), .ZN(n5195)
         );
  AOI21_X1 U6391 ( .B1(n5316), .B2(n5196), .A(n5195), .ZN(n5218) );
  NAND2_X1 U6392 ( .A1(n215), .A2(pmp_addr_i[181]), .ZN(n5197) );
  OAI21_X1 U6393 ( .B1(n1364), .B2(n5276), .A(n5197), .ZN(n10982) );
  INV_X1 U6394 ( .A(n10982), .ZN(n5207) );
  NAND2_X1 U6395 ( .A1(n5914), .A2(pmp_addr_i[184]), .ZN(n5198) );
  OAI21_X1 U6396 ( .B1(n1351), .B2(n5276), .A(n5198), .ZN(n10989) );
  INV_X1 U6397 ( .A(n10989), .ZN(n5199) );
  NOR2_X1 U6398 ( .A1(n12158), .A2(n5199), .ZN(n5213) );
  NAND2_X1 U6399 ( .A1(n215), .A2(pmp_addr_i[183]), .ZN(n5201) );
  OAI21_X1 U6400 ( .B1(n1367), .B2(n5276), .A(n5201), .ZN(n10988) );
  INV_X1 U6401 ( .A(n10988), .ZN(n5211) );
  NOR2_X1 U6402 ( .A1(n4644), .A2(n5211), .ZN(n5203) );
  NOR2_X1 U6403 ( .A1(n5213), .A2(n5203), .ZN(n5216) );
  NAND2_X1 U6404 ( .A1(n215), .A2(pmp_addr_i[182]), .ZN(n5204) );
  OAI21_X1 U6405 ( .B1(n1353), .B2(n5276), .A(n5204), .ZN(n10987) );
  INV_X1 U6406 ( .A(n10987), .ZN(n5205) );
  NOR2_X1 U6407 ( .A1(n5330), .A2(n5205), .ZN(n5210) );
  INV_X1 U6408 ( .A(n5210), .ZN(n5206) );
  NAND2_X1 U6410 ( .A1(n5208), .A2(n5207), .ZN(n5209) );
  OAI22_X1 U6411 ( .A1(n5210), .A2(n5209), .B1(n1269), .B2(n10987), .ZN(n5215)
         );
  NAND2_X1 U6412 ( .A1(n136), .A2(n5211), .ZN(n5212) );
  OAI22_X1 U6413 ( .A1(n5213), .A2(n5212), .B1(n1273), .B2(n10989), .ZN(n5214)
         );
  AOI21_X1 U6414 ( .B1(n5216), .B2(n5215), .A(n5214), .ZN(n5217) );
  OAI21_X1 U6415 ( .B1(n5218), .B2(n5318), .A(n5217), .ZN(n5320) );
  NOR2_X1 U6416 ( .A1(n5320), .A2(n5321), .ZN(n5311) );
  NAND2_X1 U6417 ( .A1(n5914), .A2(pmp_addr_i[176]), .ZN(n5219) );
  OAI21_X1 U6418 ( .B1(n1327), .B2(n5276), .A(n5219), .ZN(n10966) );
  INV_X1 U6419 ( .A(n10966), .ZN(n5220) );
  NOR2_X1 U6420 ( .A1(n6019), .A2(n5220), .ZN(n5231) );
  NAND2_X1 U6421 ( .A1(n215), .A2(pmp_addr_i[175]), .ZN(n5221) );
  OAI21_X1 U6422 ( .B1(n5276), .B2(n1339), .A(n5221), .ZN(n10965) );
  NOR2_X1 U6423 ( .A1(n12156), .A2(n10856), .ZN(n5849) );
  NOR2_X1 U6424 ( .A1(n5231), .A2(n5849), .ZN(n5305) );
  OR2_X1 U6425 ( .A1(n5227), .A2(n5056), .ZN(n5223) );
  NAND2_X1 U6426 ( .A1(n5857), .A2(pmp_cfg_i[43]), .ZN(n5278) );
  OR2_X1 U6427 ( .A1(n5278), .A2(n5222), .ZN(n5274) );
  OAI211_X1 U6428 ( .C1(n5223), .C2(n5274), .A(pmp_cfg_i[44]), .B(
        pmp_addr_i[174]), .ZN(n5224) );
  OAI21_X1 U6429 ( .B1(n5225), .B2(n5276), .A(n5224), .ZN(n10802) );
  INV_X1 U6430 ( .A(n10802), .ZN(n11015) );
  OR2_X1 U6431 ( .A1(n3100), .A2(n11015), .ZN(n5303) );
  INV_X1 U6432 ( .A(n5303), .ZN(n5839) );
  OAI21_X1 U6433 ( .B1(n5274), .B2(n5227), .A(pmp_cfg_i[44]), .ZN(n5236) );
  NAND2_X1 U6434 ( .A1(n161), .A2(pmp_addr_i[141]), .ZN(n5228) );
  OAI21_X1 U6435 ( .B1(n5236), .B2(n5056), .A(n5228), .ZN(n10803) );
  INV_X1 U6436 ( .A(n10803), .ZN(n10948) );
  NAND2_X1 U6437 ( .A1(n208), .A2(n10948), .ZN(n5904) );
  NAND2_X1 U6438 ( .A1(n5229), .A2(n11015), .ZN(n5894) );
  OAI21_X1 U6439 ( .B1(n5839), .B2(n5904), .A(n5894), .ZN(n5233) );
  NAND2_X1 U6440 ( .A1(n5974), .A2(n10856), .ZN(n5902) );
  OAI22_X1 U6441 ( .A1(n5231), .A2(n5902), .B1(instr_addr_o_18__BAR), .B2(
        n10966), .ZN(n5232) );
  AOI21_X1 U6442 ( .B1(n5305), .B2(n5233), .A(n5232), .ZN(n5310) );
  NAND2_X1 U6443 ( .A1(n161), .A2(pmp_addr_i[140]), .ZN(n5234) );
  OAI21_X1 U6444 ( .B1(n5236), .B2(n5235), .A(n5234), .ZN(n10809) );
  INV_X1 U6445 ( .A(n10809), .ZN(n10945) );
  NOR2_X1 U6446 ( .A1(n12181), .A2(n10945), .ZN(n5252) );
  INV_X1 U6447 ( .A(n5237), .ZN(n5860) );
  OAI21_X1 U6448 ( .B1(n5274), .B2(n5860), .A(pmp_cfg_i[44]), .ZN(n5244) );
  NAND2_X1 U6449 ( .A1(n161), .A2(pmp_addr_i[139]), .ZN(n5238) );
  OAI21_X1 U6450 ( .B1(n5244), .B2(n5239), .A(n5238), .ZN(n11005) );
  INV_X1 U6451 ( .A(n11005), .ZN(n10947) );
  NAND2_X1 U6452 ( .A1(n149), .A2(n10947), .ZN(n5891) );
  NOR2_X1 U6453 ( .A1(n150), .A2(n10947), .ZN(n5241) );
  NOR2_X1 U6454 ( .A1(n5252), .A2(n5241), .ZN(n5833) );
  NAND2_X1 U6455 ( .A1(n161), .A2(pmp_addr_i[138]), .ZN(n5242) );
  OAI21_X1 U6456 ( .B1(n5244), .B2(n5243), .A(n5242), .ZN(n10807) );
  INV_X1 U6457 ( .A(n10807), .ZN(n10939) );
  OR2_X1 U6458 ( .A1(n5245), .A2(n10939), .ZN(n5302) );
  NAND2_X1 U6459 ( .A1(pmp_addr_i[166]), .A2(pmp_addr_i[165]), .ZN(n5246) );
  NOR2_X1 U6460 ( .A1(n5274), .A2(n5246), .ZN(n5256) );
  AND2_X1 U6461 ( .A1(pmp_addr_i[168]), .A2(pmp_addr_i[167]), .ZN(n5247) );
  AOI21_X1 U6462 ( .B1(n5256), .B2(n5247), .A(n5255), .ZN(n5259) );
  NAND2_X1 U6463 ( .A1(n5259), .A2(pmp_addr_i[169]), .ZN(n5248) );
  OAI21_X1 U6464 ( .B1(n5276), .B2(n5249), .A(n5248), .ZN(n10806) );
  INV_X1 U6465 ( .A(n10806), .ZN(n10946) );
  NAND2_X1 U6466 ( .A1(n5250), .A2(n10939), .ZN(n5903) );
  NAND2_X1 U6467 ( .A1(n5251), .A2(n10945), .ZN(n5893) );
  OR2_X1 U6468 ( .A1(n12179), .A2(n10948), .ZN(n5919) );
  NAND4_X1 U6469 ( .A1(n5254), .A2(n5305), .A3(n5303), .A4(n5919), .ZN(n5309)
         );
  OR2_X1 U6470 ( .A1(n5256), .A2(n5255), .ZN(n5265) );
  NAND2_X1 U6471 ( .A1(n161), .A2(pmp_addr_i[135]), .ZN(n5257) );
  OAI21_X1 U6472 ( .B1(n5265), .B2(n5258), .A(n5257), .ZN(n10832) );
  INV_X1 U6473 ( .A(n10832), .ZN(n10940) );
  OR2_X1 U6474 ( .A1(n155), .A2(n10940), .ZN(n5296) );
  INV_X1 U6475 ( .A(n5296), .ZN(n5263) );
  NAND2_X1 U6476 ( .A1(n5259), .A2(pmp_addr_i[168]), .ZN(n5260) );
  OAI21_X1 U6477 ( .B1(n5276), .B2(n5261), .A(n5260), .ZN(n10833) );
  INV_X1 U6478 ( .A(n10833), .ZN(n10942) );
  OR2_X1 U6479 ( .A1(n5270), .A2(n10942), .ZN(n5294) );
  INV_X1 U6480 ( .A(n5294), .ZN(n5271) );
  NOR2_X1 U6481 ( .A1(n5263), .A2(n5271), .ZN(n5834) );
  NAND2_X1 U6482 ( .A1(n161), .A2(pmp_addr_i[134]), .ZN(n5264) );
  OAI21_X1 U6483 ( .B1(n5265), .B2(n5036), .A(n5264), .ZN(n10829) );
  INV_X1 U6484 ( .A(n10829), .ZN(n10941) );
  OR2_X1 U6485 ( .A1(n5342), .A2(n10941), .ZN(n5295) );
  NAND3_X1 U6486 ( .A1(n5274), .A2(pmp_cfg_i[44]), .A3(pmp_addr_i[165]), .ZN(
        n5266) );
  OAI21_X1 U6487 ( .B1(n5276), .B2(n5267), .A(n5266), .ZN(n10830) );
  INV_X1 U6488 ( .A(n10830), .ZN(n10954) );
  NAND2_X1 U6489 ( .A1(n5269), .A2(n10941), .ZN(n5895) );
  NAND2_X1 U6490 ( .A1(n154), .A2(n10940), .ZN(n5892) );
  NAND2_X1 U6491 ( .A1(n5270), .A2(n10942), .ZN(n5901) );
  OAI21_X1 U6492 ( .B1(n5892), .B2(n5271), .A(n5901), .ZN(n5272) );
  AOI21_X1 U6493 ( .B1(n5834), .B2(n5273), .A(n5272), .ZN(n5301) );
  NAND3_X1 U6494 ( .A1(n5274), .A2(pmp_cfg_i[44]), .A3(pmp_addr_i[164]), .ZN(
        n5275) );
  OAI21_X1 U6495 ( .B1(n5276), .B2(n1308), .A(n5275), .ZN(n10814) );
  INV_X1 U6496 ( .A(n10814), .ZN(n10952) );
  NAND2_X1 U6497 ( .A1(n5278), .A2(pmp_cfg_i[44]), .ZN(n5282) );
  NAND2_X1 U6498 ( .A1(n161), .A2(pmp_addr_i[131]), .ZN(n5279) );
  OAI21_X1 U6499 ( .B1(n5282), .B2(n5859), .A(n5279), .ZN(n10813) );
  INV_X1 U6500 ( .A(n10813), .ZN(n10963) );
  NOR2_X1 U6501 ( .A1(n5280), .A2(n10963), .ZN(n5848) );
  NAND2_X1 U6502 ( .A1(n161), .A2(pmp_addr_i[130]), .ZN(n5281) );
  OAI21_X1 U6503 ( .B1(n5282), .B2(n5026), .A(n5281), .ZN(n10960) );
  NAND2_X1 U6504 ( .A1(n161), .A2(pmp_addr_i[128]), .ZN(n5285) );
  NAND2_X1 U6505 ( .A1(n5283), .A2(pmp_addr_i[160]), .ZN(n5284) );
  NAND2_X1 U6506 ( .A1(n5285), .A2(n5284), .ZN(n10957) );
  AND2_X1 U6507 ( .A1(pmp_cfg_i[43]), .A2(pmp_addr_i[160]), .ZN(n5288) );
  NAND2_X1 U6508 ( .A1(pmp_cfg_i[44]), .A2(pmp_addr_i[161]), .ZN(n5287) );
  NAND2_X1 U6509 ( .A1(n161), .A2(pmp_addr_i[129]), .ZN(n5286) );
  OAI21_X1 U6510 ( .B1(n5288), .B2(n5287), .A(n5286), .ZN(n10956) );
  OR2_X1 U6511 ( .A1(n10957), .A2(n10956), .ZN(n5289) );
  NAND2_X1 U6512 ( .A1(n10960), .A2(n5289), .ZN(n5290) );
  INV_X1 U6513 ( .A(n10960), .ZN(n5898) );
  INV_X1 U6514 ( .A(n5289), .ZN(n5915) );
  AOI22_X1 U6515 ( .A1(n3836), .A2(n5290), .B1(n5898), .B2(n5915), .ZN(n5292)
         );
  NOR3_X1 U6516 ( .A1(n5837), .A2(n5848), .A3(n5292), .ZN(n5299) );
  NAND2_X1 U6517 ( .A1(n5293), .A2(n10963), .ZN(n5900) );
  NAND2_X1 U6518 ( .A1(instr_addr_o_6_), .A2(n10952), .ZN(n5890) );
  OAI21_X1 U6519 ( .B1(n5837), .B2(n5900), .A(n5890), .ZN(n5298) );
  OR2_X1 U6520 ( .A1(n12267), .A2(n10954), .ZN(n5835) );
  AND4_X1 U6521 ( .A1(n5296), .A2(n5835), .A3(n5295), .A4(n5294), .ZN(n5297)
         );
  OAI21_X1 U6522 ( .B1(n5299), .B2(n5298), .A(n5297), .ZN(n5300) );
  OR2_X1 U6523 ( .A1(n6002), .A2(n10946), .ZN(n5838) );
  AND4_X1 U6524 ( .A1(n5919), .A2(n5838), .A3(n5303), .A4(n5302), .ZN(n5304)
         );
  NAND2_X1 U6525 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  INV_X1 U6526 ( .A(n5312), .ZN(n5315) );
  NAND2_X1 U6527 ( .A1(n5313), .A2(n10968), .ZN(n5314) );
  NAND3_X1 U6528 ( .A1(n5316), .A2(n5315), .A3(n5314), .ZN(n5317) );
  NOR2_X1 U6529 ( .A1(n5318), .A2(n5317), .ZN(n5319) );
  OR3_X1 U6530 ( .A1(n5320), .A2(n5321), .A3(n5319), .ZN(n5322) );
  NAND2_X1 U6531 ( .A1(n11037), .A2(pmp_addr_i[226]), .ZN(n5325) );
  NOR2_X1 U6532 ( .A1(n5326), .A2(n5325), .ZN(n5352) );
  OAI22_X1 U6533 ( .A1(n11068), .A2(n5328), .B1(n5327), .B2(n5352), .ZN(n5335)
         );
  INV_X1 U6534 ( .A(n5329), .ZN(n5333) );
  XNOR2_X1 U6535 ( .A(n5330), .B(n7250), .ZN(n5332) );
  NAND3_X1 U6536 ( .A1(instr_addr_o_9_), .A2(n7275), .A3(n11062), .ZN(n5331)
         );
  INV_X1 U6537 ( .A(n5336), .ZN(n5345) );
  OR2_X1 U6538 ( .A1(n5337), .A2(n7246), .ZN(n7317) );
  NAND3_X1 U6539 ( .A1(n7317), .A2(pmp_cfg_i[58]), .A3(n5338), .ZN(n5339) );
  AOI21_X1 U6540 ( .B1(n3876), .B2(n7142), .A(n5339), .ZN(n5344) );
  NOR2_X1 U6541 ( .A1(n7151), .A2(pmp_addr_i[229]), .ZN(n5341) );
  NOR2_X1 U6542 ( .A1(n7142), .A2(n11037), .ZN(n5340) );
  AOI22_X1 U6543 ( .A1(n5342), .A2(n5341), .B1(n5899), .B2(n5340), .ZN(n5343)
         );
  INV_X1 U6544 ( .A(n5346), .ZN(n5349) );
  XNOR2_X1 U6545 ( .A(n4802), .B(n5347), .ZN(n5348) );
  AOI21_X1 U6546 ( .B1(n5349), .B2(n11050), .A(n5348), .ZN(n5361) );
  NAND3_X1 U6547 ( .A1(n5351), .A2(n5350), .A3(pmp_cfg_i[60]), .ZN(n5354) );
  INV_X1 U6548 ( .A(n5352), .ZN(n11040) );
  NOR2_X1 U6549 ( .A1(n11040), .A2(n5353), .ZN(n11057) );
  NAND2_X1 U6550 ( .A1(n11057), .A2(pmp_addr_i[228]), .ZN(n11031) );
  NAND2_X1 U6551 ( .A1(n5354), .A2(n11031), .ZN(n5360) );
  XNOR2_X1 U6552 ( .A(instr_addr_o_22_), .B(n7289), .ZN(n5359) );
  INV_X1 U6553 ( .A(n5355), .ZN(n5357) );
  NOR2_X1 U6554 ( .A1(n5356), .A2(n544), .ZN(n11066) );
  NAND2_X1 U6555 ( .A1(n11066), .A2(pmp_addr_i[233]), .ZN(n11043) );
  NAND2_X1 U6556 ( .A1(n5357), .A2(n11043), .ZN(n5358) );
  NAND4_X1 U6557 ( .A1(n5361), .A2(n5360), .A3(n5359), .A4(n5358), .ZN(n5362)
         );
  NOR2_X1 U6558 ( .A1(n5363), .A2(n5362), .ZN(n5413) );
  XNOR2_X1 U6559 ( .A(n4556), .B(n7255), .ZN(n5367) );
  XNOR2_X1 U6560 ( .A(n5365), .B(n7257), .ZN(n5366) );
  XNOR2_X1 U6561 ( .A(n4533), .B(n7296), .ZN(n5372) );
  XNOR2_X1 U6562 ( .A(n5980), .B(n7247), .ZN(n5371) );
  XNOR2_X1 U6563 ( .A(n138), .B(n7295), .ZN(n5370) );
  XNOR2_X1 U6564 ( .A(n210), .B(n7258), .ZN(n5369) );
  NAND4_X1 U6565 ( .A1(n5372), .A2(n5371), .A3(n5370), .A4(n5369), .ZN(n5373)
         );
  XNOR2_X1 U6566 ( .A(instr_addr_o_31_), .B(n7309), .ZN(n5382) );
  INV_X1 U6567 ( .A(n5374), .ZN(n5376) );
  INV_X1 U6568 ( .A(n11066), .ZN(n5375) );
  NAND2_X1 U6569 ( .A1(n5376), .A2(n5375), .ZN(n5381) );
  INV_X1 U6570 ( .A(n5377), .ZN(n5379) );
  INV_X1 U6571 ( .A(n11057), .ZN(n5378) );
  NAND2_X1 U6572 ( .A1(n5379), .A2(n5378), .ZN(n5380) );
  NAND4_X1 U6573 ( .A1(n5383), .A2(n5382), .A3(n5381), .A4(n5380), .ZN(n5395)
         );
  INV_X1 U6574 ( .A(n5384), .ZN(n11052) );
  INV_X1 U6575 ( .A(n5385), .ZN(n5386) );
  OAI211_X1 U6576 ( .C1(n11052), .C2(n5388), .A(n5387), .B(n5386), .ZN(n5394)
         );
  OR2_X1 U6577 ( .A1(n11043), .A2(n5389), .ZN(n11055) );
  NOR2_X1 U6578 ( .A1(n11055), .A2(n5390), .ZN(n11073) );
  XNOR2_X1 U6579 ( .A(instr_addr_o_23_), .B(n7249), .ZN(n5391) );
  OAI21_X1 U6580 ( .B1(n5392), .B2(n11073), .A(n5391), .ZN(n5393) );
  NOR3_X1 U6581 ( .A1(n5395), .A2(n5394), .A3(n5393), .ZN(n5411) );
  INV_X1 U6582 ( .A(n5396), .ZN(n5397) );
  NOR2_X1 U6583 ( .A1(n5398), .A2(n5397), .ZN(n5402) );
  XNOR2_X1 U6584 ( .A(n5550), .B(n7290), .ZN(n5401) );
  XNOR2_X1 U6585 ( .A(n6020), .B(n7248), .ZN(n5400) );
  XNOR2_X1 U6586 ( .A(n6019), .B(n7279), .ZN(n5399) );
  NAND4_X1 U6587 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n5409)
         );
  INV_X1 U6588 ( .A(n5403), .ZN(n5404) );
  NAND2_X1 U6589 ( .A1(n5404), .A2(n11055), .ZN(n5407) );
  INV_X1 U6590 ( .A(n5405), .ZN(n11072) );
  AOI21_X1 U6591 ( .B1(n5407), .B2(n5406), .A(n11072), .ZN(n5408) );
  NOR2_X1 U6592 ( .A1(n5409), .A2(n5408), .ZN(n5410) );
  NAND4_X1 U6593 ( .A1(n5413), .A2(n5412), .A3(n5411), .A4(n5410), .ZN(n5517)
         );
  INV_X1 U6594 ( .A(n5449), .ZN(n5416) );
  INV_X1 U6595 ( .A(n5453), .ZN(n5415) );
  INV_X1 U6596 ( .A(n5414), .ZN(n11867) );
  AOI22_X1 U6597 ( .A1(n5416), .A2(n11852), .B1(n5415), .B2(n11867), .ZN(n5432) );
  INV_X1 U6598 ( .A(n5452), .ZN(n5419) );
  INV_X1 U6599 ( .A(n5460), .ZN(n5418) );
  INV_X1 U6600 ( .A(n5417), .ZN(n11824) );
  NAND3_X1 U6602 ( .A1(instr_addr_o_13_), .A2(n5420), .A3(n11828), .ZN(n5423)
         );
  NAND3_X1 U6603 ( .A1(n5057), .A2(n5421), .A3(n11870), .ZN(n5422) );
  OAI211_X1 U6604 ( .C1(n5459), .C2(n11838), .A(n5423), .B(n5422), .ZN(n5424)
         );
  INV_X1 U6605 ( .A(n5424), .ZN(n5430) );
  INV_X1 U6606 ( .A(n5458), .ZN(n5428) );
  INV_X1 U6607 ( .A(n5425), .ZN(n5426) );
  NAND2_X1 U6608 ( .A1(n5427), .A2(n5426), .ZN(n11846) );
  OAI21_X1 U6609 ( .B1(n5428), .B2(n11831), .A(n11846), .ZN(n5429) );
  NAND2_X1 U6611 ( .A1(n12150), .A2(n6983), .ZN(n5456) );
  INV_X1 U6612 ( .A(n11835), .ZN(n5437) );
  NAND3_X1 U6613 ( .A1(instr_addr_o_12_), .A2(n5433), .A3(n11862), .ZN(n5436)
         );
  OR2_X1 U6614 ( .A1(n11870), .A2(n5434), .ZN(n11820) );
  INV_X1 U6618 ( .A(n5447), .ZN(n5439) );
  OR2_X1 U6619 ( .A1(n11846), .A2(n89), .ZN(n11858) );
  NAND2_X1 U6620 ( .A1(n5439), .A2(n11858), .ZN(n5444) );
  INV_X1 U6621 ( .A(n5446), .ZN(n5440) );
  OAI21_X1 U6622 ( .B1(n2311), .B2(n11858), .A(n5440), .ZN(n5443) );
  INV_X1 U6623 ( .A(n5457), .ZN(n5441) );
  NAND2_X1 U6624 ( .A1(n5441), .A2(n11850), .ZN(n5442) );
  NAND4_X1 U6625 ( .A1(n12186), .A2(n5444), .A3(n5443), .A4(n5442), .ZN(n5467)
         );
  NAND4_X1 U6626 ( .A1(n5449), .A2(n5448), .A3(n5447), .A4(n5446), .ZN(n5455)
         );
  NOR2_X1 U6627 ( .A1(n5455), .A2(n5454), .ZN(n5465) );
  NAND3_X1 U6628 ( .A1(n5457), .A2(n6985), .A3(n5456), .ZN(n5463) );
  NAND4_X1 U6629 ( .A1(n5461), .A2(n5460), .A3(n5459), .A4(n5458), .ZN(n5462)
         );
  NOR2_X1 U6630 ( .A1(n5463), .A2(n5462), .ZN(n5464) );
  NAND2_X1 U6631 ( .A1(n5465), .A2(n5464), .ZN(n5466) );
  OAI21_X1 U6632 ( .B1(n5468), .B2(n5467), .A(n5466), .ZN(n5515) );
  OR2_X1 U6633 ( .A1(n5469), .A2(n6935), .ZN(n7009) );
  AND3_X1 U6634 ( .A1(n7009), .A2(n5470), .A3(pmp_cfg_i[74]), .ZN(n5471) );
  OAI21_X1 U6635 ( .B1(n5976), .B2(n6983), .A(n5471), .ZN(n5472) );
  NOR2_X1 U6636 ( .A1(n5473), .A2(n5472), .ZN(n5477) );
  XNOR2_X1 U6637 ( .A(n5550), .B(n6971), .ZN(n5476) );
  XNOR2_X1 U6638 ( .A(n137), .B(n6963), .ZN(n5475) );
  XNOR2_X1 U6639 ( .A(n4556), .B(n6969), .ZN(n5474) );
  NAND4_X1 U6640 ( .A1(n5477), .A2(n5476), .A3(n5475), .A4(n5474), .ZN(n5483)
         );
  XNOR2_X1 U6641 ( .A(n4908), .B(n6948), .ZN(n5481) );
  XNOR2_X1 U6642 ( .A(n6020), .B(n6953), .ZN(n5480) );
  XNOR2_X1 U6643 ( .A(n4533), .B(n6955), .ZN(n5479) );
  XNOR2_X1 U6644 ( .A(n5985), .B(n6964), .ZN(n5478) );
  NAND4_X1 U6645 ( .A1(n5481), .A2(n5480), .A3(n5479), .A4(n5478), .ZN(n5482)
         );
  NOR2_X1 U6646 ( .A1(n5483), .A2(n5482), .ZN(n5514) );
  INV_X1 U6647 ( .A(n5484), .ZN(n5490) );
  XNOR2_X1 U6648 ( .A(n6027), .B(n6954), .ZN(n5486) );
  XNOR2_X1 U6649 ( .A(n5330), .B(n6962), .ZN(n5485) );
  AND2_X1 U6650 ( .A1(n5486), .A2(n5485), .ZN(n5489) );
  XNOR2_X1 U6651 ( .A(n12199), .B(n6972), .ZN(n5488) );
  XNOR2_X1 U6652 ( .A(n146), .B(n6970), .ZN(n5487) );
  AND4_X1 U6653 ( .A1(n5490), .A2(n5489), .A3(n5488), .A4(n5487), .ZN(n5513)
         );
  NOR2_X1 U6654 ( .A1(n5492), .A2(n5491), .ZN(n5501) );
  NOR2_X1 U6655 ( .A1(n5494), .A2(n5493), .ZN(n5500) );
  INV_X1 U6656 ( .A(n5495), .ZN(n5497) );
  NOR2_X1 U6657 ( .A1(n5497), .A2(n5496), .ZN(n5499) );
  XNOR2_X1 U6658 ( .A(instr_addr_o_31_), .B(n7004), .ZN(n5498) );
  NAND4_X1 U6659 ( .A1(n5501), .A2(n5500), .A3(n5499), .A4(n5498), .ZN(n5511)
         );
  NOR2_X1 U6660 ( .A1(n5503), .A2(n5502), .ZN(n5509) );
  NOR2_X1 U6661 ( .A1(n5505), .A2(n5504), .ZN(n5508) );
  XNOR2_X1 U6662 ( .A(instr_addr_o_22_), .B(n6956), .ZN(n5507) );
  XNOR2_X1 U6663 ( .A(n5208), .B(n6961), .ZN(n5506) );
  NAND4_X1 U6664 ( .A1(n5509), .A2(n5508), .A3(n5507), .A4(n5506), .ZN(n5510)
         );
  NOR2_X1 U6665 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  NAND4_X1 U6666 ( .A1(n5515), .A2(n5514), .A3(n5513), .A4(n5512), .ZN(n5516)
         );
  AND2_X1 U6667 ( .A1(n5516), .A2(n5517), .ZN(n6044) );
  INV_X1 U6668 ( .A(n5518), .ZN(n5523) );
  INV_X1 U6669 ( .A(n5519), .ZN(n5522) );
  INV_X1 U6670 ( .A(n5520), .ZN(n5521) );
  AND4_X1 U6671 ( .A1(n5524), .A2(n5523), .A3(n5522), .A4(n5521), .ZN(n5541)
         );
  INV_X1 U6672 ( .A(n5525), .ZN(n5528) );
  XNOR2_X1 U6673 ( .A(n6025), .B(n9594), .ZN(n5526) );
  NAND3_X1 U6674 ( .A1(n5528), .A2(n5527), .A3(n5526), .ZN(n5535) );
  INV_X1 U6675 ( .A(n5529), .ZN(n5533) );
  XNOR2_X1 U6676 ( .A(instr_addr_o_22_), .B(n9624), .ZN(n5532) );
  INV_X1 U6677 ( .A(n5530), .ZN(n5531) );
  NAND3_X1 U6678 ( .A1(n5533), .A2(n5532), .A3(n5531), .ZN(n5534) );
  NOR2_X1 U6679 ( .A1(n5535), .A2(n5534), .ZN(n5540) );
  XNOR2_X1 U6680 ( .A(instr_addr_o_31_), .B(n9635), .ZN(n5539) );
  NOR2_X1 U6681 ( .A1(n5537), .A2(n5536), .ZN(n5538) );
  NAND4_X1 U6682 ( .A1(n5541), .A2(n5540), .A3(n5539), .A4(n5538), .ZN(n5566)
         );
  XNOR2_X1 U6683 ( .A(n6019), .B(n9596), .ZN(n5545) );
  XNOR2_X1 U6684 ( .A(instr_addr_o_21_), .B(n9625), .ZN(n5544) );
  XNOR2_X1 U6685 ( .A(n5985), .B(n9589), .ZN(n5543) );
  XNOR2_X1 U6686 ( .A(n6020), .B(n9595), .ZN(n5542) );
  OR2_X1 U6687 ( .A1(n12224), .A2(n9584), .ZN(n9658) );
  NAND3_X1 U6688 ( .A1(n9658), .A2(n5547), .A3(pmp_cfg_i[34]), .ZN(n5548) );
  AOI21_X1 U6689 ( .B1(n3876), .B2(n9475), .A(n5548), .ZN(n5553) );
  INV_X1 U6690 ( .A(n5549), .ZN(n5552) );
  XNOR2_X1 U6691 ( .A(n5550), .B(n9632), .ZN(n5551) );
  AND3_X1 U6692 ( .A1(n5553), .A2(n5552), .A3(n5551), .ZN(n5556) );
  XNOR2_X1 U6693 ( .A(n5202), .B(n9618), .ZN(n5555) );
  XNOR2_X1 U6694 ( .A(n4556), .B(n9586), .ZN(n5554) );
  INV_X1 U6695 ( .A(n5557), .ZN(n5563) );
  XNOR2_X1 U6696 ( .A(instr_addr_o_20_), .B(n9588), .ZN(n5559) );
  XNOR2_X1 U6697 ( .A(n6028), .B(n9587), .ZN(n5558) );
  AND2_X1 U6698 ( .A1(n5559), .A2(n5558), .ZN(n5562) );
  XNOR2_X1 U6699 ( .A(n5980), .B(n9597), .ZN(n5561) );
  XNOR2_X1 U6700 ( .A(n146), .B(n9619), .ZN(n5560) );
  NAND4_X1 U6701 ( .A1(n5563), .A2(n5562), .A3(n5561), .A4(n5560), .ZN(n5564)
         );
  NOR3_X1 U6702 ( .A1(n5566), .A2(n5565), .A3(n5564), .ZN(n5730) );
  INV_X1 U6703 ( .A(n5612), .ZN(n5571) );
  INV_X1 U6704 ( .A(n5587), .ZN(n11934) );
  NAND2_X1 U6705 ( .A1(n11934), .A2(pmp_addr_i[138]), .ZN(n5568) );
  OR2_X1 U6706 ( .A1(n5568), .A2(n5567), .ZN(n11894) );
  NOR2_X1 U6707 ( .A1(n11894), .A2(n5569), .ZN(n5575) );
  NAND2_X1 U6708 ( .A1(n5575), .A2(pmp_addr_i[140]), .ZN(n11880) );
  INV_X1 U6709 ( .A(n5602), .ZN(n5570) );
  AOI22_X1 U6710 ( .A1(n5571), .A2(n11880), .B1(n5570), .B2(n11894), .ZN(n5585) );
  INV_X1 U6711 ( .A(n5601), .ZN(n5574) );
  INV_X1 U6712 ( .A(n11901), .ZN(n5573) );
  INV_X1 U6713 ( .A(n5600), .ZN(n5572) );
  AOI22_X1 U6714 ( .A1(n5574), .A2(n5573), .B1(n5572), .B2(n11904), .ZN(n5584)
         );
  INV_X1 U6715 ( .A(n5607), .ZN(n5577) );
  INV_X1 U6716 ( .A(n5606), .ZN(n5576) );
  INV_X1 U6717 ( .A(n5575), .ZN(n11891) );
  AOI22_X1 U6718 ( .A1(n5577), .A2(n11929), .B1(n5576), .B2(n11891), .ZN(n5583) );
  INV_X1 U6719 ( .A(n5605), .ZN(n5581) );
  INV_X1 U6720 ( .A(n5604), .ZN(n5580) );
  INV_X1 U6721 ( .A(n11894), .ZN(n5579) );
  NAND2_X1 U6722 ( .A1(n5579), .A2(n5578), .ZN(n11882) );
  AOI22_X1 U6723 ( .A1(n5581), .A2(n11916), .B1(n5580), .B2(n11882), .ZN(n5582) );
  NAND4_X1 U6724 ( .A1(n5585), .A2(n5584), .A3(n5583), .A4(n5582), .ZN(n5623)
         );
  INV_X1 U6725 ( .A(n5616), .ZN(n5588) );
  INV_X1 U6726 ( .A(n5614), .ZN(n5586) );
  AOI22_X1 U6727 ( .A1(n5588), .A2(n5587), .B1(n5586), .B2(n11921), .ZN(n5599)
         );
  NAND2_X1 U6728 ( .A1(n12150), .A2(n9639), .ZN(n5610) );
  INV_X1 U6729 ( .A(n5610), .ZN(n5590) );
  INV_X1 U6730 ( .A(n5613), .ZN(n5589) );
  AOI22_X1 U6731 ( .A1(n5590), .A2(n11910), .B1(n5589), .B2(n11897), .ZN(n5598) );
  INV_X1 U6732 ( .A(n5603), .ZN(n5592) );
  INV_X1 U6733 ( .A(n5591), .ZN(n11903) );
  NAND2_X1 U6734 ( .A1(n5592), .A2(n11903), .ZN(n5597) );
  INV_X1 U6735 ( .A(n5615), .ZN(n5595) );
  INV_X1 U6736 ( .A(n11907), .ZN(n5594) );
  INV_X1 U6737 ( .A(n11882), .ZN(n5593) );
  NAND2_X1 U6738 ( .A1(n5593), .A2(pmp_addr_i[142]), .ZN(n11889) );
  OAI21_X1 U6739 ( .B1(n5595), .B2(n5594), .A(n11889), .ZN(n5596) );
  NAND4_X1 U6740 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), .ZN(n5622)
         );
  NAND4_X1 U6741 ( .A1(n5603), .A2(n5602), .A3(n5601), .A4(n5600), .ZN(n5609)
         );
  NAND4_X1 U6742 ( .A1(n5607), .A2(n5606), .A3(n5605), .A4(n5604), .ZN(n5608)
         );
  NOR2_X1 U6743 ( .A1(n5609), .A2(n5608), .ZN(n5620) );
  INV_X1 U6744 ( .A(n9638), .ZN(n5611) );
  NAND3_X1 U6745 ( .A1(n5612), .A2(n5611), .A3(n5610), .ZN(n5618) );
  NAND4_X1 U6746 ( .A1(n5616), .A2(n5615), .A3(n5614), .A4(n5613), .ZN(n5617)
         );
  NOR2_X1 U6747 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  NAND2_X1 U6748 ( .A1(n5620), .A2(n5619), .ZN(n5621) );
  OAI21_X1 U6749 ( .B1(n5623), .B2(n5622), .A(n5621), .ZN(n5729) );
  INV_X1 U6750 ( .A(n5624), .ZN(n5631) );
  INV_X1 U6751 ( .A(n5625), .ZN(n5630) );
  INV_X1 U6752 ( .A(n5626), .ZN(n5629) );
  INV_X1 U6753 ( .A(n5627), .ZN(n5628) );
  NAND4_X1 U6754 ( .A1(n5631), .A2(n5630), .A3(n5629), .A4(n5628), .ZN(n5635)
         );
  XNOR2_X1 U6755 ( .A(instr_addr_o_31_), .B(n5632), .ZN(n5633) );
  XNOR2_X1 U6756 ( .A(n5202), .B(n6306), .ZN(n5637) );
  XNOR2_X1 U6757 ( .A(n12207), .B(n6322), .ZN(n5636) );
  NAND2_X1 U6758 ( .A1(n5637), .A2(n5636), .ZN(n5642) );
  XNOR2_X1 U6759 ( .A(instr_addr_o_28_), .B(n6319), .ZN(n5640) );
  XNOR2_X1 U6760 ( .A(instr_addr_o_20_), .B(n6314), .ZN(n5639) );
  XNOR2_X1 U6761 ( .A(n6028), .B(n6304), .ZN(n5638) );
  NAND3_X1 U6762 ( .A1(n5640), .A2(n5639), .A3(n5638), .ZN(n5641) );
  NOR2_X1 U6763 ( .A1(n5642), .A2(n5641), .ZN(n5654) );
  INV_X1 U6764 ( .A(n5643), .ZN(n5645) );
  XNOR2_X1 U6765 ( .A(n6025), .B(n6303), .ZN(n5644) );
  NAND3_X1 U6766 ( .A1(n5646), .A2(n5645), .A3(n5644), .ZN(n5652) );
  INV_X1 U6767 ( .A(n5647), .ZN(n5650) );
  XNOR2_X1 U6768 ( .A(instr_addr_o_22_), .B(n6311), .ZN(n5649) );
  NAND3_X1 U6769 ( .A1(n5650), .A2(n5649), .A3(n5648), .ZN(n5651) );
  NOR2_X1 U6770 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  NAND3_X1 U6771 ( .A1(n5655), .A2(n5654), .A3(n5653), .ZN(n5674) );
  NOR2_X1 U6772 ( .A1(n5657), .A2(n5656), .ZN(n5661) );
  XNOR2_X1 U6773 ( .A(n5183), .B(n6310), .ZN(n5660) );
  XNOR2_X1 U6774 ( .A(n6020), .B(n6313), .ZN(n5659) );
  XNOR2_X1 U6775 ( .A(n6019), .B(n6236), .ZN(n5658) );
  NAND4_X1 U6776 ( .A1(n5661), .A2(n5660), .A3(n5659), .A4(n5658), .ZN(n5673)
         );
  NAND2_X1 U6777 ( .A1(n5663), .A2(n5662), .ZN(n6051) );
  AND3_X1 U6778 ( .A1(n6051), .A2(n5664), .A3(pmp_cfg_i[18]), .ZN(n5665) );
  OAI21_X1 U6779 ( .B1(n5976), .B2(n6258), .A(n5665), .ZN(n5666) );
  NOR2_X1 U6780 ( .A1(n5667), .A2(n5666), .ZN(n5671) );
  XNOR2_X1 U6781 ( .A(n5985), .B(n6307), .ZN(n5670) );
  XNOR2_X1 U6782 ( .A(n5550), .B(n6321), .ZN(n5669) );
  XNOR2_X1 U6783 ( .A(n4556), .B(n6318), .ZN(n5668) );
  NAND4_X1 U6784 ( .A1(n5671), .A2(n5670), .A3(n5669), .A4(n5668), .ZN(n5672)
         );
  NOR3_X1 U6785 ( .A1(n5674), .A2(n5673), .A3(n5672), .ZN(n5728) );
  AND2_X1 U6786 ( .A1(n5675), .A2(n5699), .ZN(n5722) );
  NOR2_X1 U6787 ( .A1(n11151), .A2(n2039), .ZN(n11165) );
  NAND2_X1 U6788 ( .A1(n11165), .A2(pmp_addr_i[67]), .ZN(n11167) );
  OR2_X1 U6789 ( .A1(n11167), .A2(n5676), .ZN(n11162) );
  INV_X1 U6790 ( .A(n5677), .ZN(n5678) );
  OR2_X1 U6791 ( .A1(n11162), .A2(n5678), .ZN(n11192) );
  INV_X1 U6792 ( .A(n11192), .ZN(n5696) );
  INV_X1 U6793 ( .A(n5711), .ZN(n5684) );
  NOR2_X1 U6794 ( .A1(n11162), .A2(n5679), .ZN(n11177) );
  NAND2_X1 U6795 ( .A1(n11177), .A2(pmp_addr_i[70]), .ZN(n5704) );
  NAND3_X1 U6796 ( .A1(n12267), .A2(n6093), .A3(n11162), .ZN(n5682) );
  INV_X1 U6797 ( .A(n11165), .ZN(n5680) );
  NAND3_X1 U6798 ( .A1(instr_addr_o_5_), .A2(n6095), .A3(n5680), .ZN(n5681) );
  NAND3_X1 U6799 ( .A1(n5682), .A2(n11155), .A3(n5681), .ZN(n5683) );
  AOI21_X1 U6800 ( .B1(n5684), .B2(n5704), .A(n5683), .ZN(n5690) );
  NOR2_X1 U6801 ( .A1(n11192), .A2(n5685), .ZN(n11176) );
  AND2_X1 U6802 ( .A1(n11176), .A2(pmp_addr_i[75]), .ZN(n5686) );
  INV_X1 U6803 ( .A(n5686), .ZN(n11185) );
  OR2_X1 U6804 ( .A1(n5686), .A2(n6244), .ZN(n11183) );
  OAI21_X1 U6805 ( .B1(instr_addr_o_14__BAR), .B2(n11183), .A(n5720), .ZN(
        n5688) );
  OAI21_X1 U6806 ( .B1(n2056), .B2(n11185), .A(n5688), .ZN(n5689) );
  OAI211_X1 U6807 ( .C1(n5722), .C2(n5696), .A(n5690), .B(n5689), .ZN(n5727)
         );
  INV_X1 U6808 ( .A(n5721), .ZN(n5693) );
  INV_X1 U6809 ( .A(n11176), .ZN(n5692) );
  INV_X1 U6810 ( .A(n5719), .ZN(n5691) );
  AOI22_X1 U6811 ( .A1(n5693), .A2(n5692), .B1(n5691), .B2(n11167), .ZN(n5709)
         );
  INV_X1 U6812 ( .A(n5694), .ZN(n5698) );
  INV_X1 U6813 ( .A(n11177), .ZN(n5697) );
  NAND2_X1 U6814 ( .A1(n5696), .A2(n5695), .ZN(n11193) );
  INV_X1 U6815 ( .A(n5699), .ZN(n5702) );
  INV_X1 U6816 ( .A(n5714), .ZN(n5701) );
  INV_X1 U6817 ( .A(n11193), .ZN(n5700) );
  NAND2_X1 U6818 ( .A1(n5700), .A2(pmp_addr_i[78]), .ZN(n11198) );
  AOI22_X1 U6819 ( .A1(n5702), .A2(n2068), .B1(n5701), .B2(n11198), .ZN(n5707)
         );
  INV_X1 U6820 ( .A(n5703), .ZN(n5705) );
  INV_X1 U6821 ( .A(n5704), .ZN(n11173) );
  NAND2_X1 U6822 ( .A1(n11173), .A2(pmp_addr_i[71]), .ZN(n11148) );
  AND2_X1 U6823 ( .A1(n12150), .A2(n6258), .ZN(n5712) );
  AOI22_X1 U6824 ( .A1(n5705), .A2(n11148), .B1(n5712), .B2(n11151), .ZN(n5706) );
  NAND4_X1 U6825 ( .A1(n5709), .A2(n5708), .A3(n5707), .A4(n5706), .ZN(n5726)
         );
  NAND3_X1 U6826 ( .A1(n5711), .A2(n6096), .A3(n5710), .ZN(n5717) );
  INV_X1 U6827 ( .A(n5712), .ZN(n5713) );
  AND4_X1 U6828 ( .A1(n5721), .A2(n5720), .A3(n5719), .A4(n5718), .ZN(n5724)
         );
  INV_X1 U6829 ( .A(n11603), .ZN(n5731) );
  OAI22_X1 U6830 ( .A1(n11583), .A2(n5766), .B1(n5777), .B2(n5731), .ZN(n5748)
         );
  INV_X1 U6831 ( .A(n5732), .ZN(n5733) );
  OR2_X1 U6832 ( .A1(n11595), .A2(n5733), .ZN(n11613) );
  NOR2_X1 U6833 ( .A1(n11613), .A2(n1792), .ZN(n5750) );
  INV_X1 U6834 ( .A(n5750), .ZN(n11620) );
  INV_X1 U6835 ( .A(n5734), .ZN(n11616) );
  NOR2_X1 U6836 ( .A1(n11620), .A2(n11616), .ZN(n5746) );
  NAND2_X1 U6837 ( .A1(n5750), .A2(pmp_addr_i[259]), .ZN(n5757) );
  OR2_X1 U6838 ( .A1(n5757), .A2(n5735), .ZN(n11633) );
  INV_X1 U6839 ( .A(n11633), .ZN(n5736) );
  NOR2_X1 U6840 ( .A1(n5736), .A2(n8857), .ZN(n5739) );
  NOR2_X1 U6841 ( .A1(n11633), .A2(n5737), .ZN(n11635) );
  NOR2_X1 U6842 ( .A1(n11635), .A2(n8856), .ZN(n5738) );
  AOI22_X1 U6843 ( .A1(n5740), .A2(n5739), .B1(n6005), .B2(n5738), .ZN(n5745)
         );
  INV_X1 U6844 ( .A(n5741), .ZN(n5743) );
  NAND2_X1 U6845 ( .A1(n8974), .A2(n5741), .ZN(n5742) );
  OAI211_X1 U6846 ( .C1(n12150), .C2(n5743), .A(n11613), .B(n5742), .ZN(n5744)
         );
  OAI211_X1 U6847 ( .C1(n5765), .C2(n5746), .A(n5745), .B(n5744), .ZN(n5747)
         );
  NOR2_X1 U6848 ( .A1(n5748), .A2(n5747), .ZN(n5762) );
  NOR2_X1 U6849 ( .A1(n11586), .A2(n1819), .ZN(n11585) );
  INV_X1 U6850 ( .A(n5749), .ZN(n11626) );
  OAI22_X1 U6851 ( .A1(n11585), .A2(n5776), .B1(n5775), .B2(n11626), .ZN(n5753) );
  INV_X1 U6852 ( .A(n11618), .ZN(n5751) );
  OAI22_X1 U6853 ( .A1(n5751), .A2(n5774), .B1(n5773), .B2(n5750), .ZN(n5752)
         );
  NOR2_X1 U6854 ( .A1(n5753), .A2(n5752), .ZN(n5761) );
  INV_X1 U6855 ( .A(n5770), .ZN(n5755) );
  INV_X1 U6856 ( .A(n5768), .ZN(n5754) );
  AOI22_X1 U6857 ( .A1(n5755), .A2(n11587), .B1(n5754), .B2(n11605), .ZN(n5760) );
  INV_X1 U6858 ( .A(n5764), .ZN(n5758) );
  INV_X1 U6859 ( .A(n5763), .ZN(n5756) );
  AOI22_X1 U6860 ( .A1(n5758), .A2(n5757), .B1(n5756), .B2(n11586), .ZN(n5759)
         );
  NAND4_X1 U6861 ( .A1(n5762), .A2(n5761), .A3(n5760), .A4(n5759), .ZN(n5782)
         );
  NAND4_X1 U6862 ( .A1(n5766), .A2(n5765), .A3(n5764), .A4(n5763), .ZN(n5772)
         );
  NAND4_X1 U6863 ( .A1(n5770), .A2(n5769), .A3(n5768), .A4(n5767), .ZN(n5771)
         );
  NOR2_X1 U6864 ( .A1(n5772), .A2(n5771), .ZN(n5780) );
  AOI21_X1 U6865 ( .B1(n5899), .B2(n5786), .A(n9009), .ZN(n5779) );
  AND4_X1 U6866 ( .A1(n5776), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(n5778)
         );
  NAND4_X1 U6867 ( .A1(n5780), .A2(n5779), .A3(n5778), .A4(n5777), .ZN(n5781)
         );
  NAND2_X1 U6868 ( .A1(n5782), .A2(n5781), .ZN(n5828) );
  AND3_X1 U6869 ( .A1(n5783), .A2(n5784), .A3(pmp_cfg_i[66]), .ZN(n5785) );
  OAI21_X1 U6870 ( .B1(n5976), .B2(n5786), .A(n5785), .ZN(n5787) );
  NOR2_X1 U6871 ( .A1(n5788), .A2(n5787), .ZN(n5792) );
  XNOR2_X1 U6872 ( .A(n5550), .B(n9002), .ZN(n5791) );
  XNOR2_X1 U6873 ( .A(n4556), .B(n8960), .ZN(n5790) );
  XNOR2_X1 U6874 ( .A(instr_addr_o_25_), .B(n8996), .ZN(n5789) );
  NAND4_X1 U6875 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(n5798)
         );
  XNOR2_X1 U6876 ( .A(instr_addr_o_21_), .B(n8985), .ZN(n5796) );
  XNOR2_X1 U6877 ( .A(n6020), .B(n8953), .ZN(n5795) );
  XNOR2_X1 U6878 ( .A(n6019), .B(n8961), .ZN(n5794) );
  XNOR2_X1 U6879 ( .A(n5985), .B(n8950), .ZN(n5793) );
  NAND4_X1 U6880 ( .A1(n5796), .A2(n5795), .A3(n5794), .A4(n5793), .ZN(n5797)
         );
  NOR2_X1 U6881 ( .A1(n5798), .A2(n5797), .ZN(n5827) );
  INV_X1 U6882 ( .A(n5799), .ZN(n5805) );
  INV_X1 U6883 ( .A(n5800), .ZN(n5804) );
  INV_X1 U6884 ( .A(n5801), .ZN(n5802) );
  AND4_X1 U6885 ( .A1(n5805), .A2(n5804), .A3(n5803), .A4(n5802), .ZN(n5818)
         );
  INV_X1 U6886 ( .A(n5806), .ZN(n5809) );
  XNOR2_X1 U6887 ( .A(n6025), .B(n8958), .ZN(n5807) );
  INV_X1 U6888 ( .A(n5810), .ZN(n5813) );
  XNOR2_X1 U6889 ( .A(instr_addr_o_22_), .B(n8959), .ZN(n5812) );
  INV_X1 U6890 ( .A(n1744), .ZN(n5811) );
  XNOR2_X1 U6891 ( .A(instr_addr_o_31_), .B(n9007), .ZN(n5817) );
  NOR2_X1 U6892 ( .A1(n5815), .A2(n5814), .ZN(n5816) );
  INV_X1 U6893 ( .A(n5819), .ZN(n5825) );
  XNOR2_X1 U6894 ( .A(instr_addr_o_20_), .B(n9001), .ZN(n5821) );
  XNOR2_X1 U6895 ( .A(n6028), .B(n8995), .ZN(n5820) );
  AND2_X1 U6896 ( .A1(n5821), .A2(n5820), .ZN(n5824) );
  XNOR2_X1 U6897 ( .A(n4753), .B(n8952), .ZN(n5823) );
  XNOR2_X1 U6898 ( .A(n146), .B(n8951), .ZN(n5822) );
  XNOR2_X1 U6899 ( .A(n4802), .B(n10979), .ZN(n5830) );
  XNOR2_X1 U6900 ( .A(instr_addr_o_24_), .B(n10987), .ZN(n5829) );
  AND2_X1 U6901 ( .A1(n5830), .A2(n5829), .ZN(n5832) );
  XNOR2_X1 U6902 ( .A(n146), .B(n10973), .ZN(n5831) );
  NAND4_X1 U6903 ( .A1(n5834), .A2(n5833), .A3(n5832), .A4(n5831), .ZN(n5856)
         );
  INV_X1 U6904 ( .A(n5835), .ZN(n5836) );
  NOR2_X1 U6905 ( .A1(n5837), .A2(n5836), .ZN(n5846) );
  INV_X1 U6906 ( .A(n5838), .ZN(n5840) );
  NOR2_X1 U6907 ( .A1(n5840), .A2(n5839), .ZN(n5845) );
  XNOR2_X1 U6908 ( .A(instr_addr_o_31_), .B(n11007), .ZN(n5844) );
  XNOR2_X1 U6909 ( .A(instr_addr_o_21_), .B(n10980), .ZN(n5843) );
  NAND4_X1 U6910 ( .A1(n5846), .A2(n5845), .A3(n5844), .A4(n5843), .ZN(n5855)
         );
  XNOR2_X1 U6911 ( .A(instr_addr_o_22_), .B(n10981), .ZN(n5852) );
  NOR2_X1 U6912 ( .A1(n5849), .A2(n5848), .ZN(n5851) );
  XNOR2_X1 U6913 ( .A(n6025), .B(n10982), .ZN(n5850) );
  NAND4_X1 U6914 ( .A1(n5853), .A2(n5852), .A3(n5851), .A4(n5850), .ZN(n5854)
         );
  NOR3_X1 U6915 ( .A1(n5856), .A2(n5855), .A3(n5854), .ZN(n5927) );
  INV_X1 U6916 ( .A(n5857), .ZN(n5858) );
  OR2_X1 U6917 ( .A1(n11381), .A2(n5858), .ZN(n5879) );
  NOR2_X1 U6918 ( .A1(n5879), .A2(n5859), .ZN(n11375) );
  NAND2_X1 U6919 ( .A1(n11375), .A2(pmp_addr_i[164]), .ZN(n5878) );
  OR2_X1 U6920 ( .A1(n5878), .A2(n5860), .ZN(n11370) );
  INV_X1 U6921 ( .A(n5861), .ZN(n5862) );
  NOR2_X1 U6922 ( .A1(n11370), .A2(n5862), .ZN(n11364) );
  OAI21_X1 U6923 ( .B1(n5894), .B2(pmp_addr_i[173]), .A(n11364), .ZN(n5871) );
  INV_X1 U6924 ( .A(n11370), .ZN(n5863) );
  AOI21_X1 U6925 ( .B1(n5863), .B2(pmp_addr_i[171]), .A(n10809), .ZN(n5864) );
  NAND2_X1 U6926 ( .A1(instr_addr_o_14_), .A2(n5864), .ZN(n5865) );
  NAND3_X1 U6927 ( .A1(n5904), .A2(n5894), .A3(n5865), .ZN(n5870) );
  INV_X1 U6928 ( .A(pmp_addr_i[165]), .ZN(n5866) );
  OR2_X1 U6929 ( .A1(n5878), .A2(n5866), .ZN(n5872) );
  NOR2_X1 U6930 ( .A1(n5872), .A2(n5036), .ZN(n11361) );
  NAND2_X1 U6931 ( .A1(n11361), .A2(pmp_addr_i[167]), .ZN(n5875) );
  OR2_X1 U6932 ( .A1(n5875), .A2(n5867), .ZN(n11397) );
  NOR2_X1 U6933 ( .A1(n11397), .A2(n5868), .ZN(n11395) );
  OAI21_X1 U6934 ( .B1(n5903), .B2(n11395), .A(n5891), .ZN(n5869) );
  AOI22_X1 U6935 ( .A1(n5871), .A2(n5870), .B1(n5869), .B2(n11370), .ZN(n5888)
         );
  INV_X1 U6936 ( .A(n11397), .ZN(n5873) );
  INV_X1 U6937 ( .A(n5872), .ZN(n11362) );
  INV_X1 U6938 ( .A(n11364), .ZN(n5874) );
  NOR2_X1 U6939 ( .A1(n5874), .A2(n5056), .ZN(n11358) );
  AND2_X1 U6940 ( .A1(n11358), .A2(pmp_addr_i[174]), .ZN(n11392) );
  INV_X1 U6941 ( .A(n5875), .ZN(n11357) );
  OAI22_X1 U6942 ( .A1(n11392), .A2(n5902), .B1(n5901), .B2(n11357), .ZN(n5876) );
  NOR2_X1 U6943 ( .A1(n5877), .A2(n5876), .ZN(n5887) );
  INV_X1 U6944 ( .A(n5878), .ZN(n11386) );
  OAI22_X1 U6945 ( .A1(n11375), .A2(n5890), .B1(n5889), .B2(n11386), .ZN(n5885) );
  NAND2_X1 U6946 ( .A1(pmp_addr_i[160]), .A2(pmp_addr_i[161]), .ZN(n11380) );
  NAND3_X1 U6947 ( .A1(n12150), .A2(n5898), .A3(n11380), .ZN(n5883) );
  INV_X1 U6948 ( .A(n5880), .ZN(n11382) );
  INV_X1 U6949 ( .A(n5879), .ZN(n11372) );
  AOI21_X1 U6950 ( .B1(n5880), .B2(n10813), .A(n11372), .ZN(n5881) );
  OAI21_X1 U6951 ( .B1(n6015), .B2(n11382), .A(n5881), .ZN(n5882) );
  OAI211_X1 U6952 ( .C1(n5892), .C2(n11361), .A(n5883), .B(n5882), .ZN(n5884)
         );
  NAND4_X1 U6955 ( .A1(n5892), .A2(n5891), .A3(n5890), .A4(n5889), .ZN(n5897)
         );
  NOR2_X1 U6956 ( .A1(n5897), .A2(n5896), .ZN(n5907) );
  AOI21_X1 U6957 ( .B1(n5899), .B2(n5898), .A(pmp_cfg_i[43]), .ZN(n5906) );
  AND4_X1 U6958 ( .A1(n5903), .A2(n5902), .A3(n5901), .A4(n5900), .ZN(n5905)
         );
  NAND4_X1 U6959 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(n5908)
         );
  NAND2_X1 U6960 ( .A1(n5909), .A2(n5908), .ZN(n5926) );
  XNOR2_X1 U6961 ( .A(n6020), .B(n10968), .ZN(n5913) );
  XNOR2_X1 U6962 ( .A(gte_x_382_A_16_), .B(n10966), .ZN(n5912) );
  XNOR2_X1 U6963 ( .A(n5985), .B(n10989), .ZN(n5911) );
  XNOR2_X1 U6964 ( .A(n5550), .B(n11012), .ZN(n5910) );
  NAND4_X1 U6965 ( .A1(n5913), .A2(n5912), .A3(n5911), .A4(n5910), .ZN(n5924)
         );
  XNOR2_X1 U6966 ( .A(n4556), .B(n10990), .ZN(n5918) );
  OR2_X1 U6967 ( .A1(n5914), .A2(n161), .ZN(n11018) );
  NAND3_X1 U6968 ( .A1(n11018), .A2(n5915), .A3(pmp_cfg_i[42]), .ZN(n5916) );
  AOI21_X1 U6969 ( .B1(n3876), .B2(n10960), .A(n5916), .ZN(n5917) );
  NAND3_X1 U6970 ( .A1(n5919), .A2(n5918), .A3(n5917), .ZN(n5923) );
  XNOR2_X1 U6971 ( .A(n12226), .B(n10988), .ZN(n5921) );
  XNOR2_X1 U6972 ( .A(n5980), .B(n10974), .ZN(n5920) );
  NAND2_X1 U6973 ( .A1(n5921), .A2(n5920), .ZN(n5922) );
  NOR3_X1 U6974 ( .A1(n5924), .A2(n5923), .A3(n5922), .ZN(n5925) );
  NAND3_X1 U6975 ( .A1(n5927), .A2(n5926), .A3(n5925), .ZN(n6040) );
  INV_X1 U6976 ( .A(n5967), .ZN(n5930) );
  INV_X1 U6977 ( .A(n5931), .ZN(n5929) );
  INV_X1 U6978 ( .A(n12021), .ZN(n5928) );
  AOI22_X1 U6979 ( .A1(n5930), .A2(n12008), .B1(n5929), .B2(n5928), .ZN(n5939)
         );
  OAI211_X1 U6980 ( .C1(n3839), .C2(n10307), .A(n5931), .B(n5932), .ZN(n5962)
         );
  NAND2_X1 U6981 ( .A1(n5962), .A2(n12042), .ZN(n5938) );
  INV_X1 U6982 ( .A(n5932), .ZN(n5936) );
  INV_X1 U6983 ( .A(n5968), .ZN(n5934) );
  OR2_X1 U6984 ( .A1(n12042), .A2(n5933), .ZN(n5942) );
  INV_X1 U6986 ( .A(n5960), .ZN(n5941) );
  INV_X1 U6987 ( .A(n5959), .ZN(n5940) );
  AOI22_X1 U6988 ( .A1(n5941), .A2(n12014), .B1(n5940), .B2(n12041), .ZN(n5956) );
  INV_X1 U6989 ( .A(n5958), .ZN(n5945) );
  INV_X1 U6990 ( .A(n5942), .ZN(n12039) );
  NAND2_X1 U6991 ( .A1(n12039), .A2(pmp_addr_i[357]), .ZN(n12025) );
  INV_X1 U6992 ( .A(n5957), .ZN(n5944) );
  INV_X1 U6993 ( .A(n12018), .ZN(n5943) );
  AOI22_X1 U6994 ( .A1(n5945), .A2(n12025), .B1(n5944), .B2(n5943), .ZN(n5955)
         );
  INV_X1 U6995 ( .A(n5966), .ZN(n5947) );
  INV_X1 U6996 ( .A(n5965), .ZN(n5946) );
  INV_X1 U6997 ( .A(n5964), .ZN(n5952) );
  INV_X1 U6998 ( .A(n5948), .ZN(n12028) );
  OR3_X1 U6999 ( .A1(n5951), .A2(n5950), .A3(n5949), .ZN(n12057) );
  OAI21_X1 U7000 ( .B1(n5952), .B2(n12028), .A(n12057), .ZN(n5953) );
  NAND4_X1 U7001 ( .A1(n5956), .A2(n5955), .A3(n5954), .A4(n5953), .ZN(n5972)
         );
  NAND4_X1 U7002 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n5961)
         );
  NOR2_X1 U7003 ( .A1(n5962), .A2(n5961), .ZN(n5970) );
  INV_X1 U7004 ( .A(n5963), .ZN(n10311) );
  AND4_X1 U7005 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n10311), .ZN(n5969)
         );
  NAND4_X1 U7006 ( .A1(n5970), .A2(n5969), .A3(n5968), .A4(n5967), .ZN(n5971)
         );
  OAI22_X1 U7007 ( .A1(instr_addr_o_12_), .A2(n10316), .B1(n4069), .B2(n5973), 
        .ZN(n5978) );
  OAI22_X1 U7008 ( .A1(instr_addr_o_10_), .A2(n10317), .B1(n5976), .B2(n12059), 
        .ZN(n5977) );
  NOR2_X1 U7009 ( .A1(n5978), .A2(n5977), .ZN(n5984) );
  XNOR2_X1 U7010 ( .A(n4556), .B(n10278), .ZN(n5983) );
  XNOR2_X1 U7011 ( .A(n146), .B(n10266), .ZN(n5982) );
  XNOR2_X1 U7012 ( .A(n4753), .B(n10258), .ZN(n5981) );
  NAND4_X1 U7013 ( .A1(n5984), .A2(n5983), .A3(n5982), .A4(n5981), .ZN(n5992)
         );
  XNOR2_X1 U7014 ( .A(n4533), .B(n10260), .ZN(n5990) );
  XNOR2_X1 U7015 ( .A(n5985), .B(n10268), .ZN(n5989) );
  XNOR2_X1 U7016 ( .A(n5202), .B(n10269), .ZN(n5988) );
  XNOR2_X1 U7017 ( .A(instr_addr_o_29_), .B(n10277), .ZN(n5987) );
  NAND4_X1 U7018 ( .A1(n5990), .A2(n5989), .A3(n5988), .A4(n5987), .ZN(n5991)
         );
  NOR2_X1 U7019 ( .A1(n5992), .A2(n5991), .ZN(n6037) );
  OAI21_X1 U7020 ( .B1(n5993), .B2(pmp_addr_i[365]), .A(n12024), .ZN(n5995) );
  OAI21_X1 U7021 ( .B1(n6017), .B2(n10280), .A(n5993), .ZN(n5994) );
  NAND2_X1 U7022 ( .A1(n5995), .A2(n5994), .ZN(n6010) );
  OAI22_X1 U7023 ( .A1(n5997), .A2(n10315), .B1(n154), .B2(n10305), .ZN(n6000)
         );
  OAI22_X1 U7024 ( .A1(instr_addr_o_6_), .A2(n10306), .B1(n12267), .B2(n10309), 
        .ZN(n5999) );
  NOR2_X1 U7025 ( .A1(n6000), .A2(n5999), .ZN(n6009) );
  OAI22_X1 U7026 ( .A1(n3934), .A2(n10318), .B1(n12180), .B2(n10314), .ZN(
        n6007) );
  OAI22_X1 U7027 ( .A1(instr_addr_o_8_), .A2(n10322), .B1(instr_addr_o_16_), 
        .B2(n6003), .ZN(n6006) );
  NOR2_X1 U7028 ( .A1(n6007), .A2(n6006), .ZN(n6008) );
  NAND3_X1 U7029 ( .A1(n6010), .A2(n6009), .A3(n6008), .ZN(n6035) );
  OR2_X1 U7030 ( .A1(n6011), .A2(n10256), .ZN(n10333) );
  AND4_X1 U7031 ( .A1(n10333), .A2(n10319), .A3(n6012), .A4(pmp_cfg_i[90]), 
        .ZN(n6013) );
  OAI21_X1 U7032 ( .B1(n6015), .B2(n6014), .A(n6013), .ZN(n6016) );
  AOI21_X1 U7033 ( .B1(n6017), .B2(n10280), .A(n6016), .ZN(n6024) );
  XNOR2_X1 U7034 ( .A(n6018), .B(n10304), .ZN(n6023) );
  XNOR2_X1 U7035 ( .A(n6019), .B(n10298), .ZN(n6022) );
  XNOR2_X1 U7036 ( .A(n6020), .B(n10261), .ZN(n6021) );
  NAND4_X1 U7037 ( .A1(n6024), .A2(n6023), .A3(n6022), .A4(n6021), .ZN(n6034)
         );
  XNOR2_X1 U7038 ( .A(n6025), .B(n10279), .ZN(n6032) );
  XNOR2_X1 U7039 ( .A(instr_addr_o_22_), .B(n10270), .ZN(n6031) );
  XNOR2_X1 U7040 ( .A(n6027), .B(n10296), .ZN(n6030) );
  XNOR2_X1 U7041 ( .A(n6028), .B(n10259), .ZN(n6029) );
  NAND4_X1 U7042 ( .A1(n6032), .A2(n6031), .A3(n6030), .A4(n6029), .ZN(n6033)
         );
  NOR3_X1 U7043 ( .A1(n6035), .A2(n6034), .A3(n6033), .ZN(n6036) );
  AND3_X1 U7044 ( .A1(n6041), .A2(n6040), .A3(n6039), .ZN(n6042) );
  NAND4_X1 U7045 ( .A1(n6045), .A2(n6044), .A3(n6043), .A4(n6042), .ZN(n12132)
         );
  NOR2_X1 U7046 ( .A1(n6047), .A2(n6046), .ZN(n6048) );
  NAND4_X1 U7047 ( .A1(n12135), .A2(n12198), .A3(n6049), .A4(n6048), .ZN(n6050) );
  INV_X1 U7048 ( .A(data_addr_i[15]), .ZN(n9941) );
  INV_X1 U7049 ( .A(n9941), .ZN(data_addr_o_15_) );
  BUF_X1 U7050 ( .A(data_addr_i[18]), .Z(n12260) );
  INV_X1 U7051 ( .A(data_addr_i[16]), .ZN(n8089) );
  INV_X1 U7052 ( .A(n8089), .ZN(data_addr_o_16_) );
  INV_X1 U7053 ( .A(data_addr_i[31]), .ZN(n9634) );
  INV_X1 U7054 ( .A(data_addr_i[17]), .ZN(n6688) );
  INV_X1 U7055 ( .A(n6688), .ZN(data_addr_o_17_) );
  INV_X1 U7056 ( .A(n12058), .ZN(data_addr_o_4_) );
  INV_X1 U7057 ( .A(data_addr_i[10]), .ZN(n7820) );
  INV_X1 U7058 ( .A(n11291), .ZN(data_addr_o_5_) );
  INV_X1 U7059 ( .A(data_addr_i[20]), .ZN(n10295) );
  INV_X1 U7060 ( .A(n10295), .ZN(data_addr_o_20_) );
  INV_X1 U7061 ( .A(data_addr_i[11]), .ZN(n7324) );
  INV_X1 U7062 ( .A(data_addr_i[8]), .ZN(n7814) );
  INV_X1 U7063 ( .A(data_addr_i[3]), .ZN(n10473) );
  INV_X1 U7064 ( .A(n10473), .ZN(data_addr_o_3_) );
  INV_X1 U7065 ( .A(data_we_i), .ZN(n11021) );
  INV_X1 U7066 ( .A(n11021), .ZN(n11019) );
  MUX2_X1 U7067 ( .A(pmp_cfg_i[16]), .B(pmp_cfg_i[17]), .S(n11019), .Z(n6052)
         );
  AND2_X1 U7068 ( .A1(n6051), .A2(n6052), .ZN(n11154) );
  BUF_X1 U7069 ( .A(data_addr_i[19]), .Z(n10627) );
  XNOR2_X1 U7070 ( .A(n10627), .B(n6313), .ZN(n6056) );
  XNOR2_X1 U7071 ( .A(n11285), .B(n6314), .ZN(n6055) );
  XNOR2_X1 U7073 ( .A(data_addr_o_30_), .B(n6322), .ZN(n6054) );
  XNOR2_X1 U7074 ( .A(n12260), .B(n6236), .ZN(n6053) );
  NAND4_X1 U7075 ( .A1(n6056), .A2(n6055), .A3(n6054), .A4(n6053), .ZN(n6062)
         );
  XNOR2_X1 U7076 ( .A(n10614), .B(n6306), .ZN(n6060) );
  XNOR2_X1 U7078 ( .A(n10606), .B(n6307), .ZN(n6059) );
  BUF_X1 U7079 ( .A(data_addr_i[27]), .Z(n10616) );
  XNOR2_X1 U7080 ( .A(n10616), .B(n6318), .ZN(n6058) );
  XNOR2_X1 U7082 ( .A(n10635), .B(n6319), .ZN(n6057) );
  NAND4_X1 U7083 ( .A1(n6060), .A2(n6059), .A3(n6058), .A4(n6057), .ZN(n6061)
         );
  NOR2_X1 U7084 ( .A1(n6062), .A2(n6061), .ZN(n6089) );
  INV_X1 U7085 ( .A(n6688), .ZN(n6813) );
  OAI22_X1 U7086 ( .A1(n6093), .A2(n7816), .B1(n10953), .B2(n6094), .ZN(n6063)
         );
  INV_X1 U7087 ( .A(n6063), .ZN(n6067) );
  INV_X1 U7088 ( .A(n8695), .ZN(n11259) );
  INV_X1 U7089 ( .A(n6251), .ZN(n6064) );
  OAI22_X1 U7090 ( .A1(n22), .A2(n6253), .B1(n11259), .B2(n6064), .ZN(n6065)
         );
  AOI21_X1 U7091 ( .B1(n6257), .B2(n12058), .A(n6065), .ZN(n6066) );
  OAI211_X1 U7092 ( .C1(n6095), .C2(n10486), .A(n6067), .B(n6066), .ZN(n6070)
         );
  OAI22_X1 U7093 ( .A1(n6068), .A2(data_addr_o_11_), .B1(n6649), .B2(n6102), 
        .ZN(n6069) );
  OAI22_X1 U7095 ( .A1(n6090), .A2(data_addr_o_12_), .B1(data_addr_o_9_), .B2(
        n6104), .ZN(n6072) );
  INV_X1 U7096 ( .A(n7820), .ZN(n11343) );
  OAI22_X1 U7097 ( .A1(n11343), .A2(n6105), .B1(n10281), .B2(n6106), .ZN(n6071) );
  NOR2_X1 U7098 ( .A1(n6072), .A2(n6071), .ZN(n6073) );
  XNOR2_X1 U7101 ( .A(n11303), .B(n6075), .ZN(n6076) );
  NOR2_X1 U7102 ( .A1(n6077), .A2(n6076), .ZN(n6088) );
  BUF_X1 U7103 ( .A(data_addr_i[21]), .Z(n10612) );
  XNOR2_X1 U7104 ( .A(n10612), .B(n6078), .ZN(n6081) );
  BUF_X1 U7105 ( .A(data_addr_i[22]), .Z(n10638) );
  XNOR2_X1 U7106 ( .A(n10638), .B(n6079), .ZN(n6080) );
  NOR2_X1 U7107 ( .A1(n6081), .A2(n6080), .ZN(n6087) );
  XNOR2_X1 U7108 ( .A(n10898), .B(n6082), .ZN(n6085) );
  BUF_X1 U7109 ( .A(data_addr_i[24]), .Z(n10629) );
  XNOR2_X1 U7110 ( .A(n10629), .B(n6083), .ZN(n6084) );
  NOR2_X1 U7111 ( .A1(n6085), .A2(n6084), .ZN(n6086) );
  NAND2_X1 U7113 ( .A1(data_addr_o_12_), .A2(n6090), .ZN(n11179) );
  OAI21_X1 U7114 ( .B1(n7324), .B2(n6240), .A(n11179), .ZN(n11191) );
  XNOR2_X1 U7115 ( .A(n9066), .B(n6244), .ZN(n6092) );
  XNOR2_X1 U7116 ( .A(n11309), .B(n6234), .ZN(n6091) );
  NAND2_X1 U7117 ( .A1(n6092), .A2(n6091), .ZN(n6100) );
  INV_X1 U7118 ( .A(data_addr_i[7]), .ZN(n7152) );
  NAND2_X1 U7119 ( .A1(n10493), .A2(n6093), .ZN(n11149) );
  NAND2_X1 U7120 ( .A1(n11331), .A2(n6094), .ZN(n11164) );
  NAND2_X1 U7121 ( .A1(data_addr_o_5_), .A2(n6095), .ZN(n11166) );
  NAND2_X1 U7122 ( .A1(n22), .A2(n6253), .ZN(n11152) );
  OAI211_X1 U7123 ( .C1(n6251), .C2(n10651), .A(n11152), .B(n6096), .ZN(n6097)
         );
  AND2_X1 U7124 ( .A1(data_addr_o_4_), .A2(n6258), .ZN(n11150) );
  NOR2_X1 U7125 ( .A1(n6097), .A2(n11150), .ZN(n6098) );
  NAND4_X1 U7126 ( .A1(n11149), .A2(n11164), .A3(n11166), .A4(n6098), .ZN(
        n6099) );
  NOR3_X1 U7127 ( .A1(n11191), .A2(n6100), .A3(n6099), .ZN(n6111) );
  XNOR2_X1 U7129 ( .A(n9987), .B(n11196), .ZN(n6110) );
  BUF_X1 U7130 ( .A(data_addr_i[31]), .Z(n12123) );
  XNOR2_X1 U7131 ( .A(n12123), .B(n6325), .ZN(n6109) );
  AND2_X1 U7132 ( .A1(data_addr_o_17_), .A2(n6101), .ZN(n11199) );
  NAND2_X1 U7133 ( .A1(n6649), .A2(n6102), .ZN(n11175) );
  NAND2_X1 U7134 ( .A1(data_addr_o_9_), .A2(n6104), .ZN(n11174) );
  NAND2_X1 U7135 ( .A1(n10838), .A2(n6105), .ZN(n11171) );
  NAND2_X1 U7136 ( .A1(n10836), .A2(n6106), .ZN(n11178) );
  NAND4_X1 U7137 ( .A1(n11175), .A2(n11174), .A3(n11171), .A4(n11178), .ZN(
        n6107) );
  NOR2_X1 U7138 ( .A1(n11199), .A2(n6107), .ZN(n6108) );
  NAND4_X1 U7139 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n6379)
         );
  INV_X1 U7140 ( .A(n8089), .ZN(n11004) );
  NOR2_X1 U7141 ( .A1(n7990), .A2(pmp_addr_i[78]), .ZN(n6163) );
  INV_X1 U7142 ( .A(n9941), .ZN(n11227) );
  NOR2_X1 U7143 ( .A1(n10338), .A2(pmp_addr_i[77]), .ZN(n6112) );
  NOR2_X1 U7144 ( .A1(n6163), .A2(n6112), .ZN(n6114) );
  NOR2_X1 U7145 ( .A1(n10403), .A2(pmp_addr_i[80]), .ZN(n6166) );
  NOR2_X1 U7146 ( .A1(n8757), .A2(pmp_addr_i[79]), .ZN(n6113) );
  NOR2_X1 U7147 ( .A1(n6166), .A2(n6113), .ZN(n6168) );
  NAND2_X1 U7148 ( .A1(n6114), .A2(n6168), .ZN(n6172) );
  INV_X1 U7149 ( .A(data_addr_i[11]), .ZN(n9508) );
  NOR2_X1 U7150 ( .A1(n9508), .A2(pmp_addr_i[73]), .ZN(n6115) );
  NOR2_X1 U7151 ( .A1(n10005), .A2(pmp_addr_i[74]), .ZN(n6153) );
  NOR2_X1 U7152 ( .A1(n6115), .A2(n6153), .ZN(n6117) );
  NOR2_X1 U7153 ( .A1(n10342), .A2(pmp_addr_i[75]), .ZN(n6116) );
  INV_X1 U7154 ( .A(data_addr_o_14_), .ZN(n6154) );
  NOR2_X1 U7155 ( .A1(n6154), .A2(pmp_addr_i[76]), .ZN(n6157) );
  NOR2_X1 U7156 ( .A1(n6116), .A2(n6157), .ZN(n6160) );
  NAND2_X1 U7157 ( .A1(n6117), .A2(n6160), .ZN(n6118) );
  NOR2_X1 U7158 ( .A1(n6172), .A2(n6118), .ZN(n6175) );
  INV_X1 U7159 ( .A(data_addr_i[5]), .ZN(n6127) );
  NOR2_X1 U7160 ( .A1(n6127), .A2(pmp_addr_i[67]), .ZN(n6119) );
  NOR2_X1 U7161 ( .A1(n9363), .A2(pmp_addr_i[68]), .ZN(n6130) );
  NOR2_X1 U7162 ( .A1(n6119), .A2(n6130), .ZN(n6133) );
  OR2_X1 U7163 ( .A1(n10010), .A2(pmp_addr_i[65]), .ZN(n6122) );
  AND2_X1 U7164 ( .A1(n8695), .A2(pmp_addr_i[64]), .ZN(n6121) );
  AND2_X1 U7165 ( .A1(n10010), .A2(pmp_addr_i[65]), .ZN(n6120) );
  AOI21_X1 U7166 ( .B1(n6122), .B2(n6121), .A(n6120), .ZN(n6126) );
  INV_X1 U7167 ( .A(data_addr_o_4_), .ZN(n6123) );
  NOR2_X1 U7168 ( .A1(n6123), .A2(pmp_addr_i[66]), .ZN(n6125) );
  NAND2_X1 U7169 ( .A1(n6123), .A2(pmp_addr_i[66]), .ZN(n6124) );
  OAI21_X1 U7170 ( .B1(n6126), .B2(n6125), .A(n6124), .ZN(n6132) );
  NAND2_X1 U7171 ( .A1(n6127), .A2(pmp_addr_i[67]), .ZN(n6129) );
  NAND2_X1 U7172 ( .A1(n8410), .A2(pmp_addr_i[68]), .ZN(n6128) );
  OAI21_X1 U7173 ( .B1(n6130), .B2(n6129), .A(n6128), .ZN(n6131) );
  AOI21_X1 U7174 ( .B1(n6133), .B2(n6132), .A(n6131), .ZN(n6150) );
  INV_X1 U7175 ( .A(n7814), .ZN(n10494) );
  NOR2_X1 U7176 ( .A1(n29), .A2(pmp_addr_i[70]), .ZN(n6139) );
  NOR2_X1 U7177 ( .A1(n7152), .A2(pmp_addr_i[69]), .ZN(n6134) );
  NOR2_X1 U7178 ( .A1(n6139), .A2(n6134), .ZN(n6136) );
  INV_X1 U7179 ( .A(data_addr_o_9_), .ZN(n6140) );
  NOR2_X1 U7180 ( .A1(n6140), .A2(pmp_addr_i[71]), .ZN(n6135) );
  INV_X1 U7181 ( .A(n8238), .ZN(n6141) );
  NOR2_X1 U7182 ( .A1(n6141), .A2(pmp_addr_i[72]), .ZN(n6144) );
  NOR2_X1 U7183 ( .A1(n6135), .A2(n6144), .ZN(n6147) );
  NAND2_X1 U7184 ( .A1(n6136), .A2(n6147), .ZN(n6149) );
  NAND2_X1 U7185 ( .A1(n7152), .A2(pmp_addr_i[69]), .ZN(n6138) );
  NAND2_X1 U7186 ( .A1(n29), .A2(pmp_addr_i[70]), .ZN(n6137) );
  OAI21_X1 U7187 ( .B1(n6139), .B2(n6138), .A(n6137), .ZN(n6146) );
  NAND2_X1 U7188 ( .A1(n6140), .A2(pmp_addr_i[71]), .ZN(n6143) );
  NAND2_X1 U7189 ( .A1(n6141), .A2(pmp_addr_i[72]), .ZN(n6142) );
  OAI21_X1 U7190 ( .B1(n6144), .B2(n6143), .A(n6142), .ZN(n6145) );
  AOI21_X1 U7191 ( .B1(n6147), .B2(n6146), .A(n6145), .ZN(n6148) );
  OAI21_X1 U7192 ( .B1(n6150), .B2(n6149), .A(n6148), .ZN(n6174) );
  NAND2_X1 U7193 ( .A1(n7324), .A2(pmp_addr_i[73]), .ZN(n6152) );
  NAND2_X1 U7194 ( .A1(n7976), .A2(pmp_addr_i[74]), .ZN(n6151) );
  OAI21_X1 U7195 ( .B1(n6153), .B2(n6152), .A(n6151), .ZN(n6159) );
  NAND2_X1 U7196 ( .A1(n10342), .A2(pmp_addr_i[75]), .ZN(n6156) );
  NAND2_X1 U7197 ( .A1(n6154), .A2(pmp_addr_i[76]), .ZN(n6155) );
  OAI21_X1 U7198 ( .B1(n6157), .B2(n6156), .A(n6155), .ZN(n6158) );
  AOI21_X1 U7199 ( .B1(n6160), .B2(n6159), .A(n6158), .ZN(n6171) );
  NAND2_X1 U7200 ( .A1(n10338), .A2(pmp_addr_i[77]), .ZN(n6162) );
  NAND2_X1 U7201 ( .A1(n10047), .A2(pmp_addr_i[78]), .ZN(n6161) );
  OAI21_X1 U7202 ( .B1(n6163), .B2(n6162), .A(n6161), .ZN(n6169) );
  NAND2_X1 U7203 ( .A1(n8444), .A2(pmp_addr_i[79]), .ZN(n6165) );
  NAND2_X1 U7204 ( .A1(n10060), .A2(pmp_addr_i[80]), .ZN(n6164) );
  OAI21_X1 U7205 ( .B1(n6166), .B2(n6165), .A(n6164), .ZN(n6167) );
  AOI21_X1 U7206 ( .B1(n6169), .B2(n6168), .A(n6167), .ZN(n6170) );
  OAI21_X1 U7207 ( .B1(n6172), .B2(n6171), .A(n6170), .ZN(n6173) );
  AOI21_X1 U7208 ( .B1(n6175), .B2(n6174), .A(n6173), .ZN(n6233) );
  NOR2_X1 U7209 ( .A1(n10064), .A2(pmp_addr_i[85]), .ZN(n6176) );
  NOR2_X1 U7210 ( .A1(n9163), .A2(pmp_addr_i[86]), .ZN(n6201) );
  NOR2_X1 U7211 ( .A1(n6176), .A2(n6201), .ZN(n6178) );
  NOR2_X1 U7212 ( .A1(n10768), .A2(pmp_addr_i[87]), .ZN(n6177) );
  INV_X1 U7213 ( .A(data_addr_i[26]), .ZN(n6202) );
  NOR2_X1 U7214 ( .A1(n6202), .A2(pmp_addr_i[88]), .ZN(n6205) );
  NOR2_X1 U7215 ( .A1(n6177), .A2(n6205), .ZN(n6208) );
  NAND2_X1 U7216 ( .A1(n6178), .A2(n6208), .ZN(n6210) );
  INV_X1 U7217 ( .A(data_addr_i[21]), .ZN(n6192) );
  NOR2_X1 U7218 ( .A1(n6192), .A2(pmp_addr_i[83]), .ZN(n6179) );
  NOR2_X1 U7219 ( .A1(n9156), .A2(pmp_addr_i[84]), .ZN(n6195) );
  NOR2_X1 U7220 ( .A1(n6179), .A2(n6195), .ZN(n6198) );
  NOR2_X1 U7221 ( .A1(n10753), .A2(pmp_addr_i[81]), .ZN(n6180) );
  INV_X1 U7222 ( .A(data_addr_i[20]), .ZN(n6188) );
  NOR2_X1 U7223 ( .A1(n6188), .A2(pmp_addr_i[82]), .ZN(n6191) );
  NOR2_X1 U7224 ( .A1(n6180), .A2(n6191), .ZN(n6181) );
  NAND2_X1 U7225 ( .A1(n6198), .A2(n6181), .ZN(n6182) );
  NOR2_X1 U7226 ( .A1(n6210), .A2(n6182), .ZN(n6187) );
  INV_X1 U7227 ( .A(data_addr_i[27]), .ZN(n6212) );
  NOR2_X1 U7228 ( .A1(n6212), .A2(pmp_addr_i[89]), .ZN(n6183) );
  NOR2_X1 U7229 ( .A1(n8807), .A2(pmp_addr_i[90]), .ZN(n6215) );
  NOR2_X1 U7230 ( .A1(n6183), .A2(n6215), .ZN(n6185) );
  INV_X1 U7231 ( .A(data_addr_o_29_), .ZN(n6216) );
  NOR2_X1 U7232 ( .A1(n6216), .A2(pmp_addr_i[91]), .ZN(n6184) );
  NOR2_X1 U7233 ( .A1(n8814), .A2(pmp_addr_i[92]), .ZN(n6219) );
  NOR2_X1 U7234 ( .A1(n6184), .A2(n6219), .ZN(n6222) );
  NAND2_X1 U7235 ( .A1(n6185), .A2(n6222), .ZN(n6186) );
  NOR2_X1 U7236 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[93]), .ZN(n6226) );
  NOR2_X1 U7237 ( .A1(n6186), .A2(n6226), .ZN(n6229) );
  NAND2_X1 U7238 ( .A1(n6187), .A2(n6229), .ZN(n6232) );
  NAND2_X1 U7239 ( .A1(n10753), .A2(pmp_addr_i[81]), .ZN(n6190) );
  NAND2_X1 U7240 ( .A1(n6188), .A2(pmp_addr_i[82]), .ZN(n6189) );
  OAI21_X1 U7241 ( .B1(n6191), .B2(n6190), .A(n6189), .ZN(n6197) );
  NAND2_X1 U7242 ( .A1(n6192), .A2(pmp_addr_i[83]), .ZN(n6194) );
  NAND2_X1 U7243 ( .A1(n9156), .A2(pmp_addr_i[84]), .ZN(n6193) );
  OAI21_X1 U7244 ( .B1(n6195), .B2(n6194), .A(n6193), .ZN(n6196) );
  AOI21_X1 U7245 ( .B1(n6198), .B2(n6197), .A(n6196), .ZN(n6211) );
  NAND2_X1 U7246 ( .A1(n10064), .A2(pmp_addr_i[85]), .ZN(n6200) );
  NAND2_X1 U7247 ( .A1(n9163), .A2(pmp_addr_i[86]), .ZN(n6199) );
  OAI21_X1 U7248 ( .B1(n6201), .B2(n6200), .A(n6199), .ZN(n6207) );
  NAND2_X1 U7249 ( .A1(n6462), .A2(pmp_addr_i[87]), .ZN(n6204) );
  NAND2_X1 U7250 ( .A1(n6202), .A2(pmp_addr_i[88]), .ZN(n6203) );
  OAI21_X1 U7251 ( .B1(n6205), .B2(n6204), .A(n6203), .ZN(n6206) );
  AOI21_X1 U7252 ( .B1(n6208), .B2(n6207), .A(n6206), .ZN(n6209) );
  OAI21_X1 U7253 ( .B1(n6211), .B2(n6210), .A(n6209), .ZN(n6230) );
  NAND2_X1 U7254 ( .A1(n6212), .A2(pmp_addr_i[89]), .ZN(n6214) );
  NAND2_X1 U7255 ( .A1(n8807), .A2(pmp_addr_i[90]), .ZN(n6213) );
  OAI21_X1 U7256 ( .B1(n6215), .B2(n6214), .A(n6213), .ZN(n6221) );
  NAND2_X1 U7257 ( .A1(n6216), .A2(pmp_addr_i[91]), .ZN(n6218) );
  NAND2_X1 U7258 ( .A1(n8814), .A2(pmp_addr_i[92]), .ZN(n6217) );
  OAI21_X1 U7259 ( .B1(n6219), .B2(n6218), .A(n6217), .ZN(n6220) );
  AOI21_X1 U7260 ( .B1(n6222), .B2(n6221), .A(n6220), .ZN(n6227) );
  NAND2_X1 U7261 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[93]), .ZN(n6223)
         );
  NAND2_X1 U7262 ( .A1(n6223), .A2(n4301), .ZN(n6224) );
  NOR2_X1 U7263 ( .A1(n6224), .A2(pmp_addr_i[95]), .ZN(n6225) );
  OAI21_X1 U7264 ( .B1(n6227), .B2(n6226), .A(n6225), .ZN(n6228) );
  AOI21_X1 U7265 ( .B1(n6230), .B2(n6229), .A(n6228), .ZN(n6231) );
  OAI21_X1 U7266 ( .B1(n6233), .B2(n6232), .A(n6231), .ZN(n6377) );
  INV_X1 U7267 ( .A(n8089), .ZN(n10335) );
  NOR2_X1 U7268 ( .A1(n10335), .A2(n11194), .ZN(n6290) );
  INV_X1 U7269 ( .A(n9941), .ZN(n10657) );
  NOR2_X1 U7270 ( .A1(n10657), .A2(n11187), .ZN(n6235) );
  NOR2_X1 U7271 ( .A1(n6290), .A2(n6235), .ZN(n6239) );
  INV_X2 U7273 ( .A(n10297), .ZN(n10857) );
  NOR2_X1 U7274 ( .A1(n10857), .A2(n1913), .ZN(n6293) );
  NOR2_X1 U7275 ( .A1(n6813), .A2(n6101), .ZN(n6238) );
  NOR2_X1 U7276 ( .A1(n6293), .A2(n6238), .ZN(n6296) );
  NAND2_X1 U7277 ( .A1(n6239), .A2(n6296), .ZN(n6299) );
  INV_X1 U7278 ( .A(n7324), .ZN(n8246) );
  NOR2_X1 U7279 ( .A1(n8246), .A2(n6068), .ZN(n6242) );
  NOR2_X1 U7280 ( .A1(data_addr_o_12_), .A2(n6090), .ZN(n6282) );
  NOR2_X1 U7281 ( .A1(n6242), .A2(n6282), .ZN(n6246) );
  INV_X1 U7282 ( .A(data_addr_i[13]), .ZN(n10466) );
  NOR2_X1 U7284 ( .A1(n10847), .A2(n6102), .ZN(n6245) );
  INV_X1 U7285 ( .A(data_addr_i[14]), .ZN(n10518) );
  INV_X1 U7286 ( .A(n10518), .ZN(n10848) );
  NOR2_X1 U7287 ( .A1(n10848), .A2(n11184), .ZN(n6284) );
  NOR2_X1 U7288 ( .A1(n6245), .A2(n6284), .ZN(n6287) );
  NAND2_X1 U7289 ( .A1(n6246), .A2(n6287), .ZN(n6247) );
  NOR2_X1 U7290 ( .A1(n6299), .A2(n6247), .ZN(n6302) );
  NOR2_X1 U7291 ( .A1(n10486), .A2(n6095), .ZN(n6250) );
  NOR2_X1 U7292 ( .A1(data_addr_o_6_), .A2(n6094), .ZN(n6262) );
  NOR2_X1 U7293 ( .A1(n6250), .A2(n6262), .ZN(n6265) );
  INV_X1 U7294 ( .A(n10651), .ZN(data_addr_o_2_) );
  OR2_X1 U7295 ( .A1(data_addr_o_2_), .A2(n6064), .ZN(n6256) );
  INV_X1 U7296 ( .A(n6252), .ZN(n6253) );
  OR2_X1 U7297 ( .A1(n22), .A2(n6253), .ZN(n6255) );
  AND2_X1 U7298 ( .A1(n22), .A2(n6253), .ZN(n6254) );
  AOI21_X1 U7299 ( .B1(n6256), .B2(n6255), .A(n6254), .ZN(n6261) );
  INV_X1 U7300 ( .A(n6257), .ZN(n6258) );
  NOR2_X1 U7301 ( .A1(n10479), .A2(n6258), .ZN(n6260) );
  NAND2_X1 U7302 ( .A1(n10479), .A2(n6258), .ZN(n6259) );
  OAI21_X1 U7303 ( .B1(n6261), .B2(n6260), .A(n6259), .ZN(n6264) );
  OAI21_X1 U7304 ( .B1(n6262), .B2(n11166), .A(n11164), .ZN(n6263) );
  AOI21_X1 U7305 ( .B1(n6265), .B2(n6264), .A(n6263), .ZN(n6280) );
  INV_X1 U7306 ( .A(data_addr_i[9]), .ZN(n10501) );
  INV_X1 U7307 ( .A(n10501), .ZN(n8237) );
  NOR2_X1 U7308 ( .A1(n8237), .A2(n6104), .ZN(n6268) );
  INV_X1 U7309 ( .A(n7820), .ZN(n8238) );
  NOR2_X1 U7310 ( .A1(n8238), .A2(n6105), .ZN(n6274) );
  NOR2_X1 U7311 ( .A1(n6268), .A2(n6274), .ZN(n6277) );
  NOR2_X1 U7312 ( .A1(n10836), .A2(n6106), .ZN(n6273) );
  INV_X1 U7313 ( .A(n7152), .ZN(data_addr_o_7_) );
  NOR2_X1 U7314 ( .A1(data_addr_o_7_), .A2(n6093), .ZN(n6271) );
  NOR2_X1 U7315 ( .A1(n6273), .A2(n6271), .ZN(n6272) );
  NAND2_X1 U7316 ( .A1(n6277), .A2(n6272), .ZN(n6279) );
  OAI21_X1 U7317 ( .B1(n6273), .B2(n11149), .A(n11178), .ZN(n6276) );
  OAI21_X1 U7318 ( .B1(n6274), .B2(n11174), .A(n11171), .ZN(n6275) );
  AOI21_X1 U7319 ( .B1(n6277), .B2(n6276), .A(n6275), .ZN(n6278) );
  OAI21_X1 U7320 ( .B1(n6280), .B2(n6279), .A(n6278), .ZN(n6301) );
  NAND2_X1 U7321 ( .A1(n8246), .A2(n6068), .ZN(n6281) );
  OAI21_X1 U7322 ( .B1(n6282), .B2(n6281), .A(n11179), .ZN(n6286) );
  NAND2_X1 U7323 ( .A1(n10848), .A2(n11184), .ZN(n6283) );
  OAI21_X1 U7324 ( .B1(n6284), .B2(n11175), .A(n6283), .ZN(n6285) );
  AOI21_X1 U7325 ( .B1(n6287), .B2(n6286), .A(n6285), .ZN(n6298) );
  NAND2_X1 U7326 ( .A1(n10657), .A2(n11187), .ZN(n6289) );
  NAND2_X1 U7327 ( .A1(n10335), .A2(n11194), .ZN(n6288) );
  OAI21_X1 U7328 ( .B1(n6290), .B2(n6289), .A(n6288), .ZN(n6295) );
  NAND2_X1 U7329 ( .A1(n6813), .A2(n6101), .ZN(n6292) );
  NAND2_X1 U7330 ( .A1(n10857), .A2(n1913), .ZN(n6291) );
  OAI21_X1 U7331 ( .B1(n6293), .B2(n6292), .A(n6291), .ZN(n6294) );
  AOI21_X1 U7332 ( .B1(n6296), .B2(n6295), .A(n6294), .ZN(n6297) );
  OAI21_X1 U7333 ( .B1(n6299), .B2(n6298), .A(n6297), .ZN(n6300) );
  AOI21_X1 U7334 ( .B1(n6302), .B2(n6301), .A(n6300), .ZN(n6374) );
  NOR2_X1 U7335 ( .A1(n10898), .A2(n6082), .ZN(n6305) );
  BUF_X1 U7336 ( .A(data_addr_i[24]), .Z(n10899) );
  NOR2_X1 U7337 ( .A1(n10899), .A2(n6083), .ZN(n6342) );
  NOR2_X1 U7338 ( .A1(n6305), .A2(n6342), .ZN(n6309) );
  BUF_X1 U7339 ( .A(data_addr_i[25]), .Z(n9923) );
  INV_X1 U7340 ( .A(n6306), .ZN(n6343) );
  NOR2_X1 U7341 ( .A1(n9923), .A2(n6343), .ZN(n6308) );
  INV_X1 U7342 ( .A(n6307), .ZN(n6344) );
  NOR2_X1 U7343 ( .A1(n10606), .A2(n6344), .ZN(n6347) );
  NOR2_X1 U7344 ( .A1(n6308), .A2(n6347), .ZN(n6350) );
  NAND2_X1 U7345 ( .A1(n6309), .A2(n6350), .ZN(n6352) );
  BUF_X1 U7346 ( .A(data_addr_i[21]), .Z(n10891) );
  NOR2_X1 U7347 ( .A1(n10891), .A2(n6078), .ZN(n6312) );
  NOR2_X1 U7348 ( .A1(n9529), .A2(n6079), .ZN(n6336) );
  NOR2_X1 U7349 ( .A1(n6312), .A2(n6336), .ZN(n6339) );
  BUF_X1 U7350 ( .A(data_addr_i[19]), .Z(n10886) );
  INV_X1 U7351 ( .A(n6313), .ZN(n6330) );
  NOR2_X1 U7352 ( .A1(n10886), .A2(n6330), .ZN(n6315) );
  NOR2_X1 U7354 ( .A1(n10530), .A2(n1977), .ZN(n6333) );
  NOR2_X1 U7355 ( .A1(n6315), .A2(n6333), .ZN(n6316) );
  NAND2_X1 U7356 ( .A1(n6339), .A2(n6316), .ZN(n6317) );
  NOR2_X1 U7357 ( .A1(n6352), .A2(n6317), .ZN(n6329) );
  NOR2_X1 U7358 ( .A1(n11322), .A2(n2006), .ZN(n6320) );
  BUF_X1 U7359 ( .A(data_addr_i[28]), .Z(n10914) );
  NOR2_X1 U7360 ( .A1(n10914), .A2(n1985), .ZN(n6356) );
  NOR2_X1 U7361 ( .A1(n6320), .A2(n6356), .ZN(n6324) );
  BUF_X1 U7362 ( .A(data_addr_i[29]), .Z(n10918) );
  NOR2_X1 U7363 ( .A1(n10918), .A2(n6075), .ZN(n6323) );
  NOR2_X1 U7365 ( .A1(n10919), .A2(n1981), .ZN(n6359) );
  NOR2_X1 U7366 ( .A1(n6323), .A2(n6359), .ZN(n6362) );
  NAND2_X1 U7367 ( .A1(n6324), .A2(n6362), .ZN(n6328) );
  INV_X1 U7368 ( .A(n9634), .ZN(n9549) );
  NOR2_X1 U7369 ( .A1(n10662), .A2(n5632), .ZN(n6326) );
  NOR2_X1 U7370 ( .A1(n6326), .A2(pmp_addr_i[62]), .ZN(n6327) );
  INV_X1 U7371 ( .A(pmp_addr_i[63]), .ZN(n6364) );
  NAND2_X1 U7372 ( .A1(n6327), .A2(n6364), .ZN(n6367) );
  NOR2_X1 U7373 ( .A1(n6328), .A2(n6367), .ZN(n6370) );
  NAND2_X1 U7374 ( .A1(n6329), .A2(n6370), .ZN(n6373) );
  NAND2_X1 U7375 ( .A1(n10886), .A2(n6330), .ZN(n6332) );
  NAND2_X1 U7376 ( .A1(n10530), .A2(n1977), .ZN(n6331) );
  OAI21_X1 U7377 ( .B1(n6333), .B2(n6332), .A(n6331), .ZN(n6338) );
  NAND2_X1 U7378 ( .A1(n10891), .A2(n6078), .ZN(n6335) );
  NAND2_X1 U7379 ( .A1(n9915), .A2(n6079), .ZN(n6334) );
  OAI21_X1 U7380 ( .B1(n6336), .B2(n6335), .A(n6334), .ZN(n6337) );
  AOI21_X1 U7381 ( .B1(n6339), .B2(n6338), .A(n6337), .ZN(n6353) );
  NAND2_X1 U7382 ( .A1(n10898), .A2(n6082), .ZN(n6341) );
  NAND2_X1 U7383 ( .A1(n10899), .A2(n6083), .ZN(n6340) );
  OAI21_X1 U7384 ( .B1(n6342), .B2(n6341), .A(n6340), .ZN(n6349) );
  NAND2_X1 U7385 ( .A1(n9923), .A2(n6343), .ZN(n6346) );
  NAND2_X1 U7386 ( .A1(n10606), .A2(n6344), .ZN(n6345) );
  OAI21_X1 U7387 ( .B1(n6347), .B2(n6346), .A(n6345), .ZN(n6348) );
  AOI21_X1 U7388 ( .B1(n6350), .B2(n6349), .A(n6348), .ZN(n6351) );
  OAI21_X1 U7389 ( .B1(n6353), .B2(n6352), .A(n6351), .ZN(n6371) );
  NAND2_X1 U7390 ( .A1(n11322), .A2(n2006), .ZN(n6355) );
  NAND2_X1 U7391 ( .A1(n10914), .A2(n1985), .ZN(n6354) );
  OAI21_X1 U7392 ( .B1(n6356), .B2(n6355), .A(n6354), .ZN(n6361) );
  NAND2_X1 U7393 ( .A1(n10918), .A2(n6075), .ZN(n6358) );
  NAND2_X1 U7394 ( .A1(n10919), .A2(n1981), .ZN(n6357) );
  OAI21_X1 U7395 ( .B1(n6359), .B2(n6358), .A(n6357), .ZN(n6360) );
  AOI21_X1 U7396 ( .B1(n6362), .B2(n6361), .A(n6360), .ZN(n6368) );
  NAND2_X1 U7397 ( .A1(n12123), .A2(n5632), .ZN(n6363) );
  NOR2_X1 U7398 ( .A1(n6363), .A2(pmp_addr_i[62]), .ZN(n6365) );
  NAND2_X1 U7399 ( .A1(n6365), .A2(n6364), .ZN(n6366) );
  OAI21_X1 U7400 ( .B1(n6368), .B2(n6367), .A(n6366), .ZN(n6369) );
  AOI21_X1 U7401 ( .B1(n6371), .B2(n6370), .A(n6369), .ZN(n6372) );
  OAI21_X1 U7402 ( .B1(n6374), .B2(n6373), .A(n6372), .ZN(n6375) );
  NAND3_X1 U7403 ( .A1(n6377), .A2(n6376), .A3(n6375), .ZN(n6378) );
  OAI21_X1 U7404 ( .B1(n11147), .B2(n6379), .A(n6378), .ZN(n6698) );
  NOR2_X1 U7405 ( .A1(n10047), .A2(pmp_addr_i[494]), .ZN(n6380) );
  NOR2_X1 U7407 ( .A1(pmp_addr_i[495]), .A2(n8444), .ZN(n6427) );
  NOR2_X1 U7408 ( .A1(n6380), .A2(n6427), .ZN(n6430) );
  NOR2_X1 U7409 ( .A1(pmp_addr_i[492]), .A2(n11334), .ZN(n6381) );
  NOR2_X1 U7410 ( .A1(pmp_addr_i[493]), .A2(n10338), .ZN(n6424) );
  NOR2_X1 U7411 ( .A1(n6381), .A2(n6424), .ZN(n6382) );
  NAND2_X1 U7412 ( .A1(n6430), .A2(n6382), .ZN(n6432) );
  NOR2_X1 U7413 ( .A1(pmp_addr_i[488]), .A2(n10701), .ZN(n6383) );
  NOR2_X1 U7414 ( .A1(pmp_addr_i[489]), .A2(n7324), .ZN(n6415) );
  NOR2_X1 U7415 ( .A1(n6383), .A2(n6415), .ZN(n6385) );
  NOR2_X1 U7416 ( .A1(pmp_addr_i[490]), .A2(n10005), .ZN(n6384) );
  INV_X1 U7417 ( .A(data_addr_i[13]), .ZN(n10342) );
  NOR2_X1 U7418 ( .A1(pmp_addr_i[491]), .A2(n10342), .ZN(n6418) );
  NOR2_X1 U7419 ( .A1(n6384), .A2(n6418), .ZN(n6421) );
  NAND2_X1 U7420 ( .A1(n6385), .A2(n6421), .ZN(n6386) );
  NOR2_X1 U7421 ( .A1(n6432), .A2(n6386), .ZN(n6436) );
  INV_X1 U7422 ( .A(n10135), .ZN(n10351) );
  NOR2_X1 U7423 ( .A1(pmp_addr_i[482]), .A2(n10351), .ZN(n6387) );
  INV_X1 U7424 ( .A(data_addr_i[5]), .ZN(n10346) );
  NOR2_X1 U7425 ( .A1(pmp_addr_i[483]), .A2(n10346), .ZN(n6393) );
  NOR2_X1 U7426 ( .A1(n6387), .A2(n6393), .ZN(n6396) );
  INV_X1 U7427 ( .A(data_addr_o_3_), .ZN(n10010) );
  NOR2_X1 U7428 ( .A1(pmp_addr_i[481]), .A2(n10010), .ZN(n6390) );
  NAND2_X1 U7429 ( .A1(pmp_addr_i[480]), .A2(n10651), .ZN(n6389) );
  NAND2_X1 U7430 ( .A1(pmp_addr_i[481]), .A2(n10010), .ZN(n6388) );
  OAI21_X1 U7431 ( .B1(n6390), .B2(n6389), .A(n6388), .ZN(n6395) );
  NAND2_X1 U7432 ( .A1(pmp_addr_i[482]), .A2(n10351), .ZN(n6392) );
  NAND2_X1 U7433 ( .A1(pmp_addr_i[483]), .A2(n10346), .ZN(n6391) );
  OAI21_X1 U7434 ( .B1(n6393), .B2(n6392), .A(n6391), .ZN(n6394) );
  AOI21_X1 U7435 ( .B1(n6396), .B2(n6395), .A(n6394), .ZN(n6412) );
  NOR2_X1 U7436 ( .A1(pmp_addr_i[484]), .A2(n9363), .ZN(n6397) );
  INV_X1 U7437 ( .A(n7816), .ZN(n6400) );
  NOR2_X1 U7438 ( .A1(pmp_addr_i[485]), .A2(n6400), .ZN(n6403) );
  NOR2_X1 U7439 ( .A1(n6397), .A2(n6403), .ZN(n6399) );
  NOR2_X1 U7440 ( .A1(pmp_addr_i[486]), .A2(n29), .ZN(n6398) );
  NOR2_X1 U7441 ( .A1(pmp_addr_i[487]), .A2(n6140), .ZN(n6406) );
  NOR2_X1 U7442 ( .A1(n6398), .A2(n6406), .ZN(n6409) );
  NAND2_X1 U7443 ( .A1(n6399), .A2(n6409), .ZN(n6411) );
  NAND2_X1 U7444 ( .A1(pmp_addr_i[484]), .A2(n10362), .ZN(n6402) );
  NAND2_X1 U7445 ( .A1(pmp_addr_i[485]), .A2(n6400), .ZN(n6401) );
  OAI21_X1 U7446 ( .B1(n6403), .B2(n6402), .A(n6401), .ZN(n6408) );
  NAND2_X1 U7447 ( .A1(pmp_addr_i[486]), .A2(n29), .ZN(n6405) );
  NAND2_X1 U7448 ( .A1(pmp_addr_i[487]), .A2(n6140), .ZN(n6404) );
  OAI21_X1 U7449 ( .B1(n6406), .B2(n6405), .A(n6404), .ZN(n6407) );
  AOI21_X1 U7450 ( .B1(n6409), .B2(n6408), .A(n6407), .ZN(n6410) );
  OAI21_X1 U7451 ( .B1(n6412), .B2(n6411), .A(n6410), .ZN(n6435) );
  NAND2_X1 U7452 ( .A1(pmp_addr_i[488]), .A2(n6141), .ZN(n6414) );
  NAND2_X1 U7453 ( .A1(pmp_addr_i[489]), .A2(n10711), .ZN(n6413) );
  OAI21_X1 U7454 ( .B1(n6415), .B2(n6414), .A(n6413), .ZN(n6420) );
  NAND2_X1 U7455 ( .A1(pmp_addr_i[490]), .A2(n7976), .ZN(n6417) );
  NAND2_X1 U7456 ( .A1(pmp_addr_i[491]), .A2(n10342), .ZN(n6416) );
  OAI21_X1 U7457 ( .B1(n6418), .B2(n6417), .A(n6416), .ZN(n6419) );
  AOI21_X1 U7458 ( .B1(n6421), .B2(n6420), .A(n6419), .ZN(n6433) );
  NAND2_X1 U7459 ( .A1(pmp_addr_i[492]), .A2(n10000), .ZN(n6423) );
  NAND2_X1 U7460 ( .A1(pmp_addr_i[493]), .A2(n10338), .ZN(n6422) );
  OAI21_X1 U7461 ( .B1(n6424), .B2(n6423), .A(n6422), .ZN(n6429) );
  NAND2_X1 U7462 ( .A1(n7057), .A2(pmp_addr_i[494]), .ZN(n6426) );
  NAND2_X1 U7463 ( .A1(pmp_addr_i[495]), .A2(n7995), .ZN(n6425) );
  OAI21_X1 U7464 ( .B1(n6427), .B2(n6426), .A(n6425), .ZN(n6428) );
  AOI21_X1 U7465 ( .B1(n6430), .B2(n6429), .A(n6428), .ZN(n6431) );
  OAI21_X1 U7466 ( .B1(n6433), .B2(n6432), .A(n6431), .ZN(n6434) );
  AOI21_X1 U7467 ( .B1(n6436), .B2(n6435), .A(n6434), .ZN(n6495) );
  INV_X1 U7468 ( .A(n12260), .ZN(n10403) );
  NOR2_X1 U7469 ( .A1(pmp_addr_i[496]), .A2(n10403), .ZN(n6437) );
  NOR2_X1 U7470 ( .A1(pmp_addr_i[497]), .A2(n10414), .ZN(n6452) );
  NOR2_X1 U7471 ( .A1(n6437), .A2(n6452), .ZN(n6439) );
  NOR2_X1 U7472 ( .A1(pmp_addr_i[498]), .A2(n6188), .ZN(n6438) );
  NOR2_X1 U7473 ( .A1(pmp_addr_i[499]), .A2(n6192), .ZN(n6455) );
  NOR2_X1 U7474 ( .A1(n6438), .A2(n6455), .ZN(n6458) );
  NAND2_X1 U7475 ( .A1(n6439), .A2(n6458), .ZN(n6443) );
  NOR2_X1 U7476 ( .A1(pmp_addr_i[500]), .A2(n9425), .ZN(n6440) );
  NOR2_X1 U7477 ( .A1(pmp_addr_i[501]), .A2(n10064), .ZN(n6461) );
  NOR2_X1 U7478 ( .A1(n6440), .A2(n6461), .ZN(n6442) );
  NOR2_X1 U7479 ( .A1(pmp_addr_i[502]), .A2(n10428), .ZN(n6441) );
  INV_X1 U7480 ( .A(n10614), .ZN(n6462) );
  NOR2_X1 U7481 ( .A1(pmp_addr_i[503]), .A2(n6462), .ZN(n6465) );
  NOR2_X1 U7482 ( .A1(n6441), .A2(n6465), .ZN(n6468) );
  NAND2_X1 U7483 ( .A1(n6442), .A2(n6468), .ZN(n6470) );
  NOR2_X1 U7484 ( .A1(n6443), .A2(n6470), .ZN(n6449) );
  NOR2_X1 U7485 ( .A1(pmp_addr_i[504]), .A2(n10439), .ZN(n6444) );
  NOR2_X1 U7486 ( .A1(pmp_addr_i[505]), .A2(n9438), .ZN(n6474) );
  NOR2_X1 U7487 ( .A1(n6444), .A2(n6474), .ZN(n6446) );
  INV_X1 U7488 ( .A(data_addr_o_29_), .ZN(n10100) );
  NOR2_X1 U7489 ( .A1(pmp_addr_i[507]), .A2(n10100), .ZN(n6477) );
  NOR2_X1 U7490 ( .A1(pmp_addr_i[506]), .A2(n8807), .ZN(n6445) );
  NOR2_X1 U7491 ( .A1(n6477), .A2(n6445), .ZN(n6480) );
  NAND2_X1 U7492 ( .A1(n6446), .A2(n6480), .ZN(n6448) );
  INV_X1 U7493 ( .A(n9549), .ZN(n10107) );
  NOR2_X1 U7494 ( .A1(pmp_addr_i[509]), .A2(n10107), .ZN(n6483) );
  NOR2_X1 U7495 ( .A1(pmp_addr_i[508]), .A2(n8814), .ZN(n6447) );
  OR2_X1 U7496 ( .A1(n6483), .A2(n6447), .ZN(n6488) );
  NOR2_X1 U7497 ( .A1(n6448), .A2(n6488), .ZN(n6491) );
  NAND2_X1 U7498 ( .A1(n6449), .A2(n6491), .ZN(n6494) );
  INV_X1 U7499 ( .A(n12260), .ZN(n10060) );
  NAND2_X1 U7500 ( .A1(pmp_addr_i[496]), .A2(n10060), .ZN(n6451) );
  NAND2_X1 U7501 ( .A1(pmp_addr_i[497]), .A2(n9414), .ZN(n6450) );
  OAI21_X1 U7502 ( .B1(n6452), .B2(n6451), .A(n6450), .ZN(n6457) );
  NAND2_X1 U7503 ( .A1(pmp_addr_i[498]), .A2(n10754), .ZN(n6454) );
  NAND2_X1 U7504 ( .A1(pmp_addr_i[499]), .A2(n9418), .ZN(n6453) );
  OAI21_X1 U7505 ( .B1(n6455), .B2(n6454), .A(n6453), .ZN(n6456) );
  AOI21_X1 U7506 ( .B1(n6458), .B2(n6457), .A(n6456), .ZN(n6471) );
  NAND2_X1 U7507 ( .A1(pmp_addr_i[500]), .A2(n9156), .ZN(n6460) );
  NAND2_X1 U7508 ( .A1(pmp_addr_i[501]), .A2(n10064), .ZN(n6459) );
  OAI21_X1 U7509 ( .B1(n6461), .B2(n6460), .A(n6459), .ZN(n6467) );
  NAND2_X1 U7510 ( .A1(pmp_addr_i[502]), .A2(n10428), .ZN(n6464) );
  NAND2_X1 U7511 ( .A1(pmp_addr_i[503]), .A2(n6462), .ZN(n6463) );
  OAI21_X1 U7512 ( .B1(n6465), .B2(n6464), .A(n6463), .ZN(n6466) );
  AOI21_X1 U7513 ( .B1(n6468), .B2(n6467), .A(n6466), .ZN(n6469) );
  OAI21_X1 U7514 ( .B1(n6471), .B2(n6470), .A(n6469), .ZN(n6492) );
  NAND2_X1 U7515 ( .A1(pmp_addr_i[504]), .A2(n6202), .ZN(n6473) );
  NAND2_X1 U7516 ( .A1(pmp_addr_i[505]), .A2(n10096), .ZN(n6472) );
  OAI21_X1 U7517 ( .B1(n6474), .B2(n6473), .A(n6472), .ZN(n6479) );
  NAND2_X1 U7518 ( .A1(pmp_addr_i[506]), .A2(n8807), .ZN(n6476) );
  NAND2_X1 U7519 ( .A1(pmp_addr_i[507]), .A2(n10100), .ZN(n6475) );
  OAI21_X1 U7520 ( .B1(n6477), .B2(n6476), .A(n6475), .ZN(n6478) );
  AOI21_X1 U7521 ( .B1(n6480), .B2(n6479), .A(n6478), .ZN(n6489) );
  NAND2_X1 U7522 ( .A1(pmp_addr_i[508]), .A2(n8494), .ZN(n6482) );
  NAND2_X1 U7523 ( .A1(pmp_addr_i[509]), .A2(data_addr_o_31__BAR), .ZN(n6481)
         );
  OAI21_X1 U7524 ( .B1(n6483), .B2(n6482), .A(n6481), .ZN(n6486) );
  INV_X1 U7525 ( .A(n6484), .ZN(n6485) );
  NOR2_X1 U7526 ( .A1(n6486), .A2(n6485), .ZN(n6487) );
  OAI21_X1 U7527 ( .B1(n6489), .B2(n6488), .A(n6487), .ZN(n6490) );
  AOI21_X1 U7528 ( .B1(n6492), .B2(n6491), .A(n6490), .ZN(n6493) );
  OAI21_X1 U7529 ( .B1(n6495), .B2(n6494), .A(n6493), .ZN(n6625) );
  BUF_X1 U7530 ( .A(data_addr_o_20_), .Z(n10887) );
  NOR2_X1 U7531 ( .A1(n4013), .A2(n10887), .ZN(n6496) );
  INV_X1 U7532 ( .A(n6626), .ZN(n6565) );
  BUF_X1 U7533 ( .A(data_addr_i[21]), .Z(n10202) );
  NOR2_X1 U7534 ( .A1(n6565), .A2(n10202), .ZN(n6568) );
  NOR2_X1 U7535 ( .A1(n6496), .A2(n6568), .ZN(n6498) );
  INV_X1 U7536 ( .A(n6627), .ZN(n6569) );
  NOR2_X1 U7537 ( .A1(n6569), .A2(n9915), .ZN(n6497) );
  INV_X1 U7538 ( .A(n6628), .ZN(n6570) );
  NOR2_X1 U7539 ( .A1(n6570), .A2(n10737), .ZN(n6573) );
  NOR2_X1 U7540 ( .A1(n6497), .A2(n6573), .ZN(n6576) );
  NAND2_X1 U7541 ( .A1(n6498), .A2(n6576), .ZN(n6578) );
  INV_X1 U7542 ( .A(n6648), .ZN(n6557) );
  NOR2_X1 U7543 ( .A1(n6557), .A2(n10857), .ZN(n6499) );
  INV_X1 U7544 ( .A(n6644), .ZN(n6558) );
  NOR2_X1 U7545 ( .A1(n6558), .A2(n10886), .ZN(n6561) );
  NOR2_X1 U7546 ( .A1(n6499), .A2(n6561), .ZN(n6564) );
  NAND2_X1 U7547 ( .A1(n11793), .A2(n6688), .ZN(n11773) );
  INV_X1 U7548 ( .A(n11773), .ZN(n6556) );
  NAND2_X1 U7549 ( .A1(n8089), .A2(n6554), .ZN(n6659) );
  INV_X1 U7550 ( .A(n6659), .ZN(n6500) );
  NOR2_X1 U7551 ( .A1(n6556), .A2(n6500), .ZN(n6501) );
  NAND2_X1 U7552 ( .A1(n6564), .A2(n6501), .ZN(n6502) );
  NOR2_X1 U7553 ( .A1(n6578), .A2(n6502), .ZN(n6582) );
  NOR2_X1 U7554 ( .A1(n11259), .A2(n323), .ZN(n6505) );
  INV_X1 U7555 ( .A(n10473), .ZN(n10958) );
  NOR2_X1 U7556 ( .A1(n10958), .A2(n6677), .ZN(n6504) );
  NAND2_X1 U7557 ( .A1(n10958), .A2(n6677), .ZN(n11798) );
  OAI21_X1 U7558 ( .B1(n6505), .B2(n6504), .A(n11798), .ZN(n6508) );
  NAND2_X1 U7559 ( .A1(n12058), .A2(n6506), .ZN(n6680) );
  INV_X1 U7560 ( .A(n12058), .ZN(n11288) );
  AND2_X1 U7561 ( .A1(n11288), .A2(n6674), .ZN(n6507) );
  AOI21_X1 U7562 ( .B1(n6508), .B2(n6680), .A(n6507), .ZN(n6517) );
  INV_X1 U7563 ( .A(n11291), .ZN(n10824) );
  OR2_X1 U7564 ( .A1(n10824), .A2(n3887), .ZN(n6511) );
  OR2_X1 U7565 ( .A1(n10953), .A2(n3888), .ZN(n6514) );
  NAND2_X1 U7566 ( .A1(n6511), .A2(n6514), .ZN(n6516) );
  AND2_X1 U7567 ( .A1(n10824), .A2(n3887), .ZN(n6513) );
  AND2_X1 U7568 ( .A1(n10953), .A2(n3888), .ZN(n6512) );
  AOI21_X1 U7569 ( .B1(n6514), .B2(n6513), .A(n6512), .ZN(n6515) );
  OAI21_X1 U7570 ( .B1(n6517), .B2(n6516), .A(n6515), .ZN(n6524) );
  INV_X1 U7571 ( .A(n7814), .ZN(n10281) );
  NOR2_X1 U7572 ( .A1(n10281), .A2(n3909), .ZN(n6521) );
  NOR2_X1 U7573 ( .A1(n7816), .A2(n3908), .ZN(n6520) );
  NOR2_X1 U7574 ( .A1(n6521), .A2(n6520), .ZN(n6523) );
  NAND2_X1 U7575 ( .A1(n7816), .A2(n3908), .ZN(n11764) );
  NAND2_X1 U7576 ( .A1(n10281), .A2(n3909), .ZN(n11778) );
  OAI21_X1 U7577 ( .B1(n6521), .B2(n11764), .A(n11778), .ZN(n6522) );
  AOI21_X1 U7578 ( .B1(n6524), .B2(n6523), .A(n6522), .ZN(n6553) );
  OR2_X1 U7579 ( .A1(data_addr_o_9_), .A2(n6654), .ZN(n6526) );
  OR2_X1 U7580 ( .A1(n11343), .A2(n3912), .ZN(n6538) );
  NAND2_X1 U7581 ( .A1(n6526), .A2(n6538), .ZN(n6530) );
  OR2_X1 U7582 ( .A1(data_addr_o_11_), .A2(n3955), .ZN(n6529) );
  OR2_X1 U7583 ( .A1(data_addr_o_12_), .A2(n6683), .ZN(n6541) );
  NAND2_X1 U7584 ( .A1(n6529), .A2(n6541), .ZN(n6543) );
  NOR2_X1 U7585 ( .A1(n6530), .A2(n6543), .ZN(n6535) );
  OR2_X1 U7586 ( .A1(data_addr_o_13_), .A2(n3959), .ZN(n6532) );
  BUF_X1 U7587 ( .A(data_addr_o_14_), .Z(n9066) );
  OR2_X1 U7588 ( .A1(n9066), .A2(n4733), .ZN(n6546) );
  NAND2_X1 U7589 ( .A1(n6532), .A2(n6546), .ZN(n6534) );
  NOR2_X1 U7590 ( .A1(n11309), .A2(n4730), .ZN(n6651) );
  NOR2_X1 U7591 ( .A1(n6534), .A2(n6651), .ZN(n6549) );
  NAND2_X1 U7592 ( .A1(n6535), .A2(n6549), .ZN(n6552) );
  AND2_X1 U7593 ( .A1(data_addr_o_9_), .A2(n6654), .ZN(n6537) );
  AND2_X1 U7594 ( .A1(n11343), .A2(n3912), .ZN(n6536) );
  AOI21_X1 U7595 ( .B1(n6538), .B2(n6537), .A(n6536), .ZN(n6544) );
  AND2_X1 U7596 ( .A1(data_addr_o_11_), .A2(n3955), .ZN(n6540) );
  AND2_X1 U7597 ( .A1(data_addr_o_12_), .A2(n6683), .ZN(n6539) );
  AOI21_X1 U7598 ( .B1(n6541), .B2(n6540), .A(n6539), .ZN(n6542) );
  OAI21_X1 U7599 ( .B1(n6544), .B2(n6543), .A(n6542), .ZN(n6550) );
  AND2_X1 U7600 ( .A1(data_addr_o_13_), .A2(n3959), .ZN(n6545) );
  AND2_X1 U7601 ( .A1(n9066), .A2(n4733), .ZN(n11763) );
  AOI21_X1 U7602 ( .B1(n6546), .B2(n6545), .A(n11763), .ZN(n6547) );
  NAND2_X1 U7603 ( .A1(n11309), .A2(n4730), .ZN(n11806) );
  OAI21_X1 U7604 ( .B1(n6547), .B2(n6651), .A(n11806), .ZN(n6548) );
  AOI21_X1 U7605 ( .B1(n6550), .B2(n6549), .A(n6548), .ZN(n6551) );
  OAI21_X1 U7606 ( .B1(n6553), .B2(n6552), .A(n6551), .ZN(n6581) );
  NAND2_X1 U7607 ( .A1(n9987), .A2(n3965), .ZN(n11809) );
  NAND2_X1 U7608 ( .A1(n4719), .A2(n6813), .ZN(n6555) );
  OAI21_X1 U7609 ( .B1(n6556), .B2(n11809), .A(n6555), .ZN(n6563) );
  NAND2_X1 U7610 ( .A1(n6557), .A2(n10857), .ZN(n6560) );
  NAND2_X1 U7611 ( .A1(n6558), .A2(n11283), .ZN(n6559) );
  OAI21_X1 U7612 ( .B1(n6561), .B2(n6560), .A(n6559), .ZN(n6562) );
  AOI21_X1 U7613 ( .B1(n6564), .B2(n6563), .A(n6562), .ZN(n6579) );
  NAND2_X1 U7614 ( .A1(n4013), .A2(n10887), .ZN(n6567) );
  NAND2_X1 U7615 ( .A1(n6565), .A2(n10202), .ZN(n6566) );
  OAI21_X1 U7616 ( .B1(n6568), .B2(n6567), .A(n6566), .ZN(n6575) );
  NAND2_X1 U7617 ( .A1(n6569), .A2(n9915), .ZN(n6572) );
  NAND2_X1 U7618 ( .A1(n6570), .A2(n10737), .ZN(n6571) );
  OAI21_X1 U7619 ( .B1(n6573), .B2(n6572), .A(n6571), .ZN(n6574) );
  AOI21_X1 U7620 ( .B1(n6576), .B2(n6575), .A(n6574), .ZN(n6577) );
  OAI21_X1 U7621 ( .B1(n6579), .B2(n6578), .A(n6577), .ZN(n6580) );
  AOI21_X1 U7622 ( .B1(n6582), .B2(n6581), .A(n6580), .ZN(n6622) );
  INV_X1 U7623 ( .A(n6629), .ZN(n6591) );
  NOR2_X1 U7624 ( .A1(n6591), .A2(n10899), .ZN(n6583) );
  NOR2_X1 U7625 ( .A1(n4026), .A2(n9923), .ZN(n6594) );
  NOR2_X1 U7626 ( .A1(n6583), .A2(n6594), .ZN(n6585) );
  INV_X1 U7627 ( .A(n6635), .ZN(n6595) );
  BUF_X1 U7628 ( .A(data_addr_i[26]), .Z(n10904) );
  NOR2_X1 U7629 ( .A1(n6595), .A2(n10904), .ZN(n6584) );
  INV_X1 U7630 ( .A(n6663), .ZN(n6596) );
  NOR2_X1 U7631 ( .A1(n6596), .A2(n10746), .ZN(n6599) );
  NOR2_X1 U7632 ( .A1(n6584), .A2(n6599), .ZN(n6602) );
  NAND2_X1 U7633 ( .A1(n6585), .A2(n6602), .ZN(n6589) );
  NOR2_X1 U7634 ( .A1(n4045), .A2(n24), .ZN(n6611) );
  INV_X1 U7635 ( .A(n6637), .ZN(n6608) );
  NOR2_X1 U7636 ( .A1(n6608), .A2(n10919), .ZN(n6586) );
  NOR2_X1 U7637 ( .A1(n6611), .A2(n6586), .ZN(n6614) );
  INV_X1 U7638 ( .A(n6636), .ZN(n6603) );
  NOR2_X1 U7639 ( .A1(n6603), .A2(n10747), .ZN(n6587) );
  INV_X1 U7640 ( .A(n6664), .ZN(n6604) );
  NOR2_X1 U7641 ( .A1(n6604), .A2(n10918), .ZN(n6607) );
  NOR2_X1 U7642 ( .A1(n6587), .A2(n6607), .ZN(n6588) );
  NAND2_X1 U7643 ( .A1(n6614), .A2(n6588), .ZN(n6616) );
  NOR2_X1 U7644 ( .A1(n6589), .A2(n6616), .ZN(n6590) );
  NAND2_X1 U7646 ( .A1(n6590), .A2(n2589), .ZN(n6621) );
  NAND2_X1 U7647 ( .A1(n6591), .A2(n10899), .ZN(n6593) );
  NAND2_X1 U7648 ( .A1(n4026), .A2(n9923), .ZN(n6592) );
  OAI21_X1 U7649 ( .B1(n6594), .B2(n6593), .A(n6592), .ZN(n6601) );
  NAND2_X1 U7650 ( .A1(n6595), .A2(n10904), .ZN(n6598) );
  NAND2_X1 U7651 ( .A1(n6596), .A2(n10746), .ZN(n6597) );
  OAI21_X1 U7652 ( .B1(n6599), .B2(n6598), .A(n6597), .ZN(n6600) );
  AOI21_X1 U7653 ( .B1(n6602), .B2(n6601), .A(n6600), .ZN(n6617) );
  NAND2_X1 U7654 ( .A1(n6603), .A2(n10747), .ZN(n6606) );
  NAND2_X1 U7655 ( .A1(n6604), .A2(n10918), .ZN(n6605) );
  OAI21_X1 U7656 ( .B1(n6607), .B2(n6606), .A(n6605), .ZN(n6613) );
  NAND2_X1 U7657 ( .A1(n6608), .A2(n10919), .ZN(n6610) );
  NAND2_X1 U7658 ( .A1(n4045), .A2(n24), .ZN(n6609) );
  OAI21_X1 U7659 ( .B1(n6611), .B2(n6610), .A(n6609), .ZN(n6612) );
  AOI21_X1 U7660 ( .B1(n6614), .B2(n6613), .A(n6612), .ZN(n6615) );
  OAI21_X1 U7661 ( .B1(n6617), .B2(n6616), .A(n6615), .ZN(n6619) );
  NAND2_X1 U7662 ( .A1(n6619), .A2(n2589), .ZN(n6620) );
  OAI21_X1 U7663 ( .B1(n6622), .B2(n6621), .A(n6620), .ZN(n6623) );
  NAND3_X1 U7664 ( .A1(n6625), .A2(n6624), .A3(n6623), .ZN(n6694) );
  BUF_X1 U7665 ( .A(data_addr_i[21]), .Z(n11312) );
  XNOR2_X1 U7666 ( .A(n6626), .B(n11312), .ZN(n6633) );
  BUF_X1 U7667 ( .A(data_addr_i[22]), .Z(n11313) );
  XNOR2_X1 U7668 ( .A(n6627), .B(n11313), .ZN(n6632) );
  XNOR2_X1 U7670 ( .A(n6628), .B(data_addr_o_23_), .ZN(n6631) );
  XNOR2_X1 U7671 ( .A(n6629), .B(n10629), .ZN(n6630) );
  NAND4_X1 U7672 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .ZN(n6643)
         );
  XNOR2_X1 U7673 ( .A(n6634), .B(n11320), .ZN(n6641) );
  BUF_X1 U7674 ( .A(data_addr_i[26]), .Z(data_addr_o_26_) );
  XNOR2_X1 U7675 ( .A(n6635), .B(data_addr_o_26_), .ZN(n6640) );
  XNOR2_X1 U7677 ( .A(n6636), .B(n10635), .ZN(n6639) );
  XNOR2_X1 U7679 ( .A(n6637), .B(data_addr_o_30_), .ZN(n6638) );
  NAND4_X1 U7680 ( .A1(n6641), .A2(n6640), .A3(n6639), .A4(n6638), .ZN(n6642)
         );
  OR2_X1 U7681 ( .A1(n6643), .A2(n6642), .ZN(n6670) );
  BUF_X1 U7682 ( .A(data_addr_i[19]), .Z(n11283) );
  XNOR2_X1 U7683 ( .A(n6644), .B(n11283), .ZN(n6647) );
  XNOR2_X1 U7685 ( .A(n6645), .B(n9935), .ZN(n6646) );
  AND2_X1 U7686 ( .A1(n6647), .A2(n6646), .ZN(n6668) );
  XNOR2_X1 U7687 ( .A(n6648), .B(n10297), .ZN(n6662) );
  OAI22_X1 U7688 ( .A1(n6683), .A2(data_addr_o_12_), .B1(n6649), .B2(n3959), 
        .ZN(n6650) );
  NOR2_X1 U7689 ( .A1(n6651), .A2(n6650), .ZN(n6660) );
  INV_X1 U7690 ( .A(data_addr_i[14]), .ZN(n11334) );
  OAI22_X1 U7691 ( .A1(n3908), .A2(n7816), .B1(n11331), .B2(n3888), .ZN(n6652)
         );
  AOI21_X1 U7692 ( .B1(n11334), .B2(n6653), .A(n6652), .ZN(n6658) );
  OAI22_X1 U7693 ( .A1(n3912), .A2(n11343), .B1(data_addr_o_11_), .B2(n3955), 
        .ZN(n6656) );
  OAI22_X1 U7694 ( .A1(data_addr_o_9_), .A2(n6654), .B1(n9805), .B2(n3909), 
        .ZN(n6655) );
  NOR2_X1 U7695 ( .A1(n6656), .A2(n6655), .ZN(n6657) );
  NAND4_X1 U7696 ( .A1(n6660), .A2(n6659), .A3(n6658), .A4(n6657), .ZN(n6661)
         );
  NOR2_X1 U7697 ( .A1(n6662), .A2(n6661), .ZN(n6667) );
  BUF_X1 U7698 ( .A(data_addr_i[27]), .Z(n11322) );
  XNOR2_X1 U7699 ( .A(n6663), .B(n11322), .ZN(n6666) );
  BUF_X1 U7700 ( .A(data_addr_i[29]), .Z(n11303) );
  XNOR2_X1 U7701 ( .A(n6664), .B(n11303), .ZN(n6665) );
  NAND4_X1 U7702 ( .A1(n6668), .A2(n6667), .A3(n6666), .A4(n6665), .ZN(n6669)
         );
  XNOR2_X1 U7704 ( .A(n6671), .B(n12123), .ZN(n6692) );
  NAND2_X1 U7705 ( .A1(data_addr_o_10_), .A2(n3912), .ZN(n11760) );
  OAI21_X1 U7706 ( .B1(n10501), .B2(n6672), .A(n11760), .ZN(n11770) );
  AOI21_X1 U7707 ( .B1(n11259), .B2(n323), .A(n6673), .ZN(n6675) );
  NAND2_X1 U7708 ( .A1(data_addr_o_4_), .A2(n6674), .ZN(n11766) );
  NAND4_X1 U7709 ( .A1(n11764), .A2(n6675), .A3(n11766), .A4(n11798), .ZN(
        n6676) );
  NOR3_X1 U7710 ( .A1(n11770), .A2(n11763), .A3(n6676), .ZN(n6687) );
  NAND2_X1 U7711 ( .A1(data_addr_o_6_), .A2(n3888), .ZN(n11782) );
  NAND2_X1 U7712 ( .A1(data_addr_o_5_), .A2(n3887), .ZN(n11783) );
  AND2_X1 U7713 ( .A1(n11782), .A2(n11783), .ZN(n6682) );
  INV_X1 U7714 ( .A(n11291), .ZN(n11255) );
  OAI22_X1 U7715 ( .A1(n10958), .A2(n6677), .B1(n11259), .B2(n323), .ZN(n6678)
         );
  INV_X1 U7716 ( .A(n6678), .ZN(n6679) );
  OAI211_X1 U7717 ( .C1(n11255), .C2(n3887), .A(n6680), .B(n6679), .ZN(n11800)
         );
  INV_X1 U7718 ( .A(n11800), .ZN(n6681) );
  NAND2_X1 U7719 ( .A1(n8246), .A2(n3955), .ZN(n11777) );
  NAND4_X1 U7720 ( .A1(n6682), .A2(n6681), .A3(n11777), .A4(n11778), .ZN(n6685) );
  NAND2_X1 U7721 ( .A1(n6649), .A2(n3959), .ZN(n11788) );
  NAND2_X1 U7722 ( .A1(data_addr_o_12_), .A2(n6683), .ZN(n11801) );
  NAND2_X1 U7723 ( .A1(n11788), .A2(n11801), .ZN(n6684) );
  NOR2_X1 U7724 ( .A1(n6685), .A2(n6684), .ZN(n6686) );
  NAND4_X1 U7725 ( .A1(n6687), .A2(n6686), .A3(n11809), .A4(n11806), .ZN(n6690) );
  XNOR2_X1 U7726 ( .A(n11793), .B(n7995), .ZN(n6689) );
  NOR2_X1 U7727 ( .A1(n6690), .A2(n6689), .ZN(n6691) );
  NAND3_X1 U7728 ( .A1(n11759), .A2(n6692), .A3(n6691), .ZN(n6693) );
  NAND2_X1 U7729 ( .A1(n6694), .A2(n6693), .ZN(n6697) );
  MUX2_X1 U7730 ( .A(pmp_cfg_i[120]), .B(pmp_cfg_i[121]), .S(n11019), .Z(n6696) );
  AND2_X1 U7731 ( .A1(n6695), .A2(n6696), .ZN(n11812) );
  AOI22_X1 U7732 ( .A1(n11154), .A2(n6698), .B1(n6697), .B2(n11812), .ZN(n9341) );
  INV_X1 U7733 ( .A(data_addr_o_14_), .ZN(n10000) );
  NOR2_X1 U7734 ( .A1(pmp_addr_i[300]), .A2(n10000), .ZN(n6699) );
  NOR2_X1 U7735 ( .A1(pmp_addr_i[301]), .A2(n10338), .ZN(n6742) );
  NOR2_X1 U7736 ( .A1(n6699), .A2(n6742), .ZN(n6701) );
  NOR2_X1 U7737 ( .A1(pmp_addr_i[302]), .A2(n10047), .ZN(n6700) );
  NOR2_X1 U7738 ( .A1(pmp_addr_i[303]), .A2(n7995), .ZN(n6745) );
  NOR2_X1 U7739 ( .A1(n6700), .A2(n6745), .ZN(n6748) );
  NAND2_X1 U7740 ( .A1(n6701), .A2(n6748), .ZN(n6750) );
  NOR2_X1 U7741 ( .A1(pmp_addr_i[296]), .A2(n6141), .ZN(n6702) );
  NOR2_X1 U7742 ( .A1(pmp_addr_i[297]), .A2(n9508), .ZN(n6733) );
  NOR2_X1 U7743 ( .A1(n6702), .A2(n6733), .ZN(n6704) );
  NOR2_X1 U7744 ( .A1(pmp_addr_i[298]), .A2(n7976), .ZN(n6703) );
  NOR2_X1 U7746 ( .A1(pmp_addr_i[299]), .A2(n11006), .ZN(n6736) );
  NOR2_X1 U7747 ( .A1(n6703), .A2(n6736), .ZN(n6739) );
  NAND2_X1 U7748 ( .A1(n6704), .A2(n6739), .ZN(n6705) );
  NOR2_X1 U7749 ( .A1(n6750), .A2(n6705), .ZN(n6754) );
  NOR2_X1 U7750 ( .A1(pmp_addr_i[290]), .A2(n10351), .ZN(n6706) );
  NOR2_X1 U7751 ( .A1(pmp_addr_i[291]), .A2(n10346), .ZN(n6712) );
  NOR2_X1 U7752 ( .A1(n6706), .A2(n6712), .ZN(n6715) );
  INV_X1 U7753 ( .A(n22), .ZN(n9350) );
  NOR2_X1 U7754 ( .A1(pmp_addr_i[289]), .A2(n9350), .ZN(n6709) );
  NAND2_X1 U7755 ( .A1(pmp_addr_i[288]), .A2(n10651), .ZN(n6708) );
  NAND2_X1 U7756 ( .A1(pmp_addr_i[289]), .A2(n9350), .ZN(n6707) );
  OAI21_X1 U7757 ( .B1(n6709), .B2(n6708), .A(n6707), .ZN(n6714) );
  NAND2_X1 U7758 ( .A1(pmp_addr_i[290]), .A2(n10351), .ZN(n6711) );
  NAND2_X1 U7759 ( .A1(pmp_addr_i[291]), .A2(n10346), .ZN(n6710) );
  OAI21_X1 U7760 ( .B1(n6712), .B2(n6711), .A(n6710), .ZN(n6713) );
  AOI21_X1 U7761 ( .B1(n6715), .B2(n6714), .A(n6713), .ZN(n6730) );
  NOR2_X1 U7762 ( .A1(pmp_addr_i[292]), .A2(n10362), .ZN(n6716) );
  NOR2_X1 U7763 ( .A1(pmp_addr_i[293]), .A2(n6400), .ZN(n6721) );
  NOR2_X1 U7764 ( .A1(n6716), .A2(n6721), .ZN(n6718) );
  NOR2_X1 U7765 ( .A1(pmp_addr_i[294]), .A2(n29), .ZN(n6717) );
  INV_X1 U7766 ( .A(data_addr_o_9_), .ZN(n9367) );
  NOR2_X1 U7767 ( .A1(pmp_addr_i[295]), .A2(n9367), .ZN(n6724) );
  NOR2_X1 U7768 ( .A1(n6717), .A2(n6724), .ZN(n6727) );
  NAND2_X1 U7769 ( .A1(n6718), .A2(n6727), .ZN(n6729) );
  NAND2_X1 U7770 ( .A1(pmp_addr_i[292]), .A2(n9363), .ZN(n6720) );
  NAND2_X1 U7771 ( .A1(pmp_addr_i[293]), .A2(n10697), .ZN(n6719) );
  OAI21_X1 U7772 ( .B1(n6721), .B2(n6720), .A(n6719), .ZN(n6726) );
  NAND2_X1 U7773 ( .A1(pmp_addr_i[294]), .A2(n29), .ZN(n6723) );
  NAND2_X1 U7774 ( .A1(pmp_addr_i[295]), .A2(n6140), .ZN(n6722) );
  OAI21_X1 U7775 ( .B1(n6724), .B2(n6723), .A(n6722), .ZN(n6725) );
  AOI21_X1 U7776 ( .B1(n6727), .B2(n6726), .A(n6725), .ZN(n6728) );
  OAI21_X1 U7777 ( .B1(n6730), .B2(n6729), .A(n6728), .ZN(n6753) );
  NAND2_X1 U7778 ( .A1(pmp_addr_i[296]), .A2(n6141), .ZN(n6732) );
  NAND2_X1 U7779 ( .A1(pmp_addr_i[297]), .A2(n9508), .ZN(n6731) );
  OAI21_X1 U7780 ( .B1(n6733), .B2(n6732), .A(n6731), .ZN(n6738) );
  NAND2_X1 U7781 ( .A1(pmp_addr_i[298]), .A2(n7472), .ZN(n6735) );
  NAND2_X1 U7782 ( .A1(pmp_addr_i[299]), .A2(n10342), .ZN(n6734) );
  OAI21_X1 U7783 ( .B1(n6736), .B2(n6735), .A(n6734), .ZN(n6737) );
  AOI21_X1 U7784 ( .B1(n6739), .B2(n6738), .A(n6737), .ZN(n6751) );
  NAND2_X1 U7785 ( .A1(pmp_addr_i[300]), .A2(n6154), .ZN(n6741) );
  NAND2_X1 U7786 ( .A1(pmp_addr_i[301]), .A2(n9125), .ZN(n6740) );
  OAI21_X1 U7787 ( .B1(n6742), .B2(n6741), .A(n6740), .ZN(n6747) );
  NAND2_X1 U7788 ( .A1(pmp_addr_i[302]), .A2(n7990), .ZN(n6744) );
  NAND2_X1 U7789 ( .A1(pmp_addr_i[303]), .A2(n8444), .ZN(n6743) );
  OAI21_X1 U7790 ( .B1(n6745), .B2(n6744), .A(n6743), .ZN(n6746) );
  AOI21_X1 U7791 ( .B1(n6748), .B2(n6747), .A(n6746), .ZN(n6749) );
  OAI21_X1 U7792 ( .B1(n6751), .B2(n6750), .A(n6749), .ZN(n6752) );
  AOI21_X1 U7793 ( .B1(n6754), .B2(n6753), .A(n6752), .ZN(n6812) );
  NOR2_X1 U7794 ( .A1(pmp_addr_i[304]), .A2(n10403), .ZN(n6755) );
  NOR2_X1 U7795 ( .A1(pmp_addr_i[305]), .A2(n10414), .ZN(n6770) );
  NOR2_X1 U7796 ( .A1(n6755), .A2(n6770), .ZN(n6757) );
  NOR2_X1 U7797 ( .A1(pmp_addr_i[306]), .A2(n6188), .ZN(n6756) );
  NOR2_X1 U7798 ( .A1(pmp_addr_i[307]), .A2(n6192), .ZN(n6773) );
  NOR2_X1 U7799 ( .A1(n6756), .A2(n6773), .ZN(n6776) );
  NAND2_X1 U7800 ( .A1(n6757), .A2(n6776), .ZN(n6761) );
  NOR2_X1 U7801 ( .A1(pmp_addr_i[308]), .A2(n9425), .ZN(n6758) );
  INV_X1 U7802 ( .A(n10737), .ZN(n10064) );
  NOR2_X1 U7803 ( .A1(pmp_addr_i[309]), .A2(n10064), .ZN(n6779) );
  NOR2_X1 U7804 ( .A1(n6758), .A2(n6779), .ZN(n6760) );
  NOR2_X1 U7805 ( .A1(pmp_addr_i[310]), .A2(n9163), .ZN(n6759) );
  NOR2_X1 U7806 ( .A1(pmp_addr_i[311]), .A2(n6462), .ZN(n6782) );
  NOR2_X1 U7807 ( .A1(n6759), .A2(n6782), .ZN(n6785) );
  NAND2_X1 U7808 ( .A1(n6760), .A2(n6785), .ZN(n6787) );
  NOR2_X1 U7809 ( .A1(n6761), .A2(n6787), .ZN(n6767) );
  NOR2_X1 U7810 ( .A1(pmp_addr_i[312]), .A2(n10439), .ZN(n6762) );
  NOR2_X1 U7811 ( .A1(pmp_addr_i[313]), .A2(n10096), .ZN(n6791) );
  NOR2_X1 U7812 ( .A1(n6762), .A2(n6791), .ZN(n6764) );
  NOR2_X1 U7813 ( .A1(pmp_addr_i[314]), .A2(n10443), .ZN(n6763) );
  NOR2_X1 U7814 ( .A1(pmp_addr_i[315]), .A2(n10100), .ZN(n6794) );
  NOR2_X1 U7815 ( .A1(n6763), .A2(n6794), .ZN(n6797) );
  NAND2_X1 U7816 ( .A1(n6764), .A2(n6797), .ZN(n6766) );
  NOR2_X1 U7817 ( .A1(pmp_addr_i[316]), .A2(n8494), .ZN(n6765) );
  NOR2_X1 U7818 ( .A1(pmp_addr_i[317]), .A2(data_addr_o_31__BAR), .ZN(n6800)
         );
  OR2_X1 U7819 ( .A1(n6765), .A2(n6800), .ZN(n6805) );
  NOR2_X1 U7820 ( .A1(n6766), .A2(n6805), .ZN(n6808) );
  NAND2_X1 U7821 ( .A1(n6767), .A2(n6808), .ZN(n6811) );
  NAND2_X1 U7823 ( .A1(pmp_addr_i[304]), .A2(n12184), .ZN(n6769) );
  NAND2_X1 U7824 ( .A1(pmp_addr_i[305]), .A2(n10414), .ZN(n6768) );
  OAI21_X1 U7825 ( .B1(n6770), .B2(n6769), .A(n6768), .ZN(n6775) );
  NAND2_X1 U7826 ( .A1(pmp_addr_i[306]), .A2(n6188), .ZN(n6772) );
  NAND2_X1 U7827 ( .A1(pmp_addr_i[307]), .A2(n9418), .ZN(n6771) );
  OAI21_X1 U7828 ( .B1(n6773), .B2(n6772), .A(n6771), .ZN(n6774) );
  AOI21_X1 U7829 ( .B1(n6776), .B2(n6775), .A(n6774), .ZN(n6788) );
  NAND2_X1 U7830 ( .A1(pmp_addr_i[308]), .A2(n9425), .ZN(n6778) );
  NAND2_X1 U7831 ( .A1(pmp_addr_i[309]), .A2(n10064), .ZN(n6777) );
  OAI21_X1 U7832 ( .B1(n6779), .B2(n6778), .A(n6777), .ZN(n6784) );
  NAND2_X1 U7833 ( .A1(pmp_addr_i[310]), .A2(n10428), .ZN(n6781) );
  NAND2_X1 U7834 ( .A1(pmp_addr_i[311]), .A2(n6462), .ZN(n6780) );
  OAI21_X1 U7835 ( .B1(n6782), .B2(n6781), .A(n6780), .ZN(n6783) );
  AOI21_X1 U7836 ( .B1(n6785), .B2(n6784), .A(n6783), .ZN(n6786) );
  OAI21_X1 U7837 ( .B1(n6788), .B2(n6787), .A(n6786), .ZN(n6809) );
  NAND2_X1 U7838 ( .A1(pmp_addr_i[312]), .A2(n6202), .ZN(n6790) );
  NAND2_X1 U7839 ( .A1(pmp_addr_i[313]), .A2(n10096), .ZN(n6789) );
  OAI21_X1 U7840 ( .B1(n6791), .B2(n6790), .A(n6789), .ZN(n6796) );
  NAND2_X1 U7841 ( .A1(pmp_addr_i[314]), .A2(n10443), .ZN(n6793) );
  NAND2_X1 U7842 ( .A1(pmp_addr_i[315]), .A2(n10100), .ZN(n6792) );
  OAI21_X1 U7843 ( .B1(n6794), .B2(n6793), .A(n6792), .ZN(n6795) );
  AOI21_X1 U7844 ( .B1(n6797), .B2(n6796), .A(n6795), .ZN(n6806) );
  NAND2_X1 U7845 ( .A1(pmp_addr_i[316]), .A2(n8814), .ZN(n6799) );
  NAND2_X1 U7846 ( .A1(pmp_addr_i[317]), .A2(data_addr_o_31__BAR), .ZN(n6798)
         );
  OAI21_X1 U7847 ( .B1(n6800), .B2(n6799), .A(n6798), .ZN(n6803) );
  INV_X1 U7848 ( .A(n6801), .ZN(n6802) );
  NOR2_X1 U7849 ( .A1(n6803), .A2(n6802), .ZN(n6804) );
  OAI21_X1 U7850 ( .B1(n6806), .B2(n6805), .A(n6804), .ZN(n6807) );
  AOI21_X1 U7851 ( .B1(n6809), .B2(n6808), .A(n6807), .ZN(n6810) );
  OAI21_X1 U7852 ( .B1(n6812), .B2(n6811), .A(n6810), .ZN(n6936) );
  INV_X1 U7853 ( .A(n11821), .ZN(n6875) );
  NOR2_X1 U7855 ( .A1(n6875), .A2(n11014), .ZN(n6814) );
  NOR2_X1 U7856 ( .A1(n2283), .A2(n6813), .ZN(n6876) );
  NOR2_X1 U7857 ( .A1(n6814), .A2(n6876), .ZN(n6816) );
  NOR2_X1 U7858 ( .A1(n2216), .A2(n10857), .ZN(n6815) );
  NOR2_X1 U7859 ( .A1(n2208), .A2(n10886), .ZN(n6880) );
  NOR2_X1 U7860 ( .A1(n6815), .A2(n6880), .ZN(n6883) );
  NAND2_X1 U7861 ( .A1(n6816), .A2(n6883), .ZN(n6820) );
  NOR2_X1 U7862 ( .A1(n2166), .A2(n10887), .ZN(n6817) );
  NOR2_X1 U7863 ( .A1(n2170), .A2(n10891), .ZN(n6886) );
  NOR2_X1 U7864 ( .A1(n6817), .A2(n6886), .ZN(n6819) );
  BUF_X1 U7865 ( .A(data_addr_i[22]), .Z(n9915) );
  NOR2_X1 U7866 ( .A1(n2162), .A2(n9915), .ZN(n6818) );
  NOR2_X1 U7867 ( .A1(n2190), .A2(n10737), .ZN(n6889) );
  NOR2_X1 U7868 ( .A1(n6818), .A2(n6889), .ZN(n6892) );
  NAND2_X1 U7869 ( .A1(n6819), .A2(n6892), .ZN(n6894) );
  NOR2_X1 U7870 ( .A1(n6820), .A2(n6894), .ZN(n6898) );
  NAND2_X1 U7871 ( .A1(n6865), .A2(n11334), .ZN(n6951) );
  INV_X1 U7872 ( .A(n6951), .ZN(n6821) );
  NAND2_X1 U7873 ( .A1(n6866), .A2(n9941), .ZN(n6952) );
  INV_X1 U7874 ( .A(n6952), .ZN(n6868) );
  NOR2_X1 U7875 ( .A1(n6821), .A2(n6868), .ZN(n6871) );
  INV_X1 U7876 ( .A(data_addr_o_12_), .ZN(n10005) );
  NAND2_X1 U7877 ( .A1(n6859), .A2(n10005), .ZN(n6944) );
  OR2_X1 U7878 ( .A1(n8246), .A2(n6982), .ZN(n6823) );
  NAND2_X1 U7879 ( .A1(n6944), .A2(n6823), .ZN(n6824) );
  NAND2_X1 U7880 ( .A1(n6862), .A2(n11006), .ZN(n6945) );
  INV_X1 U7881 ( .A(n6945), .ZN(n6863) );
  NOR2_X1 U7882 ( .A1(n6824), .A2(n6863), .ZN(n6825) );
  NAND2_X1 U7883 ( .A1(n6871), .A2(n6825), .ZN(n6874) );
  INV_X1 U7884 ( .A(n6984), .ZN(n6826) );
  NOR2_X1 U7885 ( .A1(n10129), .A2(n6826), .ZN(n6829) );
  INV_X1 U7886 ( .A(n10473), .ZN(n10130) );
  INV_X1 U7887 ( .A(n6989), .ZN(n6827) );
  NOR2_X1 U7888 ( .A1(n10130), .A2(n6827), .ZN(n6828) );
  NAND2_X1 U7889 ( .A1(n10130), .A2(n6827), .ZN(n11833) );
  OAI21_X1 U7890 ( .B1(n6829), .B2(n6828), .A(n11833), .ZN(n6832) );
  NAND2_X1 U7891 ( .A1(n12058), .A2(n6830), .ZN(n6992) );
  AND2_X1 U7892 ( .A1(n10135), .A2(n6983), .ZN(n6831) );
  AOI21_X1 U7893 ( .B1(n6832), .B2(n6992), .A(n6831), .ZN(n6840) );
  OR2_X1 U7894 ( .A1(n10824), .A2(n6996), .ZN(n6835) );
  OR2_X1 U7895 ( .A1(n10655), .A2(n6937), .ZN(n6837) );
  NAND2_X1 U7896 ( .A1(n6835), .A2(n6837), .ZN(n6839) );
  AND2_X1 U7897 ( .A1(n10824), .A2(n6996), .ZN(n6836) );
  AND2_X1 U7898 ( .A1(n10655), .A2(n6937), .ZN(n11857) );
  AOI21_X1 U7899 ( .B1(n6837), .B2(n6836), .A(n11857), .ZN(n6838) );
  OAI21_X1 U7900 ( .B1(n6840), .B2(n6839), .A(n6838), .ZN(n6858) );
  OR2_X1 U7902 ( .A1(n10494), .A2(n6999), .ZN(n6849) );
  OR2_X1 U7903 ( .A1(n7816), .A2(n6995), .ZN(n6843) );
  NAND2_X1 U7904 ( .A1(n6849), .A2(n6843), .ZN(n6846) );
  OR2_X1 U7905 ( .A1(data_addr_o_9_), .A2(n6998), .ZN(n6845) );
  INV_X1 U7906 ( .A(n7820), .ZN(n10838) );
  OR2_X1 U7907 ( .A1(n10838), .A2(n6981), .ZN(n6852) );
  NAND2_X1 U7908 ( .A1(n6845), .A2(n6852), .ZN(n6854) );
  NOR2_X1 U7909 ( .A1(n6846), .A2(n6854), .ZN(n6857) );
  AND2_X1 U7910 ( .A1(data_addr_o_7_), .A2(n6995), .ZN(n6848) );
  AND2_X1 U7911 ( .A1(n10494), .A2(n6999), .ZN(n6847) );
  AOI21_X1 U7912 ( .B1(n6849), .B2(n6848), .A(n6847), .ZN(n6855) );
  AND2_X1 U7913 ( .A1(data_addr_o_9_), .A2(n6998), .ZN(n6851) );
  AND2_X1 U7914 ( .A1(n10838), .A2(n6981), .ZN(n6850) );
  AOI21_X1 U7915 ( .B1(n6852), .B2(n6851), .A(n6850), .ZN(n6853) );
  OAI21_X1 U7916 ( .B1(n6855), .B2(n6854), .A(n6853), .ZN(n6856) );
  AOI21_X1 U7917 ( .B1(n6858), .B2(n6857), .A(n6856), .ZN(n6873) );
  AND2_X1 U7918 ( .A1(data_addr_o_11_), .A2(n6982), .ZN(n6861) );
  OR2_X1 U7919 ( .A1(n6859), .A2(n7472), .ZN(n11861) );
  INV_X1 U7920 ( .A(n11861), .ZN(n6860) );
  AOI21_X1 U7921 ( .B1(n6944), .B2(n6861), .A(n6860), .ZN(n6864) );
  OR2_X1 U7922 ( .A1(n6862), .A2(n11006), .ZN(n11826) );
  OAI21_X1 U7923 ( .B1(n6864), .B2(n6863), .A(n11826), .ZN(n6870) );
  NOR2_X1 U7924 ( .A1(n6865), .A2(n10518), .ZN(n11868) );
  INV_X1 U7925 ( .A(n11868), .ZN(n6867) );
  OR2_X1 U7926 ( .A1(n6866), .A2(n9941), .ZN(n11869) );
  OAI21_X1 U7927 ( .B1(n6868), .B2(n6867), .A(n11869), .ZN(n6869) );
  AOI21_X1 U7928 ( .B1(n6871), .B2(n6870), .A(n6869), .ZN(n6872) );
  OAI21_X1 U7929 ( .B1(n6874), .B2(n6873), .A(n6872), .ZN(n6897) );
  NAND2_X1 U7930 ( .A1(n6875), .A2(n11014), .ZN(n6877) );
  OR2_X1 U7931 ( .A1(n6947), .A2(n8444), .ZN(n11823) );
  OAI21_X1 U7932 ( .B1(n6877), .B2(n6876), .A(n11823), .ZN(n6882) );
  NAND2_X1 U7933 ( .A1(n2216), .A2(n10857), .ZN(n6879) );
  NAND2_X1 U7934 ( .A1(n2208), .A2(n11283), .ZN(n6878) );
  OAI21_X1 U7935 ( .B1(n6880), .B2(n6879), .A(n6878), .ZN(n6881) );
  AOI21_X1 U7936 ( .B1(n6883), .B2(n6882), .A(n6881), .ZN(n6895) );
  NAND2_X1 U7937 ( .A1(n2166), .A2(data_addr_o_20_), .ZN(n6885) );
  NAND2_X1 U7938 ( .A1(n2170), .A2(n10891), .ZN(n6884) );
  OAI21_X1 U7939 ( .B1(n6886), .B2(n6885), .A(n6884), .ZN(n6891) );
  NAND2_X1 U7940 ( .A1(n2162), .A2(n9915), .ZN(n6888) );
  NAND2_X1 U7941 ( .A1(n2190), .A2(n10737), .ZN(n6887) );
  OAI21_X1 U7942 ( .B1(n6889), .B2(n6888), .A(n6887), .ZN(n6890) );
  AOI21_X1 U7943 ( .B1(n6892), .B2(n6891), .A(n6890), .ZN(n6893) );
  OAI21_X1 U7944 ( .B1(n6895), .B2(n6894), .A(n6893), .ZN(n6896) );
  AOI21_X1 U7945 ( .B1(n6898), .B2(n6897), .A(n6896), .ZN(n6933) );
  NOR2_X1 U7946 ( .A1(n2154), .A2(n10904), .ZN(n6899) );
  NOR2_X1 U7947 ( .A1(n2176), .A2(n10746), .ZN(n6912) );
  NOR2_X1 U7948 ( .A1(n6899), .A2(n6912), .ZN(n6915) );
  BUF_X1 U7949 ( .A(data_addr_i[24]), .Z(n10738) );
  NOR2_X1 U7950 ( .A1(n2159), .A2(n10738), .ZN(n6900) );
  NOR2_X1 U7951 ( .A1(n2193), .A2(n9923), .ZN(n6909) );
  NOR2_X1 U7952 ( .A1(n6900), .A2(n6909), .ZN(n6901) );
  NAND2_X1 U7953 ( .A1(n6915), .A2(n6901), .ZN(n6905) );
  NOR2_X1 U7954 ( .A1(n2200), .A2(n12123), .ZN(n6922) );
  NOR2_X1 U7955 ( .A1(n2143), .A2(n10919), .ZN(n6902) );
  NOR2_X1 U7956 ( .A1(n6922), .A2(n6902), .ZN(n6925) );
  NOR2_X1 U7957 ( .A1(n2149), .A2(n10747), .ZN(n6903) );
  INV_X1 U7958 ( .A(n6971), .ZN(n6916) );
  NOR2_X1 U7959 ( .A1(n6916), .A2(data_addr_o_29_), .ZN(n6919) );
  NOR2_X1 U7960 ( .A1(n6903), .A2(n6919), .ZN(n6904) );
  NAND2_X1 U7961 ( .A1(n6925), .A2(n6904), .ZN(n6927) );
  NOR2_X1 U7962 ( .A1(n6905), .A2(n6927), .ZN(n6906) );
  NOR2_X1 U7963 ( .A1(pmp_addr_i[287]), .A2(pmp_addr_i[286]), .ZN(n6929) );
  NAND2_X1 U7964 ( .A1(n6906), .A2(n6929), .ZN(n6932) );
  NAND2_X1 U7965 ( .A1(n2159), .A2(n10738), .ZN(n6908) );
  NAND2_X1 U7966 ( .A1(n2193), .A2(n9923), .ZN(n6907) );
  OAI21_X1 U7967 ( .B1(n6909), .B2(n6908), .A(n6907), .ZN(n6914) );
  NAND2_X1 U7968 ( .A1(n2154), .A2(n10904), .ZN(n6911) );
  NAND2_X1 U7969 ( .A1(n2176), .A2(n10746), .ZN(n6910) );
  OAI21_X1 U7970 ( .B1(n6912), .B2(n6911), .A(n6910), .ZN(n6913) );
  AOI21_X1 U7971 ( .B1(n6915), .B2(n6914), .A(n6913), .ZN(n6928) );
  NAND2_X1 U7972 ( .A1(n2149), .A2(n10747), .ZN(n6918) );
  NAND2_X1 U7973 ( .A1(n6916), .A2(data_addr_o_29_), .ZN(n6917) );
  OAI21_X1 U7974 ( .B1(n6919), .B2(n6918), .A(n6917), .ZN(n6924) );
  NAND2_X1 U7975 ( .A1(n2143), .A2(n10919), .ZN(n6921) );
  NAND2_X1 U7976 ( .A1(n2200), .A2(n12123), .ZN(n6920) );
  OAI21_X1 U7977 ( .B1(n6922), .B2(n6921), .A(n6920), .ZN(n6923) );
  AOI21_X1 U7978 ( .B1(n6925), .B2(n6924), .A(n6923), .ZN(n6926) );
  OAI21_X1 U7979 ( .B1(n6928), .B2(n6927), .A(n6926), .ZN(n6930) );
  NAND2_X1 U7980 ( .A1(n6930), .A2(n6929), .ZN(n6931) );
  OAI21_X1 U7981 ( .B1(n6933), .B2(n6932), .A(n6931), .ZN(n6934) );
  NAND3_X1 U7982 ( .A1(n6936), .A2(n6935), .A3(n6934), .ZN(n7012) );
  OAI22_X1 U7983 ( .A1(n6995), .A2(n7816), .B1(n10953), .B2(n6937), .ZN(n6938)
         );
  AOI21_X1 U7984 ( .B1(n6141), .B2(n6939), .A(n6938), .ZN(n6943) );
  OAI22_X1 U7985 ( .A1(data_addr_o_9_), .A2(n6998), .B1(n10494), .B2(n6999), 
        .ZN(n6941) );
  NOR2_X1 U7986 ( .A1(data_addr_o_11_), .A2(n6982), .ZN(n6940) );
  NOR2_X1 U7987 ( .A1(n6941), .A2(n6940), .ZN(n6942) );
  NAND4_X1 U7988 ( .A1(n6945), .A2(n6944), .A3(n6943), .A4(n6942), .ZN(n6946)
         );
  AOI21_X1 U7989 ( .B1(n6947), .B2(n8757), .A(n6946), .ZN(n6950) );
  XNOR2_X1 U7990 ( .A(n6948), .B(n10967), .ZN(n6949) );
  AND4_X1 U7991 ( .A1(n6952), .A2(n6951), .A3(n6950), .A4(n6949), .ZN(n6980)
         );
  BUF_X1 U7992 ( .A(data_addr_i[19]), .Z(n9846) );
  XNOR2_X1 U7993 ( .A(n6953), .B(n9846), .ZN(n6960) );
  XNOR2_X1 U7994 ( .A(n6954), .B(n9935), .ZN(n6959) );
  XNOR2_X1 U7995 ( .A(n6955), .B(n10202), .ZN(n6958) );
  BUF_X1 U7996 ( .A(data_addr_i[22]), .Z(n9529) );
  XNOR2_X1 U7997 ( .A(n6956), .B(n9529), .ZN(n6957) );
  AND4_X1 U7998 ( .A1(n6960), .A2(n6959), .A3(n6958), .A4(n6957), .ZN(n6979)
         );
  XNOR2_X1 U7999 ( .A(n6961), .B(n10898), .ZN(n6968) );
  XNOR2_X1 U8000 ( .A(n6962), .B(n10629), .ZN(n6967) );
  BUF_X1 U8001 ( .A(data_addr_i[25]), .Z(n10903) );
  XNOR2_X1 U8002 ( .A(n6963), .B(n10903), .ZN(n6966) );
  BUF_X1 U8003 ( .A(data_addr_i[26]), .Z(n10267) );
  XNOR2_X1 U8004 ( .A(n6964), .B(n10267), .ZN(n6965) );
  AND4_X1 U8005 ( .A1(n6968), .A2(n6967), .A3(n6966), .A4(n6965), .ZN(n6978)
         );
  BUF_X1 U8006 ( .A(data_addr_i[27]), .Z(n9886) );
  XNOR2_X1 U8007 ( .A(n6969), .B(n9886), .ZN(n6976) );
  XNOR2_X1 U8008 ( .A(n6970), .B(n10635), .ZN(n6975) );
  BUF_X1 U8009 ( .A(data_addr_i[29]), .Z(n9955) );
  XNOR2_X1 U8010 ( .A(n6971), .B(n9955), .ZN(n6974) );
  XNOR2_X1 U8011 ( .A(n6972), .B(data_addr_o_30_), .ZN(n6973) );
  AND4_X1 U8012 ( .A1(n6976), .A2(n6975), .A3(n6974), .A4(n6973), .ZN(n6977)
         );
  NAND4_X1 U8013 ( .A1(n6980), .A2(n6979), .A3(n6978), .A4(n6977), .ZN(n11876)
         );
  NAND2_X1 U8014 ( .A1(data_addr_o_10_), .A2(n6981), .ZN(n11839) );
  NAND2_X1 U8015 ( .A1(n10508), .A2(n6982), .ZN(n11851) );
  NAND2_X1 U8016 ( .A1(data_addr_o_4_), .A2(n6983), .ZN(n11830) );
  INV_X1 U8017 ( .A(n6985), .ZN(n6986) );
  AOI21_X1 U8018 ( .B1(n11259), .B2(n6826), .A(n6986), .ZN(n6987) );
  NAND3_X1 U8019 ( .A1(n11830), .A2(n6987), .A3(n11833), .ZN(n6988) );
  NOR2_X1 U8020 ( .A1(n11857), .A2(n6988), .ZN(n6994) );
  OAI22_X1 U8021 ( .A1(n10958), .A2(n6827), .B1(n11259), .B2(n6826), .ZN(n6990) );
  INV_X1 U8022 ( .A(n6990), .ZN(n6991) );
  OAI211_X1 U8023 ( .C1(n11255), .C2(n6996), .A(n6992), .B(n6991), .ZN(n6993)
         );
  INV_X1 U8024 ( .A(n6993), .ZN(n11837) );
  NAND4_X1 U8025 ( .A1(n11839), .A2(n11851), .A3(n6994), .A4(n11837), .ZN(
        n7001) );
  NAND2_X1 U8026 ( .A1(data_addr_o_7_), .A2(n6995), .ZN(n11841) );
  NAND2_X1 U8027 ( .A1(data_addr_o_5_), .A2(n6996), .ZN(n6997) );
  AND2_X1 U8028 ( .A1(n11841), .A2(n6997), .ZN(n11843) );
  NAND2_X1 U8029 ( .A1(data_addr_o_9_), .A2(n6998), .ZN(n11847) );
  NAND2_X1 U8030 ( .A1(n10836), .A2(n6999), .ZN(n11848) );
  NAND3_X1 U8031 ( .A1(n11843), .A2(n11847), .A3(n11848), .ZN(n7000) );
  NOR2_X1 U8032 ( .A1(n7001), .A2(n7000), .ZN(n7002) );
  NAND4_X1 U8033 ( .A1(n11823), .A2(n7002), .A3(n11826), .A4(n11861), .ZN(
        n7003) );
  NOR2_X1 U8034 ( .A1(n11868), .A2(n7003), .ZN(n7007) );
  XNOR2_X1 U8035 ( .A(n11821), .B(n11004), .ZN(n7006) );
  XNOR2_X1 U8036 ( .A(n7004), .B(n12123), .ZN(n7005) );
  NAND4_X1 U8037 ( .A1(n7007), .A2(n7006), .A3(n7005), .A4(n11869), .ZN(n7008)
         );
  OR2_X1 U8038 ( .A1(n11876), .A2(n7008), .ZN(n7011) );
  OR2_X1 U8039 ( .A1(n11019), .A2(pmp_cfg_i[72]), .ZN(n7010) );
  OAI211_X1 U8040 ( .C1(pmp_cfg_i[73]), .C2(n11021), .A(n7009), .B(n7010), 
        .ZN(n11827) );
  AOI21_X1 U8041 ( .B1(n7012), .B2(n7011), .A(n11827), .ZN(n8088) );
  INV_X1 U8042 ( .A(n11004), .ZN(n7057) );
  NOR2_X1 U8043 ( .A1(n7057), .A2(pmp_addr_i[238]), .ZN(n7013) );
  NOR2_X1 U8044 ( .A1(n7995), .A2(pmp_addr_i[239]), .ZN(n7060) );
  NOR2_X1 U8045 ( .A1(n7013), .A2(n7060), .ZN(n7063) );
  NOR2_X1 U8046 ( .A1(pmp_addr_i[236]), .A2(n10000), .ZN(n7014) );
  NOR2_X1 U8047 ( .A1(pmp_addr_i[237]), .A2(n9125), .ZN(n7056) );
  NOR2_X1 U8048 ( .A1(n7014), .A2(n7056), .ZN(n7015) );
  NAND2_X1 U8049 ( .A1(n7063), .A2(n7015), .ZN(n7066) );
  NOR2_X1 U8050 ( .A1(pmp_addr_i[232]), .A2(n10701), .ZN(n7016) );
  NOR2_X1 U8051 ( .A1(pmp_addr_i[233]), .A2(n9508), .ZN(n7047) );
  NOR2_X1 U8052 ( .A1(n7016), .A2(n7047), .ZN(n7018) );
  NOR2_X1 U8053 ( .A1(pmp_addr_i[234]), .A2(n7472), .ZN(n7017) );
  NOR2_X1 U8054 ( .A1(pmp_addr_i[235]), .A2(n11006), .ZN(n7050) );
  NOR2_X1 U8055 ( .A1(n7017), .A2(n7050), .ZN(n7053) );
  NAND2_X1 U8056 ( .A1(n7018), .A2(n7053), .ZN(n7019) );
  NOR2_X1 U8057 ( .A1(n7066), .A2(n7019), .ZN(n7069) );
  NOR2_X1 U8058 ( .A1(pmp_addr_i[227]), .A2(n11291), .ZN(n7026) );
  NOR2_X1 U8059 ( .A1(pmp_addr_i[226]), .A2(n8406), .ZN(n7020) );
  NOR2_X1 U8060 ( .A1(n7026), .A2(n7020), .ZN(n7029) );
  NOR2_X1 U8061 ( .A1(pmp_addr_i[225]), .A2(n9350), .ZN(n7023) );
  NAND2_X1 U8062 ( .A1(pmp_addr_i[224]), .A2(n10651), .ZN(n7022) );
  NAND2_X1 U8063 ( .A1(pmp_addr_i[225]), .A2(n9350), .ZN(n7021) );
  OAI21_X1 U8064 ( .B1(n7023), .B2(n7022), .A(n7021), .ZN(n7028) );
  NAND2_X1 U8065 ( .A1(pmp_addr_i[226]), .A2(n10351), .ZN(n7025) );
  NAND2_X1 U8066 ( .A1(pmp_addr_i[227]), .A2(n6127), .ZN(n7024) );
  OAI21_X1 U8067 ( .B1(n7026), .B2(n7025), .A(n7024), .ZN(n7027) );
  AOI21_X1 U8068 ( .B1(n7029), .B2(n7028), .A(n7027), .ZN(n7044) );
  NOR2_X1 U8069 ( .A1(pmp_addr_i[228]), .A2(n10362), .ZN(n7030) );
  NOR2_X1 U8070 ( .A1(pmp_addr_i[229]), .A2(n7152), .ZN(n7035) );
  NOR2_X1 U8071 ( .A1(n7030), .A2(n7035), .ZN(n7032) );
  NOR2_X1 U8072 ( .A1(pmp_addr_i[230]), .A2(n8735), .ZN(n7031) );
  NOR2_X1 U8073 ( .A1(pmp_addr_i[231]), .A2(n9367), .ZN(n7038) );
  NOR2_X1 U8074 ( .A1(n7031), .A2(n7038), .ZN(n7041) );
  NAND2_X1 U8075 ( .A1(n7032), .A2(n7041), .ZN(n7043) );
  NAND2_X1 U8076 ( .A1(pmp_addr_i[228]), .A2(n10362), .ZN(n7034) );
  NAND2_X1 U8077 ( .A1(pmp_addr_i[229]), .A2(n10697), .ZN(n7033) );
  OAI21_X1 U8078 ( .B1(n7035), .B2(n7034), .A(n7033), .ZN(n7040) );
  NAND2_X1 U8079 ( .A1(pmp_addr_i[230]), .A2(n29), .ZN(n7037) );
  NAND2_X1 U8080 ( .A1(pmp_addr_i[231]), .A2(n9367), .ZN(n7036) );
  OAI21_X1 U8081 ( .B1(n7038), .B2(n7037), .A(n7036), .ZN(n7039) );
  AOI21_X1 U8082 ( .B1(n7041), .B2(n7040), .A(n7039), .ZN(n7042) );
  OAI21_X1 U8083 ( .B1(n7044), .B2(n7043), .A(n7042), .ZN(n7068) );
  NAND2_X1 U8084 ( .A1(pmp_addr_i[232]), .A2(n6141), .ZN(n7046) );
  NAND2_X1 U8085 ( .A1(pmp_addr_i[233]), .A2(n7324), .ZN(n7045) );
  OAI21_X1 U8086 ( .B1(n7047), .B2(n7046), .A(n7045), .ZN(n7052) );
  NAND2_X1 U8087 ( .A1(pmp_addr_i[234]), .A2(n7472), .ZN(n7049) );
  NAND2_X1 U8088 ( .A1(pmp_addr_i[235]), .A2(n11006), .ZN(n7048) );
  OAI21_X1 U8089 ( .B1(n7050), .B2(n7049), .A(n7048), .ZN(n7051) );
  AOI21_X1 U8090 ( .B1(n7053), .B2(n7052), .A(n7051), .ZN(n7065) );
  NAND2_X1 U8091 ( .A1(pmp_addr_i[236]), .A2(n10000), .ZN(n7055) );
  NAND2_X1 U8092 ( .A1(pmp_addr_i[237]), .A2(n9125), .ZN(n7054) );
  OAI21_X1 U8093 ( .B1(n7056), .B2(n7055), .A(n7054), .ZN(n7062) );
  NAND2_X1 U8094 ( .A1(n7057), .A2(pmp_addr_i[238]), .ZN(n7059) );
  NAND2_X1 U8095 ( .A1(n7995), .A2(pmp_addr_i[239]), .ZN(n7058) );
  OAI21_X1 U8096 ( .B1(n7060), .B2(n7059), .A(n7058), .ZN(n7061) );
  AOI21_X1 U8097 ( .B1(n7063), .B2(n7062), .A(n7061), .ZN(n7064) );
  OAI21_X1 U8098 ( .B1(n7066), .B2(n7065), .A(n7064), .ZN(n7067) );
  AOI21_X1 U8099 ( .B1(n7069), .B2(n7068), .A(n7067), .ZN(n7125) );
  NOR2_X1 U8100 ( .A1(n9156), .A2(pmp_addr_i[244]), .ZN(n7070) );
  NOR2_X1 U8101 ( .A1(n10764), .A2(pmp_addr_i[245]), .ZN(n7094) );
  NOR2_X1 U8102 ( .A1(n7070), .A2(n7094), .ZN(n7072) );
  NOR2_X1 U8103 ( .A1(n10428), .A2(pmp_addr_i[246]), .ZN(n7071) );
  NOR2_X1 U8104 ( .A1(n7071), .A2(n7097), .ZN(n7100) );
  NAND2_X1 U8105 ( .A1(n7072), .A2(n7100), .ZN(n7102) );
  NOR2_X1 U8106 ( .A1(n6192), .A2(pmp_addr_i[243]), .ZN(n7088) );
  NOR2_X1 U8107 ( .A1(n10754), .A2(pmp_addr_i[242]), .ZN(n7073) );
  NOR2_X1 U8108 ( .A1(n7088), .A2(n7073), .ZN(n7091) );
  NOR2_X1 U8109 ( .A1(n10414), .A2(pmp_addr_i[241]), .ZN(n7085) );
  NOR2_X1 U8110 ( .A1(n10060), .A2(pmp_addr_i[240]), .ZN(n7074) );
  NOR2_X1 U8111 ( .A1(n7085), .A2(n7074), .ZN(n7075) );
  NAND2_X1 U8112 ( .A1(n7091), .A2(n7075), .ZN(n7076) );
  NOR2_X1 U8113 ( .A1(n7102), .A2(n7076), .ZN(n7082) );
  NOR2_X1 U8114 ( .A1(n10439), .A2(pmp_addr_i[248]), .ZN(n7077) );
  NOR2_X1 U8115 ( .A1(n6212), .A2(pmp_addr_i[249]), .ZN(n7106) );
  NOR2_X1 U8116 ( .A1(n7077), .A2(n7106), .ZN(n7079) );
  NOR2_X1 U8117 ( .A1(n10443), .A2(pmp_addr_i[250]), .ZN(n7078) );
  NOR2_X1 U8118 ( .A1(n10782), .A2(pmp_addr_i[251]), .ZN(n7109) );
  NOR2_X1 U8119 ( .A1(n7078), .A2(n7109), .ZN(n7112) );
  NAND2_X1 U8120 ( .A1(n7079), .A2(n7112), .ZN(n7081) );
  NOR2_X1 U8121 ( .A1(n8814), .A2(pmp_addr_i[252]), .ZN(n7080) );
  NOR2_X1 U8122 ( .A1(n10107), .A2(pmp_addr_i[253]), .ZN(n7115) );
  OR2_X1 U8123 ( .A1(n7080), .A2(n7115), .ZN(n7119) );
  NOR2_X1 U8124 ( .A1(n7081), .A2(n7119), .ZN(n7122) );
  NAND2_X1 U8125 ( .A1(n7082), .A2(n7122), .ZN(n7124) );
  NAND2_X1 U8126 ( .A1(n10060), .A2(pmp_addr_i[240]), .ZN(n7084) );
  NAND2_X1 U8127 ( .A1(n9414), .A2(pmp_addr_i[241]), .ZN(n7083) );
  OAI21_X1 U8128 ( .B1(n7085), .B2(n7084), .A(n7083), .ZN(n7090) );
  NAND2_X1 U8129 ( .A1(n10754), .A2(pmp_addr_i[242]), .ZN(n7087) );
  NAND2_X1 U8130 ( .A1(n9418), .A2(pmp_addr_i[243]), .ZN(n7086) );
  OAI21_X1 U8131 ( .B1(n7088), .B2(n7087), .A(n7086), .ZN(n7089) );
  AOI21_X1 U8132 ( .B1(n7091), .B2(n7090), .A(n7089), .ZN(n7103) );
  NAND2_X1 U8133 ( .A1(n9425), .A2(pmp_addr_i[244]), .ZN(n7093) );
  NAND2_X1 U8134 ( .A1(n10764), .A2(pmp_addr_i[245]), .ZN(n7092) );
  OAI21_X1 U8135 ( .B1(n7094), .B2(n7093), .A(n7092), .ZN(n7099) );
  NAND2_X1 U8136 ( .A1(n10428), .A2(pmp_addr_i[246]), .ZN(n7096) );
  OAI21_X1 U8137 ( .B1(n7097), .B2(n7096), .A(n7095), .ZN(n7098) );
  AOI21_X1 U8138 ( .B1(n7100), .B2(n7099), .A(n7098), .ZN(n7101) );
  OAI21_X1 U8139 ( .B1(n7103), .B2(n7102), .A(n7101), .ZN(n7123) );
  NAND2_X1 U8140 ( .A1(n6202), .A2(pmp_addr_i[248]), .ZN(n7105) );
  NAND2_X1 U8141 ( .A1(n9438), .A2(pmp_addr_i[249]), .ZN(n7104) );
  OAI21_X1 U8142 ( .B1(n7106), .B2(n7105), .A(n7104), .ZN(n7111) );
  NAND2_X1 U8143 ( .A1(n8807), .A2(pmp_addr_i[250]), .ZN(n7108) );
  NAND2_X1 U8144 ( .A1(n6216), .A2(pmp_addr_i[251]), .ZN(n7107) );
  OAI21_X1 U8145 ( .B1(n7109), .B2(n7108), .A(n7107), .ZN(n7110) );
  AOI21_X1 U8146 ( .B1(n7112), .B2(n7111), .A(n7110), .ZN(n7120) );
  NAND2_X1 U8147 ( .A1(n8814), .A2(pmp_addr_i[252]), .ZN(n7114) );
  NAND2_X1 U8148 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[253]), .ZN(n7113)
         );
  OAI21_X1 U8149 ( .B1(n7115), .B2(n7114), .A(n7113), .ZN(n7117) );
  NOR2_X1 U8150 ( .A1(n7117), .A2(n1703), .ZN(n7118) );
  OAI21_X1 U8151 ( .B1(n7120), .B2(n7119), .A(n7118), .ZN(n7121) );
  NOR2_X1 U8152 ( .A1(n11004), .A2(n7301), .ZN(n7174) );
  NOR2_X1 U8153 ( .A1(data_addr_o_15_), .A2(n7280), .ZN(n7127) );
  NOR2_X1 U8154 ( .A1(n7174), .A2(n7127), .ZN(n7129) );
  NOR2_X1 U8155 ( .A1(n10967), .A2(n430), .ZN(n7177) );
  NAND2_X1 U8156 ( .A1(n8757), .A2(n7175), .ZN(n7285) );
  INV_X1 U8157 ( .A(n7285), .ZN(n7128) );
  NOR2_X1 U8158 ( .A1(n7177), .A2(n7128), .ZN(n7180) );
  NAND2_X1 U8159 ( .A1(n7129), .A2(n7180), .ZN(n7183) );
  INV_X1 U8160 ( .A(n7324), .ZN(n10508) );
  NOR2_X1 U8161 ( .A1(n10508), .A2(n7266), .ZN(n7132) );
  INV_X1 U8162 ( .A(data_addr_i[12]), .ZN(n9947) );
  NOR2_X1 U8163 ( .A1(n31), .A2(n7273), .ZN(n7167) );
  NOR2_X1 U8164 ( .A1(n7132), .A2(n7167), .ZN(n7134) );
  NOR2_X1 U8165 ( .A1(n10847), .A2(n425), .ZN(n7283) );
  NOR2_X1 U8166 ( .A1(n10848), .A2(n7281), .ZN(n7169) );
  NOR2_X1 U8167 ( .A1(n7283), .A2(n7169), .ZN(n7172) );
  NAND2_X1 U8168 ( .A1(n7134), .A2(n7172), .ZN(n7135) );
  NOR2_X1 U8169 ( .A1(n7183), .A2(n7135), .ZN(n7186) );
  OAI22_X1 U8170 ( .A1(n7137), .A2(n10953), .B1(n11255), .B2(n7136), .ZN(n7282) );
  INV_X1 U8171 ( .A(n7282), .ZN(n7150) );
  INV_X1 U8172 ( .A(n7304), .ZN(n7138) );
  OR2_X1 U8173 ( .A1(n10129), .A2(n7138), .ZN(n7141) );
  OR2_X1 U8174 ( .A1(n22), .A2(n7303), .ZN(n7140) );
  AND2_X1 U8175 ( .A1(n22), .A2(n7303), .ZN(n7139) );
  AOI21_X1 U8176 ( .B1(n7141), .B2(n7140), .A(n7139), .ZN(n7144) );
  INV_X1 U8177 ( .A(n12058), .ZN(n10479) );
  NOR2_X1 U8178 ( .A1(n10479), .A2(n7268), .ZN(n7143) );
  NAND2_X1 U8179 ( .A1(n10479), .A2(n7268), .ZN(n11038) );
  OAI21_X1 U8180 ( .B1(n7144), .B2(n7143), .A(n11038), .ZN(n7149) );
  NOR2_X1 U8181 ( .A1(n11331), .A2(n7137), .ZN(n7147) );
  INV_X1 U8182 ( .A(n11291), .ZN(n10486) );
  NAND2_X1 U8183 ( .A1(n10486), .A2(n7136), .ZN(n11033) );
  NAND2_X1 U8184 ( .A1(n11331), .A2(n7137), .ZN(n11056) );
  OAI21_X1 U8185 ( .B1(n7147), .B2(n11033), .A(n11056), .ZN(n7148) );
  AOI21_X1 U8186 ( .B1(n7150), .B2(n7149), .A(n7148), .ZN(n7166) );
  NOR2_X1 U8187 ( .A1(n10494), .A2(n7274), .ZN(n7159) );
  NAND2_X1 U8188 ( .A1(n7152), .A2(n7310), .ZN(n7272) );
  INV_X1 U8189 ( .A(n7272), .ZN(n7153) );
  NOR2_X1 U8190 ( .A1(n7159), .A2(n7153), .ZN(n7157) );
  INV_X1 U8191 ( .A(n10501), .ZN(n10504) );
  NOR2_X1 U8192 ( .A1(n10504), .A2(n7275), .ZN(n7156) );
  NOR2_X1 U8193 ( .A1(n10838), .A2(n7265), .ZN(n7160) );
  NOR2_X1 U8194 ( .A1(n7156), .A2(n7160), .ZN(n7163) );
  NAND2_X1 U8195 ( .A1(n7157), .A2(n7163), .ZN(n7165) );
  INV_X1 U8196 ( .A(n7152), .ZN(n10493) );
  NAND2_X1 U8197 ( .A1(n10493), .A2(n477), .ZN(n7158) );
  NAND2_X1 U8198 ( .A1(n10494), .A2(n7274), .ZN(n11067) );
  OAI21_X1 U8199 ( .B1(n7159), .B2(n7158), .A(n11067), .ZN(n7162) );
  NAND2_X1 U8200 ( .A1(n10504), .A2(n7275), .ZN(n11064) );
  NAND2_X1 U8201 ( .A1(n10838), .A2(n7265), .ZN(n11069) );
  OAI21_X1 U8202 ( .B1(n7160), .B2(n11064), .A(n11069), .ZN(n7161) );
  AOI21_X1 U8203 ( .B1(n7163), .B2(n7162), .A(n7161), .ZN(n7164) );
  OAI21_X1 U8204 ( .B1(n7166), .B2(n7165), .A(n7164), .ZN(n7185) );
  NAND2_X1 U8205 ( .A1(n10508), .A2(n7266), .ZN(n11065) );
  NAND2_X1 U8206 ( .A1(n31), .A2(n7273), .ZN(n11042) );
  OAI21_X1 U8207 ( .B1(n7167), .B2(n11065), .A(n11042), .ZN(n7171) );
  NAND2_X1 U8208 ( .A1(n10847), .A2(n425), .ZN(n11059) );
  NAND2_X1 U8209 ( .A1(n10848), .A2(n7281), .ZN(n7168) );
  OAI21_X1 U8210 ( .B1(n7169), .B2(n11059), .A(n7168), .ZN(n7170) );
  AOI21_X1 U8211 ( .B1(n7172), .B2(n7171), .A(n7170), .ZN(n7182) );
  NAND2_X1 U8212 ( .A1(data_addr_o_15_), .A2(n7280), .ZN(n11074) );
  NAND2_X1 U8213 ( .A1(n11004), .A2(n7301), .ZN(n7173) );
  OAI21_X1 U8214 ( .B1(n7174), .B2(n11074), .A(n7173), .ZN(n7179) );
  NAND2_X1 U8215 ( .A1(data_addr_o_17_), .A2(n439), .ZN(n11030) );
  NAND2_X1 U8216 ( .A1(n11298), .A2(n430), .ZN(n7176) );
  OAI21_X1 U8217 ( .B1(n7177), .B2(n11030), .A(n7176), .ZN(n7178) );
  AOI21_X1 U8218 ( .B1(n7180), .B2(n7179), .A(n7178), .ZN(n7181) );
  OAI21_X1 U8219 ( .B1(n7183), .B2(n7182), .A(n7181), .ZN(n7184) );
  AOI21_X1 U8220 ( .B1(n7186), .B2(n7185), .A(n7184), .ZN(n7244) );
  INV_X1 U8221 ( .A(n7249), .ZN(n7211) );
  NOR2_X1 U8222 ( .A1(data_addr_o_23_), .A2(n7211), .ZN(n7187) );
  NOR2_X1 U8223 ( .A1(n10738), .A2(n356), .ZN(n7214) );
  NOR2_X1 U8224 ( .A1(n7187), .A2(n7214), .ZN(n7189) );
  NOR2_X1 U8225 ( .A1(n10903), .A2(n391), .ZN(n7188) );
  NOR2_X1 U8226 ( .A1(n10267), .A2(n353), .ZN(n7217) );
  NOR2_X1 U8227 ( .A1(n7188), .A2(n7217), .ZN(n7220) );
  NAND2_X1 U8228 ( .A1(n7189), .A2(n7220), .ZN(n7222) );
  NOR2_X1 U8229 ( .A1(n10202), .A2(n365), .ZN(n7190) );
  NOR2_X1 U8230 ( .A1(n9529), .A2(n358), .ZN(n7207) );
  NOR2_X1 U8231 ( .A1(n7190), .A2(n7207), .ZN(n7210) );
  INV_X1 U8232 ( .A(n7248), .ZN(n7201) );
  NOR2_X1 U8233 ( .A1(n9846), .A2(n7201), .ZN(n7191) );
  BUF_X1 U8234 ( .A(data_addr_i[20]), .Z(n11285) );
  NOR2_X1 U8235 ( .A1(n11285), .A2(n5347), .ZN(n7204) );
  NOR2_X1 U8236 ( .A1(n7191), .A2(n7204), .ZN(n7192) );
  NAND2_X1 U8237 ( .A1(n7210), .A2(n7192), .ZN(n7193) );
  NOR2_X1 U8238 ( .A1(n7222), .A2(n7193), .ZN(n7200) );
  NOR2_X1 U8239 ( .A1(n9886), .A2(n371), .ZN(n7194) );
  NOR2_X1 U8240 ( .A1(n10635), .A2(n347), .ZN(n7226) );
  NOR2_X1 U8241 ( .A1(n7194), .A2(n7226), .ZN(n7196) );
  NOR2_X1 U8242 ( .A1(n9955), .A2(n375), .ZN(n7195) );
  NOR2_X1 U8243 ( .A1(n10919), .A2(n343), .ZN(n7229) );
  NOR2_X1 U8244 ( .A1(n7195), .A2(n7229), .ZN(n7232) );
  NAND2_X1 U8245 ( .A1(n7196), .A2(n7232), .ZN(n7199) );
  NOR2_X1 U8246 ( .A1(n10662), .A2(n398), .ZN(n7197) );
  NOR2_X1 U8247 ( .A1(n7197), .A2(pmp_addr_i[222]), .ZN(n7198) );
  INV_X1 U8248 ( .A(pmp_addr_i[223]), .ZN(n7234) );
  NAND2_X1 U8249 ( .A1(n7198), .A2(n7234), .ZN(n7237) );
  NOR2_X1 U8250 ( .A1(n7199), .A2(n7237), .ZN(n7240) );
  NAND2_X1 U8251 ( .A1(n7200), .A2(n7240), .ZN(n7243) );
  NAND2_X1 U8252 ( .A1(n9846), .A2(n7201), .ZN(n7203) );
  NAND2_X1 U8253 ( .A1(n11285), .A2(n5347), .ZN(n7202) );
  OAI21_X1 U8254 ( .B1(n7204), .B2(n7203), .A(n7202), .ZN(n7209) );
  NAND2_X1 U8255 ( .A1(n10202), .A2(n365), .ZN(n7206) );
  NAND2_X1 U8256 ( .A1(n9529), .A2(n358), .ZN(n7205) );
  OAI21_X1 U8257 ( .B1(n7207), .B2(n7206), .A(n7205), .ZN(n7208) );
  AOI21_X1 U8258 ( .B1(n7210), .B2(n7209), .A(n7208), .ZN(n7223) );
  NAND2_X1 U8259 ( .A1(data_addr_o_23_), .A2(n7211), .ZN(n7213) );
  NAND2_X1 U8260 ( .A1(n10629), .A2(n356), .ZN(n7212) );
  OAI21_X1 U8261 ( .B1(n7214), .B2(n7213), .A(n7212), .ZN(n7219) );
  NAND2_X1 U8262 ( .A1(n10903), .A2(n391), .ZN(n7216) );
  NAND2_X1 U8263 ( .A1(n10267), .A2(n353), .ZN(n7215) );
  OAI21_X1 U8264 ( .B1(n7217), .B2(n7216), .A(n7215), .ZN(n7218) );
  AOI21_X1 U8265 ( .B1(n7220), .B2(n7219), .A(n7218), .ZN(n7221) );
  OAI21_X1 U8266 ( .B1(n7223), .B2(n7222), .A(n7221), .ZN(n7241) );
  NAND2_X1 U8267 ( .A1(n9886), .A2(n371), .ZN(n7225) );
  NAND2_X1 U8268 ( .A1(n10914), .A2(n347), .ZN(n7224) );
  OAI21_X1 U8269 ( .B1(n7226), .B2(n7225), .A(n7224), .ZN(n7231) );
  NAND2_X1 U8270 ( .A1(n9955), .A2(n375), .ZN(n7228) );
  NAND2_X1 U8271 ( .A1(n10919), .A2(n343), .ZN(n7227) );
  OAI21_X1 U8272 ( .B1(n7229), .B2(n7228), .A(n7227), .ZN(n7230) );
  AOI21_X1 U8273 ( .B1(n7232), .B2(n7231), .A(n7230), .ZN(n7238) );
  NAND2_X1 U8274 ( .A1(n12123), .A2(n398), .ZN(n7233) );
  NOR2_X1 U8275 ( .A1(n7233), .A2(pmp_addr_i[222]), .ZN(n7235) );
  NAND2_X1 U8276 ( .A1(n7235), .A2(n7234), .ZN(n7236) );
  OAI21_X1 U8277 ( .B1(n7238), .B2(n7237), .A(n7236), .ZN(n7239) );
  AOI21_X1 U8278 ( .B1(n7241), .B2(n7240), .A(n7239), .ZN(n7242) );
  OAI21_X1 U8279 ( .B1(n7244), .B2(n7243), .A(n7242), .ZN(n7245) );
  XNOR2_X1 U8280 ( .A(data_addr_o_30_), .B(n7247), .ZN(n7254) );
  XNOR2_X1 U8281 ( .A(n10627), .B(n7248), .ZN(n7253) );
  XNOR2_X1 U8282 ( .A(data_addr_o_23_), .B(n7249), .ZN(n7252) );
  XNOR2_X1 U8283 ( .A(n10629), .B(n7250), .ZN(n7251) );
  NAND4_X1 U8284 ( .A1(n7254), .A2(n7253), .A3(n7252), .A4(n7251), .ZN(n7264)
         );
  XNOR2_X1 U8285 ( .A(n10616), .B(n7255), .ZN(n7262) );
  XNOR2_X1 U8286 ( .A(n11285), .B(n7256), .ZN(n7261) );
  XNOR2_X1 U8287 ( .A(n10614), .B(n7257), .ZN(n7260) );
  XNOR2_X1 U8288 ( .A(n10606), .B(n7258), .ZN(n7259) );
  NAND4_X1 U8289 ( .A1(n7262), .A2(n7261), .A3(n7260), .A4(n7259), .ZN(n7263)
         );
  NOR2_X1 U8290 ( .A1(n7264), .A2(n7263), .ZN(n7300) );
  OAI22_X1 U8291 ( .A1(n7266), .A2(data_addr_o_11_), .B1(n11343), .B2(n7265), 
        .ZN(n7278) );
  INV_X1 U8292 ( .A(n7267), .ZN(n7303) );
  OAI22_X1 U8293 ( .A1(n11288), .A2(n7268), .B1(n10818), .B2(n7303), .ZN(n7270) );
  OAI21_X1 U8294 ( .B1(data_addr_o_2_), .B2(n7138), .A(pmp_cfg_i[60]), .ZN(
        n7269) );
  NOR2_X1 U8295 ( .A1(n7270), .A2(n7269), .ZN(n7271) );
  OAI211_X1 U8296 ( .C1(n7273), .C2(data_addr_o_12_), .A(n7272), .B(n7271), 
        .ZN(n7277) );
  OAI22_X1 U8297 ( .A1(data_addr_o_9_), .A2(n7275), .B1(n10281), .B2(n7274), 
        .ZN(n7276) );
  NOR3_X1 U8298 ( .A1(n7278), .A2(n7277), .A3(n7276), .ZN(n7288) );
  XNOR2_X1 U8299 ( .A(n10967), .B(n7279), .ZN(n7287) );
  OAI22_X1 U8300 ( .A1(n7281), .A2(data_addr_o_14_), .B1(data_addr_o_15_), 
        .B2(n7280), .ZN(n7284) );
  NOR3_X1 U8301 ( .A1(n7284), .A2(n7283), .A3(n7282), .ZN(n7286) );
  NAND4_X1 U8302 ( .A1(n7288), .A2(n7287), .A3(n7286), .A4(n7285), .ZN(n7294)
         );
  XNOR2_X1 U8303 ( .A(n10638), .B(n7289), .ZN(n7292) );
  XNOR2_X1 U8304 ( .A(n9955), .B(n7290), .ZN(n7291) );
  NAND2_X1 U8305 ( .A1(n7292), .A2(n7291), .ZN(n7293) );
  NOR2_X1 U8306 ( .A1(n7294), .A2(n7293), .ZN(n7299) );
  XNOR2_X1 U8307 ( .A(n10635), .B(n7295), .ZN(n7298) );
  XNOR2_X1 U8308 ( .A(n10612), .B(n7296), .ZN(n7297) );
  NAND4_X1 U8309 ( .A1(n7300), .A2(n7299), .A3(n7298), .A4(n7297), .ZN(n11082)
         );
  XNOR2_X1 U8310 ( .A(n9987), .B(n7301), .ZN(n7308) );
  OAI21_X1 U8311 ( .B1(n11334), .B2(n7302), .A(n11074), .ZN(n11076) );
  INV_X1 U8312 ( .A(data_addr_i[2]), .ZN(n8695) );
  NAND2_X1 U8313 ( .A1(data_addr_o_3_), .A2(n7303), .ZN(n11034) );
  OAI211_X1 U8314 ( .C1(n7304), .C2(n8695), .A(n11038), .B(n11034), .ZN(n7305)
         );
  INV_X1 U8315 ( .A(n7305), .ZN(n7306) );
  NAND3_X1 U8316 ( .A1(n11059), .A2(n7306), .A3(n11033), .ZN(n7307) );
  NOR3_X1 U8317 ( .A1(n7308), .A2(n11076), .A3(n7307), .ZN(n7315) );
  XNOR2_X1 U8318 ( .A(n12123), .B(n7309), .ZN(n7314) );
  NAND3_X1 U8319 ( .A1(n11064), .A2(n11042), .A3(n11056), .ZN(n7312) );
  NAND2_X1 U8320 ( .A1(n11069), .A2(n11065), .ZN(n7311) );
  OAI21_X1 U8321 ( .B1(n6400), .B2(n7310), .A(n11067), .ZN(n11032) );
  NOR3_X1 U8322 ( .A1(n7312), .A2(n7311), .A3(n11032), .ZN(n7313) );
  NAND4_X1 U8323 ( .A1(n7315), .A2(n7314), .A3(n7313), .A4(n11030), .ZN(n7316)
         );
  MUX2_X1 U8324 ( .A(pmp_cfg_i[56]), .B(pmp_cfg_i[57]), .S(n11019), .Z(n7318)
         );
  AND2_X1 U8325 ( .A1(n7317), .A2(n7318), .ZN(n11047) );
  NAND2_X1 U8326 ( .A1(n7319), .A2(n11047), .ZN(n8086) );
  NOR2_X1 U8327 ( .A1(n10335), .A2(n7556), .ZN(n7368) );
  NAND2_X1 U8328 ( .A1(n9941), .A2(n7367), .ZN(n7554) );
  INV_X1 U8329 ( .A(n7554), .ZN(n7321) );
  NOR2_X1 U8330 ( .A1(n7368), .A2(n7321), .ZN(n7323) );
  NOR2_X1 U8331 ( .A1(n11298), .A2(n4252), .ZN(n7371) );
  NOR2_X1 U8332 ( .A1(data_addr_o_17_), .A2(n4251), .ZN(n7570) );
  NOR2_X1 U8333 ( .A1(n7371), .A2(n7570), .ZN(n7374) );
  NAND2_X1 U8334 ( .A1(n7323), .A2(n7374), .ZN(n7377) );
  INV_X1 U8335 ( .A(n7325), .ZN(n7360) );
  NOR2_X1 U8336 ( .A1(data_addr_o_11_), .A2(n7360), .ZN(n7327) );
  NOR2_X1 U8337 ( .A1(data_addr_o_12_), .A2(n4242), .ZN(n7361) );
  NOR2_X1 U8338 ( .A1(n7327), .A2(n7361), .ZN(n7330) );
  NOR2_X1 U8339 ( .A1(n10847), .A2(n7564), .ZN(n7329) );
  NAND2_X1 U8340 ( .A1(n11334), .A2(n7362), .ZN(n7555) );
  INV_X1 U8341 ( .A(n7555), .ZN(n7363) );
  NOR2_X1 U8342 ( .A1(n7329), .A2(n7363), .ZN(n7366) );
  NAND2_X1 U8343 ( .A1(n7330), .A2(n7366), .ZN(n7331) );
  NOR2_X1 U8344 ( .A1(n7377), .A2(n7331), .ZN(n7380) );
  NOR2_X1 U8345 ( .A1(n10824), .A2(n4182), .ZN(n7334) );
  NOR2_X1 U8346 ( .A1(n11331), .A2(n7563), .ZN(n7341) );
  NOR2_X1 U8347 ( .A1(n7334), .A2(n7341), .ZN(n7344) );
  OR2_X1 U8348 ( .A1(data_addr_o_2_), .A2(n157), .ZN(n7338) );
  INV_X1 U8349 ( .A(n10473), .ZN(n10818) );
  OR2_X1 U8350 ( .A1(n10818), .A2(n7606), .ZN(n7337) );
  AND2_X1 U8351 ( .A1(n10818), .A2(n7606), .ZN(n7336) );
  AOI21_X1 U8352 ( .B1(n7338), .B2(n7337), .A(n7336), .ZN(n7340) );
  NOR2_X1 U8353 ( .A1(n10135), .A2(n4816), .ZN(n7339) );
  NAND2_X1 U8354 ( .A1(n10479), .A2(n4816), .ZN(n11726) );
  OAI21_X1 U8355 ( .B1(n7340), .B2(n7339), .A(n11726), .ZN(n7343) );
  NAND2_X1 U8356 ( .A1(n10824), .A2(n4182), .ZN(n11725) );
  NAND2_X1 U8357 ( .A1(data_addr_o_6_), .A2(n7563), .ZN(n11732) );
  OAI21_X1 U8358 ( .B1(n7341), .B2(n11725), .A(n11732), .ZN(n7342) );
  AOI21_X1 U8359 ( .B1(n7344), .B2(n7343), .A(n7342), .ZN(n7359) );
  NOR2_X1 U8360 ( .A1(n8237), .A2(n4203), .ZN(n7347) );
  NOR2_X1 U8361 ( .A1(n8238), .A2(n4205), .ZN(n7353) );
  NOR2_X1 U8362 ( .A1(n7347), .A2(n7353), .ZN(n7356) );
  INV_X1 U8363 ( .A(n7814), .ZN(n10836) );
  NOR2_X1 U8364 ( .A1(n10836), .A2(n4201), .ZN(n7352) );
  NOR2_X1 U8365 ( .A1(n7816), .A2(n7557), .ZN(n7350) );
  NOR2_X1 U8366 ( .A1(n7352), .A2(n7350), .ZN(n7351) );
  NAND2_X1 U8367 ( .A1(n7356), .A2(n7351), .ZN(n7358) );
  NAND2_X1 U8368 ( .A1(n7816), .A2(n7557), .ZN(n11748) );
  NAND2_X1 U8369 ( .A1(n10836), .A2(n4201), .ZN(n11723) );
  OAI21_X1 U8370 ( .B1(n7352), .B2(n11748), .A(n11723), .ZN(n7355) );
  NAND2_X1 U8371 ( .A1(data_addr_o_9_), .A2(n4203), .ZN(n11747) );
  NAND2_X1 U8372 ( .A1(n8238), .A2(n4205), .ZN(n11745) );
  OAI21_X1 U8373 ( .B1(n7353), .B2(n11747), .A(n11745), .ZN(n7354) );
  AOI21_X1 U8374 ( .B1(n7356), .B2(n7355), .A(n7354), .ZN(n7357) );
  OAI21_X1 U8375 ( .B1(n7359), .B2(n7358), .A(n7357), .ZN(n7379) );
  NAND2_X1 U8376 ( .A1(n10508), .A2(n7360), .ZN(n11724) );
  NAND2_X1 U8377 ( .A1(data_addr_o_12_), .A2(n4242), .ZN(n11712) );
  OAI21_X1 U8378 ( .B1(n7361), .B2(n11724), .A(n11712), .ZN(n7365) );
  NAND2_X1 U8379 ( .A1(n10847), .A2(n7564), .ZN(n11709) );
  NAND2_X1 U8380 ( .A1(n10848), .A2(n4807), .ZN(n11699) );
  OAI21_X1 U8381 ( .B1(n7363), .B2(n11709), .A(n11699), .ZN(n7364) );
  AOI21_X1 U8382 ( .B1(n7366), .B2(n7365), .A(n7364), .ZN(n7376) );
  NAND2_X1 U8383 ( .A1(n10657), .A2(n4810), .ZN(n11700) );
  NAND2_X1 U8384 ( .A1(n10335), .A2(n7556), .ZN(n11719) );
  OAI21_X1 U8385 ( .B1(n7368), .B2(n11700), .A(n11719), .ZN(n7373) );
  NAND2_X1 U8386 ( .A1(n6813), .A2(n4251), .ZN(n7370) );
  NAND2_X1 U8387 ( .A1(n10967), .A2(n4252), .ZN(n7369) );
  OAI21_X1 U8388 ( .B1(n7371), .B2(n7370), .A(n7369), .ZN(n7372) );
  AOI21_X1 U8389 ( .B1(n7374), .B2(n7373), .A(n7372), .ZN(n7375) );
  OAI21_X1 U8390 ( .B1(n7377), .B2(n7376), .A(n7375), .ZN(n7378) );
  AOI21_X1 U8391 ( .B1(n7380), .B2(n7379), .A(n7378), .ZN(n7436) );
  NOR2_X1 U8392 ( .A1(n10898), .A2(n4340), .ZN(n7381) );
  NOR2_X1 U8393 ( .A1(n10738), .A2(n4341), .ZN(n7407) );
  NOR2_X1 U8394 ( .A1(n7381), .A2(n7407), .ZN(n7383) );
  NOR2_X1 U8395 ( .A1(n9923), .A2(n4345), .ZN(n7382) );
  NOR2_X1 U8396 ( .A1(n10904), .A2(n4346), .ZN(n7410) );
  NOR2_X1 U8397 ( .A1(n7382), .A2(n7410), .ZN(n7413) );
  NAND2_X1 U8398 ( .A1(n7383), .A2(n7413), .ZN(n7415) );
  NOR2_X1 U8399 ( .A1(n10202), .A2(n4332), .ZN(n7384) );
  NOR2_X1 U8400 ( .A1(n9915), .A2(n4333), .ZN(n7401) );
  NOR2_X1 U8401 ( .A1(n7384), .A2(n7401), .ZN(n7404) );
  NOR2_X1 U8402 ( .A1(n9846), .A2(n4327), .ZN(n7386) );
  NOR2_X1 U8403 ( .A1(data_addr_o_20_), .A2(n4328), .ZN(n7398) );
  NOR2_X1 U8404 ( .A1(n7386), .A2(n7398), .ZN(n7387) );
  NAND2_X1 U8405 ( .A1(n7404), .A2(n7387), .ZN(n7388) );
  NOR2_X1 U8406 ( .A1(n7415), .A2(n7388), .ZN(n7395) );
  NOR2_X1 U8407 ( .A1(n9886), .A2(n4307), .ZN(n7389) );
  NOR2_X1 U8408 ( .A1(n10914), .A2(n4308), .ZN(n7419) );
  NOR2_X1 U8409 ( .A1(n7389), .A2(n7419), .ZN(n7391) );
  NOR2_X1 U8410 ( .A1(n9955), .A2(n4312), .ZN(n7390) );
  NOR2_X1 U8411 ( .A1(n10919), .A2(n4313), .ZN(n7422) );
  NOR2_X1 U8412 ( .A1(n7390), .A2(n7422), .ZN(n7425) );
  NAND2_X1 U8413 ( .A1(n7391), .A2(n7425), .ZN(n7394) );
  NOR2_X1 U8414 ( .A1(n10662), .A2(n4320), .ZN(n7392) );
  NOR2_X1 U8415 ( .A1(n7392), .A2(pmp_addr_i[94]), .ZN(n7393) );
  NAND2_X1 U8416 ( .A1(n7393), .A2(n4303), .ZN(n7429) );
  NOR2_X1 U8417 ( .A1(n7394), .A2(n7429), .ZN(n7432) );
  NAND2_X1 U8418 ( .A1(n7395), .A2(n7432), .ZN(n7435) );
  NAND2_X1 U8419 ( .A1(n9846), .A2(n4327), .ZN(n7397) );
  NAND2_X1 U8420 ( .A1(n10887), .A2(n4328), .ZN(n7396) );
  OAI21_X1 U8421 ( .B1(n7398), .B2(n7397), .A(n7396), .ZN(n7403) );
  NAND2_X1 U8422 ( .A1(n10202), .A2(n4332), .ZN(n7400) );
  NAND2_X1 U8423 ( .A1(n9915), .A2(n4333), .ZN(n7399) );
  OAI21_X1 U8424 ( .B1(n7401), .B2(n7400), .A(n7399), .ZN(n7402) );
  AOI21_X1 U8425 ( .B1(n7404), .B2(n7403), .A(n7402), .ZN(n7416) );
  NAND2_X1 U8426 ( .A1(n10898), .A2(n4340), .ZN(n7406) );
  NAND2_X1 U8427 ( .A1(n10738), .A2(n4341), .ZN(n7405) );
  OAI21_X1 U8428 ( .B1(n7407), .B2(n7406), .A(n7405), .ZN(n7412) );
  NAND2_X1 U8429 ( .A1(n9923), .A2(n4345), .ZN(n7409) );
  NAND2_X1 U8430 ( .A1(n10904), .A2(n4346), .ZN(n7408) );
  OAI21_X1 U8431 ( .B1(n7410), .B2(n7409), .A(n7408), .ZN(n7411) );
  AOI21_X1 U8432 ( .B1(n7413), .B2(n7412), .A(n7411), .ZN(n7414) );
  OAI21_X1 U8433 ( .B1(n7416), .B2(n7415), .A(n7414), .ZN(n7433) );
  NAND2_X1 U8434 ( .A1(n9886), .A2(n4307), .ZN(n7418) );
  NAND2_X1 U8435 ( .A1(n10914), .A2(n4308), .ZN(n7417) );
  OAI21_X1 U8436 ( .B1(n7419), .B2(n7418), .A(n7417), .ZN(n7424) );
  NAND2_X1 U8437 ( .A1(n9955), .A2(n4312), .ZN(n7421) );
  NAND2_X1 U8438 ( .A1(n10919), .A2(n4313), .ZN(n7420) );
  OAI21_X1 U8439 ( .B1(n7422), .B2(n7421), .A(n7420), .ZN(n7423) );
  AOI21_X1 U8440 ( .B1(n7425), .B2(n7424), .A(n7423), .ZN(n7430) );
  NAND2_X1 U8441 ( .A1(n12123), .A2(n4320), .ZN(n7426) );
  NOR2_X1 U8442 ( .A1(n7426), .A2(pmp_addr_i[94]), .ZN(n7427) );
  NAND2_X1 U8443 ( .A1(n7427), .A2(n4303), .ZN(n7428) );
  OAI21_X1 U8444 ( .B1(n7430), .B2(n7429), .A(n7428), .ZN(n7431) );
  AOI21_X1 U8445 ( .B1(n7433), .B2(n7432), .A(n7431), .ZN(n7434) );
  OAI21_X1 U8446 ( .B1(n7436), .B2(n7435), .A(n7434), .ZN(n7553) );
  INV_X1 U8447 ( .A(data_addr_o_16_), .ZN(n7482) );
  NOR2_X1 U8448 ( .A1(n7482), .A2(pmp_addr_i[110]), .ZN(n7485) );
  NOR2_X1 U8449 ( .A1(n10721), .A2(pmp_addr_i[109]), .ZN(n7437) );
  NOR2_X1 U8450 ( .A1(n7485), .A2(n7437), .ZN(n7439) );
  NOR2_X1 U8451 ( .A1(n12184), .A2(pmp_addr_i[112]), .ZN(n7488) );
  NOR2_X1 U8452 ( .A1(n8757), .A2(pmp_addr_i[111]), .ZN(n7438) );
  NOR2_X1 U8453 ( .A1(n7488), .A2(n7438), .ZN(n7490) );
  NAND2_X1 U8454 ( .A1(n7439), .A2(n7490), .ZN(n7493) );
  NOR2_X1 U8455 ( .A1(n9508), .A2(pmp_addr_i[105]), .ZN(n7440) );
  INV_X1 U8456 ( .A(n10499), .ZN(n7472) );
  NOR2_X1 U8457 ( .A1(n7472), .A2(pmp_addr_i[106]), .ZN(n7475) );
  NOR2_X1 U8458 ( .A1(n7440), .A2(n7475), .ZN(n7442) );
  NOR2_X1 U8459 ( .A1(n10342), .A2(pmp_addr_i[107]), .ZN(n7441) );
  NOR2_X1 U8460 ( .A1(n11334), .A2(pmp_addr_i[108]), .ZN(n7478) );
  NOR2_X1 U8461 ( .A1(n7441), .A2(n7478), .ZN(n7481) );
  NAND2_X1 U8462 ( .A1(n7442), .A2(n7481), .ZN(n7443) );
  NOR2_X1 U8463 ( .A1(n7493), .A2(n7443), .ZN(n7496) );
  OR2_X1 U8464 ( .A1(pmp_addr_i[97]), .A2(n10010), .ZN(n7446) );
  AND2_X1 U8465 ( .A1(pmp_addr_i[96]), .A2(n10651), .ZN(n7445) );
  AND2_X1 U8466 ( .A1(pmp_addr_i[97]), .A2(n10010), .ZN(n7444) );
  AOI21_X1 U8467 ( .B1(n7446), .B2(n7445), .A(n7444), .ZN(n7449) );
  NOR2_X1 U8468 ( .A1(pmp_addr_i[98]), .A2(n8406), .ZN(n7448) );
  NAND2_X1 U8469 ( .A1(pmp_addr_i[98]), .A2(n6123), .ZN(n7447) );
  OAI21_X1 U8470 ( .B1(n7449), .B2(n7448), .A(n7447), .ZN(n7456) );
  NOR2_X1 U8471 ( .A1(n6127), .A2(pmp_addr_i[99]), .ZN(n7450) );
  NOR2_X1 U8472 ( .A1(n8410), .A2(pmp_addr_i[100]), .ZN(n7453) );
  NOR2_X1 U8473 ( .A1(n7450), .A2(n7453), .ZN(n7455) );
  NAND2_X1 U8474 ( .A1(n6127), .A2(pmp_addr_i[99]), .ZN(n7452) );
  NAND2_X1 U8475 ( .A1(n10362), .A2(pmp_addr_i[100]), .ZN(n7451) );
  OAI21_X1 U8476 ( .B1(n7453), .B2(n7452), .A(n7451), .ZN(n7454) );
  AOI21_X1 U8477 ( .B1(n7456), .B2(n7455), .A(n7454), .ZN(n7471) );
  NOR2_X1 U8478 ( .A1(n29), .A2(pmp_addr_i[102]), .ZN(n7462) );
  NOR2_X1 U8479 ( .A1(n10697), .A2(pmp_addr_i[101]), .ZN(n7457) );
  NOR2_X1 U8480 ( .A1(n7462), .A2(n7457), .ZN(n7459) );
  NOR2_X1 U8481 ( .A1(n10501), .A2(pmp_addr_i[103]), .ZN(n7458) );
  NOR2_X1 U8482 ( .A1(n7964), .A2(pmp_addr_i[104]), .ZN(n7465) );
  NOR2_X1 U8483 ( .A1(n7458), .A2(n7465), .ZN(n7468) );
  NAND2_X1 U8484 ( .A1(n7459), .A2(n7468), .ZN(n7470) );
  NAND2_X1 U8485 ( .A1(n10697), .A2(pmp_addr_i[101]), .ZN(n7461) );
  NAND2_X1 U8486 ( .A1(n8735), .A2(pmp_addr_i[102]), .ZN(n7460) );
  OAI21_X1 U8487 ( .B1(n7462), .B2(n7461), .A(n7460), .ZN(n7467) );
  NAND2_X1 U8488 ( .A1(n10501), .A2(pmp_addr_i[103]), .ZN(n7464) );
  NAND2_X1 U8489 ( .A1(n6141), .A2(pmp_addr_i[104]), .ZN(n7463) );
  OAI21_X1 U8490 ( .B1(n7465), .B2(n7464), .A(n7463), .ZN(n7466) );
  AOI21_X1 U8491 ( .B1(n7468), .B2(n7467), .A(n7466), .ZN(n7469) );
  OAI21_X1 U8492 ( .B1(n7471), .B2(n7470), .A(n7469), .ZN(n7495) );
  NAND2_X1 U8493 ( .A1(n7324), .A2(pmp_addr_i[105]), .ZN(n7474) );
  NAND2_X1 U8494 ( .A1(n7472), .A2(pmp_addr_i[106]), .ZN(n7473) );
  OAI21_X1 U8495 ( .B1(n7475), .B2(n7474), .A(n7473), .ZN(n7480) );
  NAND2_X1 U8496 ( .A1(n11006), .A2(pmp_addr_i[107]), .ZN(n7477) );
  NAND2_X1 U8497 ( .A1(n6154), .A2(pmp_addr_i[108]), .ZN(n7476) );
  OAI21_X1 U8498 ( .B1(n7478), .B2(n7477), .A(n7476), .ZN(n7479) );
  AOI21_X1 U8499 ( .B1(n7481), .B2(n7480), .A(n7479), .ZN(n7492) );
  NAND2_X1 U8500 ( .A1(n10721), .A2(pmp_addr_i[109]), .ZN(n7484) );
  NAND2_X1 U8501 ( .A1(n7482), .A2(pmp_addr_i[110]), .ZN(n7483) );
  OAI21_X1 U8502 ( .B1(n7485), .B2(n7484), .A(n7483), .ZN(n7491) );
  NAND2_X1 U8503 ( .A1(n8444), .A2(pmp_addr_i[111]), .ZN(n7487) );
  NAND2_X1 U8504 ( .A1(n10060), .A2(pmp_addr_i[112]), .ZN(n7486) );
  OAI21_X1 U8505 ( .B1(n7488), .B2(n7487), .A(n7486), .ZN(n7489) );
  AOI21_X1 U8506 ( .B1(n7496), .B2(n7495), .A(n7494), .ZN(n7550) );
  NOR2_X1 U8507 ( .A1(n10424), .A2(pmp_addr_i[117]), .ZN(n7497) );
  NOR2_X1 U8508 ( .A1(n9163), .A2(pmp_addr_i[118]), .ZN(n7520) );
  NOR2_X1 U8509 ( .A1(n7497), .A2(n7520), .ZN(n7499) );
  NOR2_X1 U8510 ( .A1(n10429), .A2(pmp_addr_i[119]), .ZN(n7498) );
  NOR2_X1 U8511 ( .A1(n10439), .A2(pmp_addr_i[120]), .ZN(n7523) );
  NOR2_X1 U8512 ( .A1(n7498), .A2(n7523), .ZN(n7526) );
  NAND2_X1 U8513 ( .A1(n7499), .A2(n7526), .ZN(n7528) );
  NOR2_X1 U8514 ( .A1(n9418), .A2(pmp_addr_i[115]), .ZN(n7500) );
  NOR2_X1 U8515 ( .A1(n9156), .A2(pmp_addr_i[116]), .ZN(n7514) );
  NOR2_X1 U8516 ( .A1(n7500), .A2(n7514), .ZN(n7517) );
  NOR2_X1 U8517 ( .A1(n9414), .A2(pmp_addr_i[113]), .ZN(n7501) );
  NOR2_X1 U8518 ( .A1(n6188), .A2(pmp_addr_i[114]), .ZN(n7511) );
  NOR2_X1 U8519 ( .A1(n7501), .A2(n7511), .ZN(n7502) );
  NAND2_X1 U8520 ( .A1(n7517), .A2(n7502), .ZN(n7503) );
  NOR2_X1 U8521 ( .A1(n7528), .A2(n7503), .ZN(n7508) );
  NOR2_X1 U8522 ( .A1(n9438), .A2(pmp_addr_i[121]), .ZN(n7504) );
  NOR2_X1 U8523 ( .A1(n10443), .A2(pmp_addr_i[122]), .ZN(n7532) );
  NOR2_X1 U8524 ( .A1(n7504), .A2(n7532), .ZN(n7506) );
  NOR2_X1 U8525 ( .A1(n6216), .A2(pmp_addr_i[123]), .ZN(n7505) );
  NOR2_X1 U8526 ( .A1(n8494), .A2(pmp_addr_i[124]), .ZN(n7535) );
  NOR2_X1 U8527 ( .A1(n7505), .A2(n7535), .ZN(n7538) );
  NAND2_X1 U8528 ( .A1(n7506), .A2(n7538), .ZN(n7507) );
  NOR2_X1 U8529 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[125]), .ZN(n7543)
         );
  NOR2_X1 U8530 ( .A1(n7507), .A2(n7543), .ZN(n7546) );
  NAND2_X1 U8531 ( .A1(n7508), .A2(n7546), .ZN(n7549) );
  NAND2_X1 U8532 ( .A1(n10414), .A2(pmp_addr_i[113]), .ZN(n7510) );
  NAND2_X1 U8533 ( .A1(n10754), .A2(pmp_addr_i[114]), .ZN(n7509) );
  OAI21_X1 U8534 ( .B1(n7511), .B2(n7510), .A(n7509), .ZN(n7516) );
  NAND2_X1 U8535 ( .A1(n9418), .A2(pmp_addr_i[115]), .ZN(n7513) );
  NAND2_X1 U8536 ( .A1(n9425), .A2(pmp_addr_i[116]), .ZN(n7512) );
  OAI21_X1 U8537 ( .B1(n7514), .B2(n7513), .A(n7512), .ZN(n7515) );
  AOI21_X1 U8538 ( .B1(n7517), .B2(n7516), .A(n7515), .ZN(n7529) );
  NAND2_X1 U8539 ( .A1(n10424), .A2(pmp_addr_i[117]), .ZN(n7519) );
  NAND2_X1 U8540 ( .A1(n10428), .A2(pmp_addr_i[118]), .ZN(n7518) );
  OAI21_X1 U8541 ( .B1(n7520), .B2(n7519), .A(n7518), .ZN(n7525) );
  NAND2_X1 U8542 ( .A1(n10429), .A2(pmp_addr_i[119]), .ZN(n7522) );
  NAND2_X1 U8543 ( .A1(n10439), .A2(pmp_addr_i[120]), .ZN(n7521) );
  OAI21_X1 U8544 ( .B1(n7523), .B2(n7522), .A(n7521), .ZN(n7524) );
  AOI21_X1 U8545 ( .B1(n7526), .B2(n7525), .A(n7524), .ZN(n7527) );
  OAI21_X1 U8546 ( .B1(n7529), .B2(n7528), .A(n7527), .ZN(n7547) );
  NAND2_X1 U8547 ( .A1(n9438), .A2(pmp_addr_i[121]), .ZN(n7531) );
  NAND2_X1 U8548 ( .A1(n10443), .A2(pmp_addr_i[122]), .ZN(n7530) );
  OAI21_X1 U8549 ( .B1(n7532), .B2(n7531), .A(n7530), .ZN(n7537) );
  NAND2_X1 U8550 ( .A1(n6216), .A2(pmp_addr_i[123]), .ZN(n7534) );
  NAND2_X1 U8551 ( .A1(n8494), .A2(pmp_addr_i[124]), .ZN(n7533) );
  OAI21_X1 U8552 ( .B1(n7535), .B2(n7534), .A(n7533), .ZN(n7536) );
  AOI21_X1 U8553 ( .B1(n7538), .B2(n7537), .A(n7536), .ZN(n7544) );
  NAND2_X1 U8554 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[125]), .ZN(n7540)
         );
  INV_X1 U8555 ( .A(pmp_addr_i[126]), .ZN(n7539) );
  NAND2_X1 U8556 ( .A1(n7540), .A2(n7539), .ZN(n7541) );
  NOR2_X1 U8557 ( .A1(n7541), .A2(pmp_addr_i[127]), .ZN(n7542) );
  OAI21_X1 U8558 ( .B1(n7544), .B2(n7543), .A(n7542), .ZN(n7545) );
  AOI21_X1 U8559 ( .B1(n7547), .B2(n7546), .A(n7545), .ZN(n7548) );
  OAI21_X1 U8560 ( .B1(n7550), .B2(n7549), .A(n7548), .ZN(n7552) );
  OAI211_X1 U8561 ( .C1(n7556), .C2(n9987), .A(n7555), .B(n7554), .ZN(n7567)
         );
  OAI22_X1 U8562 ( .A1(n7557), .A2(n7816), .B1(n11255), .B2(n4182), .ZN(n7558)
         );
  INV_X1 U8563 ( .A(n7558), .ZN(n7562) );
  OAI22_X1 U8564 ( .A1(n10958), .A2(n7606), .B1(n10129), .B2(n157), .ZN(n7559)
         );
  AOI21_X1 U8565 ( .B1(n7560), .B2(n12058), .A(n7559), .ZN(n7561) );
  OAI211_X1 U8566 ( .C1(n7563), .C2(n10953), .A(n7562), .B(n7561), .ZN(n7566)
         );
  OAI22_X1 U8567 ( .A1(n4242), .A2(data_addr_o_12_), .B1(data_addr_o_13_), 
        .B2(n7564), .ZN(n7565) );
  NOR3_X1 U8568 ( .A1(n7567), .A2(n7566), .A3(n7565), .ZN(n7576) );
  OAI22_X1 U8569 ( .A1(data_addr_o_9_), .A2(n4203), .B1(n10281), .B2(n4201), 
        .ZN(n7569) );
  OAI22_X1 U8570 ( .A1(n4205), .A2(n11343), .B1(data_addr_o_11_), .B2(n7360), 
        .ZN(n7568) );
  NOR3_X1 U8571 ( .A1(n7570), .A2(n7569), .A3(n7568), .ZN(n7575) );
  XNOR2_X1 U8572 ( .A(n10967), .B(n7571), .ZN(n7574) );
  XNOR2_X1 U8573 ( .A(n10627), .B(n7572), .ZN(n7573) );
  XNOR2_X1 U8575 ( .A(n10635), .B(n7577), .ZN(n7580) );
  XNOR2_X1 U8576 ( .A(data_addr_o_30_), .B(n7578), .ZN(n7579) );
  XNOR2_X1 U8579 ( .A(n9935), .B(n7583), .ZN(n7590) );
  XNOR2_X1 U8580 ( .A(n10612), .B(n7584), .ZN(n7589) );
  XNOR2_X1 U8581 ( .A(n10638), .B(n7585), .ZN(n7588) );
  XNOR2_X1 U8582 ( .A(data_addr_o_23_), .B(n7586), .ZN(n7587) );
  NAND4_X1 U8583 ( .A1(n7590), .A2(n7589), .A3(n7588), .A4(n7587), .ZN(n7600)
         );
  XNOR2_X1 U8584 ( .A(n10629), .B(n7591), .ZN(n7598) );
  XNOR2_X1 U8585 ( .A(n10614), .B(n7592), .ZN(n7597) );
  XNOR2_X1 U8586 ( .A(n10606), .B(n7593), .ZN(n7596) );
  XNOR2_X1 U8587 ( .A(n10616), .B(n7594), .ZN(n7595) );
  NAND4_X1 U8588 ( .A1(n7598), .A2(n7597), .A3(n7596), .A4(n7595), .ZN(n7599)
         );
  NOR2_X1 U8589 ( .A1(n7600), .A2(n7599), .ZN(n7601) );
  AND2_X1 U8590 ( .A1(n7602), .A2(n7601), .ZN(n11697) );
  XNOR2_X1 U8591 ( .A(n9955), .B(n7603), .ZN(n11742) );
  NAND2_X1 U8592 ( .A1(n11712), .A2(n11709), .ZN(n7610) );
  INV_X1 U8593 ( .A(n7604), .ZN(n7605) );
  AOI21_X1 U8594 ( .B1(n11259), .B2(n157), .A(n7605), .ZN(n7607) );
  NAND2_X1 U8595 ( .A1(data_addr_o_3_), .A2(n7606), .ZN(n11734) );
  AND3_X1 U8596 ( .A1(n11726), .A2(n7607), .A3(n11734), .ZN(n7608) );
  NAND4_X1 U8597 ( .A1(n11748), .A2(n11725), .A3(n11732), .A4(n7608), .ZN(
        n7609) );
  NOR2_X1 U8598 ( .A1(n7610), .A2(n7609), .ZN(n7611) );
  NAND4_X1 U8599 ( .A1(n7611), .A2(n11719), .A3(n11700), .A4(n11699), .ZN(
        n7613) );
  AND2_X1 U8600 ( .A1(data_addr_o_17_), .A2(n4251), .ZN(n11698) );
  NAND4_X1 U8601 ( .A1(n11745), .A2(n11724), .A3(n11747), .A4(n11723), .ZN(
        n7612) );
  NOR3_X1 U8602 ( .A1(n7613), .A2(n11698), .A3(n7612), .ZN(n7616) );
  XNOR2_X1 U8603 ( .A(n12123), .B(n7614), .ZN(n7615) );
  NAND4_X1 U8604 ( .A1(n11697), .A2(n11742), .A3(n7616), .A4(n7615), .ZN(n7617) );
  NAND2_X1 U8605 ( .A1(n7618), .A2(n7617), .ZN(n7621) );
  MUX2_X1 U8606 ( .A(pmp_cfg_i[24]), .B(pmp_cfg_i[25]), .S(n11019), .Z(n7620)
         );
  AND2_X1 U8607 ( .A1(n7619), .A2(n7620), .ZN(n11739) );
  NAND2_X1 U8608 ( .A1(n7621), .A2(n11739), .ZN(n8085) );
  XNOR2_X1 U8609 ( .A(n11285), .B(n7863), .ZN(n7625) );
  XNOR2_X1 U8610 ( .A(n10612), .B(n7859), .ZN(n7624) );
  XNOR2_X1 U8611 ( .A(n10638), .B(n7860), .ZN(n7623) );
  XNOR2_X1 U8612 ( .A(n10898), .B(n7852), .ZN(n7622) );
  NAND4_X1 U8613 ( .A1(n7625), .A2(n7624), .A3(n7623), .A4(n7622), .ZN(n7631)
         );
  XNOR2_X1 U8614 ( .A(n10629), .B(n7853), .ZN(n7629) );
  XNOR2_X1 U8615 ( .A(n10614), .B(n7855), .ZN(n7628) );
  XNOR2_X1 U8616 ( .A(n10606), .B(n7856), .ZN(n7627) );
  XNOR2_X1 U8617 ( .A(n10616), .B(n7867), .ZN(n7626) );
  NAND4_X1 U8618 ( .A1(n7629), .A2(n7628), .A3(n7627), .A4(n7626), .ZN(n7630)
         );
  NOR2_X1 U8619 ( .A1(n7631), .A2(n7630), .ZN(n7645) );
  OAI22_X1 U8620 ( .A1(n7648), .A2(n7816), .B1(n10655), .B2(n7656), .ZN(n7634)
         );
  OAI22_X1 U8621 ( .A1(data_addr_o_9_), .A2(n7667), .B1(n10836), .B2(n7632), 
        .ZN(n7633) );
  AOI211_X1 U8622 ( .C1(n8444), .C2(n7787), .A(n7634), .B(n7633), .ZN(n7641)
         );
  OAI22_X1 U8623 ( .A1(n7659), .A2(n11343), .B1(data_addr_o_11_), .B2(n7660), 
        .ZN(n7635) );
  NOR2_X1 U8624 ( .A1(data_addr_o_12_), .A2(n7646), .ZN(n7833) );
  OR2_X1 U8625 ( .A1(n7635), .A2(n7833), .ZN(n7637) );
  NOR2_X1 U8626 ( .A1(n6649), .A2(n7647), .ZN(n7794) );
  OAI22_X1 U8627 ( .A1(n7652), .A2(n9066), .B1(n11227), .B2(n7651), .ZN(n7636)
         );
  NOR3_X1 U8628 ( .A1(n7637), .A2(n7794), .A3(n7636), .ZN(n7640) );
  XNOR2_X1 U8629 ( .A(n11298), .B(n7786), .ZN(n7639) );
  XNOR2_X1 U8630 ( .A(n10627), .B(n7862), .ZN(n7638) );
  AND4_X1 U8631 ( .A1(n7641), .A2(n7640), .A3(n7639), .A4(n7638), .ZN(n7644)
         );
  XNOR2_X1 U8632 ( .A(n10635), .B(n7868), .ZN(n7643) );
  XNOR2_X1 U8633 ( .A(n10919), .B(n7871), .ZN(n7642) );
  NAND4_X1 U8634 ( .A1(n7645), .A2(n7644), .A3(n7643), .A4(n7642), .ZN(n11083)
         );
  NAND2_X1 U8635 ( .A1(data_addr_o_12_), .A2(n7646), .ZN(n11126) );
  NAND2_X1 U8636 ( .A1(n6649), .A2(n7647), .ZN(n11117) );
  AND2_X1 U8637 ( .A1(n11126), .A2(n11117), .ZN(n7654) );
  NAND2_X1 U8638 ( .A1(n7816), .A2(n7648), .ZN(n11107) );
  XNOR2_X1 U8639 ( .A(n10958), .B(n11097), .ZN(n7650) );
  XNOR2_X1 U8640 ( .A(n11288), .B(n11101), .ZN(n7649) );
  AND3_X1 U8641 ( .A1(n11107), .A2(n7650), .A3(n7649), .ZN(n7653) );
  NAND2_X1 U8642 ( .A1(n10657), .A2(n7651), .ZN(n11095) );
  NAND2_X1 U8643 ( .A1(data_addr_o_14_), .A2(n7652), .ZN(n11113) );
  NAND4_X1 U8644 ( .A1(n7654), .A2(n7653), .A3(n11095), .A4(n11113), .ZN(n7665) );
  XNOR2_X1 U8645 ( .A(n9987), .B(n7655), .ZN(n7664) );
  NAND2_X1 U8646 ( .A1(n10655), .A2(n7656), .ZN(n11084) );
  XNOR2_X1 U8647 ( .A(n11259), .B(n7800), .ZN(n7657) );
  AND3_X1 U8648 ( .A1(n11084), .A2(n7658), .A3(n7657), .ZN(n7662) );
  NAND2_X1 U8649 ( .A1(n10838), .A2(n7659), .ZN(n11112) );
  NAND2_X1 U8650 ( .A1(data_addr_o_11_), .A2(n7660), .ZN(n11091) );
  XNOR2_X1 U8651 ( .A(n10824), .B(n7797), .ZN(n7661) );
  NAND4_X1 U8652 ( .A1(n7662), .A2(n11112), .A3(n11091), .A4(n7661), .ZN(n7663) );
  NOR3_X1 U8653 ( .A1(n7665), .A2(n7664), .A3(n7663), .ZN(n7670) );
  XNOR2_X1 U8654 ( .A(n11303), .B(n7870), .ZN(n11136) );
  XNOR2_X1 U8655 ( .A(n12123), .B(n7874), .ZN(n7669) );
  AND2_X1 U8656 ( .A1(data_addr_o_17_), .A2(n7666), .ZN(n11135) );
  NAND2_X1 U8657 ( .A1(data_addr_o_9_), .A2(n7667), .ZN(n11124) );
  OAI21_X1 U8658 ( .B1(n7814), .B2(n7815), .A(n11124), .ZN(n11093) );
  NOR2_X1 U8659 ( .A1(n11135), .A2(n11093), .ZN(n7668) );
  NAND4_X1 U8660 ( .A1(n7670), .A2(n11136), .A3(n7669), .A4(n7668), .ZN(n7926)
         );
  NOR2_X1 U8661 ( .A1(n7482), .A2(n7715), .ZN(n7718) );
  NOR2_X1 U8662 ( .A1(n10721), .A2(pmp_addr_i[461]), .ZN(n7671) );
  NOR2_X1 U8663 ( .A1(n7718), .A2(n7671), .ZN(n7673) );
  NOR2_X1 U8664 ( .A1(n10297), .A2(pmp_addr_i[464]), .ZN(n7721) );
  NOR2_X1 U8665 ( .A1(n7995), .A2(pmp_addr_i[463]), .ZN(n7672) );
  NOR2_X1 U8666 ( .A1(n7721), .A2(n7672), .ZN(n7723) );
  NAND2_X1 U8667 ( .A1(n7673), .A2(n7723), .ZN(n7727) );
  NOR2_X1 U8668 ( .A1(n9508), .A2(pmp_addr_i[457]), .ZN(n7674) );
  NOR2_X1 U8669 ( .A1(n7472), .A2(pmp_addr_i[458]), .ZN(n7708) );
  NOR2_X1 U8670 ( .A1(n7674), .A2(n7708), .ZN(n7676) );
  NOR2_X1 U8671 ( .A1(n10342), .A2(pmp_addr_i[459]), .ZN(n7675) );
  NOR2_X1 U8672 ( .A1(n11334), .A2(pmp_addr_i[460]), .ZN(n7711) );
  NOR2_X1 U8673 ( .A1(n7675), .A2(n7711), .ZN(n7714) );
  NAND2_X1 U8674 ( .A1(n7676), .A2(n7714), .ZN(n7677) );
  NOR2_X1 U8675 ( .A1(n7727), .A2(n7677), .ZN(n7730) );
  NOR2_X1 U8676 ( .A1(n10346), .A2(pmp_addr_i[451]), .ZN(n7678) );
  NOR2_X1 U8677 ( .A1(n8410), .A2(pmp_addr_i[452]), .ZN(n7687) );
  NOR2_X1 U8678 ( .A1(n7678), .A2(n7687), .ZN(n7690) );
  OR2_X1 U8679 ( .A1(pmp_addr_i[449]), .A2(n10473), .ZN(n7681) );
  AND2_X1 U8680 ( .A1(n10651), .A2(pmp_addr_i[448]), .ZN(n7680) );
  AND2_X1 U8681 ( .A1(pmp_addr_i[449]), .A2(n10010), .ZN(n7679) );
  AOI21_X1 U8682 ( .B1(n7681), .B2(n7680), .A(n7679), .ZN(n7684) );
  NOR2_X1 U8683 ( .A1(pmp_addr_i[450]), .A2(n8406), .ZN(n7683) );
  NAND2_X1 U8684 ( .A1(pmp_addr_i[450]), .A2(n10351), .ZN(n7682) );
  OAI21_X1 U8685 ( .B1(n7684), .B2(n7683), .A(n7682), .ZN(n7689) );
  NAND2_X1 U8686 ( .A1(n10346), .A2(pmp_addr_i[451]), .ZN(n7686) );
  NAND2_X1 U8687 ( .A1(n10362), .A2(pmp_addr_i[452]), .ZN(n7685) );
  OAI21_X1 U8688 ( .B1(n7687), .B2(n7686), .A(n7685), .ZN(n7688) );
  AOI21_X1 U8689 ( .B1(n7690), .B2(n7689), .A(n7688), .ZN(n7705) );
  NOR2_X1 U8690 ( .A1(n29), .A2(pmp_addr_i[454]), .ZN(n7696) );
  NOR2_X1 U8691 ( .A1(n6400), .A2(pmp_addr_i[453]), .ZN(n7691) );
  NOR2_X1 U8692 ( .A1(n7696), .A2(n7691), .ZN(n7693) );
  NOR2_X1 U8693 ( .A1(n10501), .A2(pmp_addr_i[455]), .ZN(n7692) );
  NOR2_X1 U8694 ( .A1(n7820), .A2(pmp_addr_i[456]), .ZN(n7699) );
  NOR2_X1 U8695 ( .A1(n7692), .A2(n7699), .ZN(n7702) );
  NAND2_X1 U8696 ( .A1(n7693), .A2(n7702), .ZN(n7704) );
  NAND2_X1 U8697 ( .A1(n6400), .A2(pmp_addr_i[453]), .ZN(n7695) );
  NAND2_X1 U8698 ( .A1(n8735), .A2(pmp_addr_i[454]), .ZN(n7694) );
  OAI21_X1 U8699 ( .B1(n7696), .B2(n7695), .A(n7694), .ZN(n7701) );
  NAND2_X1 U8700 ( .A1(n10501), .A2(pmp_addr_i[455]), .ZN(n7698) );
  NAND2_X1 U8701 ( .A1(n7964), .A2(pmp_addr_i[456]), .ZN(n7697) );
  OAI21_X1 U8702 ( .B1(n7699), .B2(n7698), .A(n7697), .ZN(n7700) );
  AOI21_X1 U8703 ( .B1(n7702), .B2(n7701), .A(n7700), .ZN(n7703) );
  OAI21_X1 U8704 ( .B1(n7705), .B2(n7704), .A(n7703), .ZN(n7729) );
  NAND2_X1 U8705 ( .A1(n9508), .A2(pmp_addr_i[457]), .ZN(n7707) );
  NAND2_X1 U8706 ( .A1(n7472), .A2(pmp_addr_i[458]), .ZN(n7706) );
  OAI21_X1 U8707 ( .B1(n7708), .B2(n7707), .A(n7706), .ZN(n7713) );
  NAND2_X1 U8708 ( .A1(n10342), .A2(pmp_addr_i[459]), .ZN(n7710) );
  NAND2_X1 U8709 ( .A1(n11334), .A2(pmp_addr_i[460]), .ZN(n7709) );
  OAI21_X1 U8710 ( .B1(n7711), .B2(n7710), .A(n7709), .ZN(n7712) );
  AOI21_X1 U8711 ( .B1(n7714), .B2(n7713), .A(n7712), .ZN(n7726) );
  NAND2_X1 U8712 ( .A1(n10721), .A2(pmp_addr_i[461]), .ZN(n7717) );
  NAND2_X1 U8713 ( .A1(n7990), .A2(n7715), .ZN(n7716) );
  OAI21_X1 U8714 ( .B1(n7718), .B2(n7717), .A(n7716), .ZN(n7724) );
  NAND2_X1 U8715 ( .A1(n8444), .A2(pmp_addr_i[463]), .ZN(n7720) );
  NAND2_X1 U8716 ( .A1(n12184), .A2(pmp_addr_i[464]), .ZN(n7719) );
  OAI21_X1 U8717 ( .B1(n7721), .B2(n7720), .A(n7719), .ZN(n7722) );
  AOI21_X1 U8718 ( .B1(n7724), .B2(n7723), .A(n7722), .ZN(n7725) );
  OAI21_X1 U8719 ( .B1(n7727), .B2(n7726), .A(n7725), .ZN(n7728) );
  AOI21_X1 U8720 ( .B1(n7730), .B2(n7729), .A(n7728), .ZN(n7783) );
  NOR2_X1 U8721 ( .A1(n10424), .A2(pmp_addr_i[469]), .ZN(n7731) );
  NOR2_X1 U8722 ( .A1(n9163), .A2(pmp_addr_i[470]), .ZN(n7754) );
  NOR2_X1 U8723 ( .A1(n7731), .A2(n7754), .ZN(n7733) );
  NOR2_X1 U8724 ( .A1(n10429), .A2(pmp_addr_i[471]), .ZN(n7732) );
  NOR2_X1 U8725 ( .A1(n6202), .A2(pmp_addr_i[472]), .ZN(n7757) );
  NOR2_X1 U8726 ( .A1(n7732), .A2(n7757), .ZN(n7760) );
  NAND2_X1 U8727 ( .A1(n7733), .A2(n7760), .ZN(n7762) );
  NOR2_X1 U8728 ( .A1(n9418), .A2(pmp_addr_i[467]), .ZN(n7734) );
  NOR2_X1 U8729 ( .A1(n9156), .A2(pmp_addr_i[468]), .ZN(n7748) );
  NOR2_X1 U8730 ( .A1(n7734), .A2(n7748), .ZN(n7751) );
  NOR2_X1 U8731 ( .A1(n9414), .A2(pmp_addr_i[465]), .ZN(n7735) );
  NOR2_X1 U8732 ( .A1(n10754), .A2(pmp_addr_i[466]), .ZN(n7745) );
  NOR2_X1 U8733 ( .A1(n7735), .A2(n7745), .ZN(n7736) );
  NAND2_X1 U8734 ( .A1(n7751), .A2(n7736), .ZN(n7737) );
  NOR2_X1 U8735 ( .A1(n7762), .A2(n7737), .ZN(n7742) );
  NOR2_X1 U8736 ( .A1(n6212), .A2(pmp_addr_i[473]), .ZN(n7738) );
  NOR2_X1 U8737 ( .A1(n10443), .A2(pmp_addr_i[474]), .ZN(n7766) );
  NOR2_X1 U8738 ( .A1(n7738), .A2(n7766), .ZN(n7740) );
  NOR2_X1 U8739 ( .A1(n6216), .A2(pmp_addr_i[475]), .ZN(n7739) );
  NOR2_X1 U8740 ( .A1(n8494), .A2(pmp_addr_i[476]), .ZN(n7769) );
  NOR2_X1 U8741 ( .A1(n7739), .A2(n7769), .ZN(n7772) );
  NAND2_X1 U8742 ( .A1(n7740), .A2(n7772), .ZN(n7741) );
  NOR2_X1 U8743 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[477]), .ZN(n7776)
         );
  NOR2_X1 U8744 ( .A1(n7741), .A2(n7776), .ZN(n7779) );
  NAND2_X1 U8745 ( .A1(n7742), .A2(n7779), .ZN(n7782) );
  NAND2_X1 U8746 ( .A1(n10414), .A2(pmp_addr_i[465]), .ZN(n7744) );
  NAND2_X1 U8747 ( .A1(n10754), .A2(pmp_addr_i[466]), .ZN(n7743) );
  OAI21_X1 U8748 ( .B1(n7745), .B2(n7744), .A(n7743), .ZN(n7750) );
  NAND2_X1 U8749 ( .A1(n6192), .A2(pmp_addr_i[467]), .ZN(n7747) );
  NAND2_X1 U8750 ( .A1(n9156), .A2(pmp_addr_i[468]), .ZN(n7746) );
  OAI21_X1 U8751 ( .B1(n7748), .B2(n7747), .A(n7746), .ZN(n7749) );
  AOI21_X1 U8752 ( .B1(n7751), .B2(n7750), .A(n7749), .ZN(n7763) );
  NAND2_X1 U8753 ( .A1(n10424), .A2(pmp_addr_i[469]), .ZN(n7753) );
  NAND2_X1 U8754 ( .A1(n10428), .A2(pmp_addr_i[470]), .ZN(n7752) );
  OAI21_X1 U8755 ( .B1(n7754), .B2(n7753), .A(n7752), .ZN(n7759) );
  NAND2_X1 U8756 ( .A1(n10429), .A2(pmp_addr_i[471]), .ZN(n7756) );
  NAND2_X1 U8757 ( .A1(n6202), .A2(pmp_addr_i[472]), .ZN(n7755) );
  OAI21_X1 U8758 ( .B1(n7757), .B2(n7756), .A(n7755), .ZN(n7758) );
  AOI21_X1 U8759 ( .B1(n7760), .B2(n7759), .A(n7758), .ZN(n7761) );
  OAI21_X1 U8760 ( .B1(n7763), .B2(n7762), .A(n7761), .ZN(n7780) );
  NAND2_X1 U8761 ( .A1(n6212), .A2(pmp_addr_i[473]), .ZN(n7765) );
  NAND2_X1 U8762 ( .A1(n8807), .A2(pmp_addr_i[474]), .ZN(n7764) );
  OAI21_X1 U8763 ( .B1(n7766), .B2(n7765), .A(n7764), .ZN(n7771) );
  NAND2_X1 U8764 ( .A1(n10782), .A2(pmp_addr_i[475]), .ZN(n7768) );
  NAND2_X1 U8765 ( .A1(n8494), .A2(pmp_addr_i[476]), .ZN(n7767) );
  OAI21_X1 U8766 ( .B1(n7769), .B2(n7768), .A(n7767), .ZN(n7770) );
  AOI21_X1 U8767 ( .B1(n7772), .B2(n7771), .A(n7770), .ZN(n7777) );
  NAND2_X1 U8768 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[477]), .ZN(n7773)
         );
  NAND2_X1 U8769 ( .A1(n7773), .A2(n4007), .ZN(n7774) );
  NOR2_X1 U8770 ( .A1(n7774), .A2(pmp_addr_i[479]), .ZN(n7775) );
  OAI21_X1 U8771 ( .B1(n7777), .B2(n7776), .A(n7775), .ZN(n7778) );
  AOI21_X1 U8772 ( .B1(n7780), .B2(n7779), .A(n7778), .ZN(n7781) );
  OAI21_X1 U8773 ( .B1(n7783), .B2(n7782), .A(n7781), .ZN(n7924) );
  NOR2_X1 U8774 ( .A1(data_addr_o_16_), .A2(n7655), .ZN(n7839) );
  NOR2_X1 U8775 ( .A1(n11309), .A2(n7651), .ZN(n7785) );
  NOR2_X1 U8776 ( .A1(n7839), .A2(n7785), .ZN(n7789) );
  NOR2_X1 U8777 ( .A1(n10967), .A2(n2438), .ZN(n7842) );
  NOR2_X1 U8778 ( .A1(n6813), .A2(n7666), .ZN(n7788) );
  NOR2_X1 U8779 ( .A1(n7842), .A2(n7788), .ZN(n7844) );
  NAND2_X1 U8780 ( .A1(n7789), .A2(n7844), .ZN(n7848) );
  NOR2_X1 U8781 ( .A1(data_addr_o_11_), .A2(n7660), .ZN(n7792) );
  NOR2_X1 U8782 ( .A1(n7792), .A2(n7833), .ZN(n7795) );
  NOR2_X1 U8783 ( .A1(data_addr_o_14_), .A2(n7652), .ZN(n7834) );
  NOR2_X1 U8784 ( .A1(n7794), .A2(n7834), .ZN(n7837) );
  NAND2_X1 U8785 ( .A1(n7795), .A2(n7837), .ZN(n7796) );
  NOR2_X1 U8786 ( .A1(n7848), .A2(n7796), .ZN(n7851) );
  NOR2_X1 U8787 ( .A1(data_addr_o_5_), .A2(n11122), .ZN(n7799) );
  NOR2_X1 U8788 ( .A1(n10358), .A2(n7656), .ZN(n7810) );
  NOR2_X1 U8789 ( .A1(n7799), .A2(n7810), .ZN(n7813) );
  INV_X1 U8790 ( .A(n10651), .ZN(n10129) );
  INV_X1 U8791 ( .A(n7800), .ZN(n7801) );
  OR2_X1 U8792 ( .A1(n10129), .A2(n7801), .ZN(n7805) );
  INV_X1 U8793 ( .A(n11097), .ZN(n7802) );
  OR2_X1 U8794 ( .A1(n10130), .A2(n7802), .ZN(n7804) );
  AND2_X1 U8795 ( .A1(n10130), .A2(n7802), .ZN(n7803) );
  AOI21_X1 U8796 ( .B1(n7805), .B2(n7804), .A(n7803), .ZN(n7808) );
  INV_X1 U8797 ( .A(n12058), .ZN(n10135) );
  NOR2_X1 U8798 ( .A1(n10135), .A2(n11103), .ZN(n7807) );
  NAND2_X1 U8799 ( .A1(n10135), .A2(n11103), .ZN(n7806) );
  OAI21_X1 U8800 ( .B1(n7808), .B2(n7807), .A(n7806), .ZN(n7812) );
  NAND2_X1 U8801 ( .A1(n10486), .A2(n11122), .ZN(n7809) );
  OAI21_X1 U8802 ( .B1(n7810), .B2(n7809), .A(n11084), .ZN(n7811) );
  AOI21_X1 U8803 ( .B1(n7813), .B2(n7812), .A(n7811), .ZN(n7832) );
  INV_X1 U8804 ( .A(n7814), .ZN(n9805) );
  NOR2_X1 U8805 ( .A1(n9805), .A2(n7632), .ZN(n7825) );
  NOR2_X1 U8806 ( .A1(n7816), .A2(n7648), .ZN(n7818) );
  NOR2_X1 U8807 ( .A1(n7825), .A2(n7818), .ZN(n7823) );
  NOR2_X1 U8808 ( .A1(data_addr_o_9_), .A2(n7667), .ZN(n7822) );
  NOR2_X1 U8809 ( .A1(data_addr_o_10_), .A2(n7659), .ZN(n7826) );
  NOR2_X1 U8810 ( .A1(n7822), .A2(n7826), .ZN(n7829) );
  NAND2_X1 U8811 ( .A1(n7823), .A2(n7829), .ZN(n7831) );
  NAND2_X1 U8812 ( .A1(n9805), .A2(n7632), .ZN(n7824) );
  OAI21_X1 U8813 ( .B1(n7825), .B2(n11107), .A(n7824), .ZN(n7828) );
  OAI21_X1 U8814 ( .B1(n7826), .B2(n11124), .A(n11112), .ZN(n7827) );
  AOI21_X1 U8815 ( .B1(n7829), .B2(n7828), .A(n7827), .ZN(n7830) );
  OAI21_X1 U8816 ( .B1(n7832), .B2(n7831), .A(n7830), .ZN(n7850) );
  OAI21_X1 U8817 ( .B1(n7833), .B2(n11091), .A(n11126), .ZN(n7836) );
  OAI21_X1 U8818 ( .B1(n7834), .B2(n11117), .A(n11113), .ZN(n7835) );
  AOI21_X1 U8819 ( .B1(n7837), .B2(n7836), .A(n7835), .ZN(n7847) );
  NAND2_X1 U8820 ( .A1(data_addr_o_16_), .A2(n7655), .ZN(n7838) );
  OAI21_X1 U8821 ( .B1(n7839), .B2(n11095), .A(n7838), .ZN(n7845) );
  NAND2_X1 U8822 ( .A1(n6813), .A2(n7666), .ZN(n7841) );
  NAND2_X1 U8823 ( .A1(n10967), .A2(n2438), .ZN(n7840) );
  OAI21_X1 U8824 ( .B1(n7842), .B2(n7841), .A(n7840), .ZN(n7843) );
  AOI21_X1 U8825 ( .B1(n7845), .B2(n7844), .A(n7843), .ZN(n7846) );
  OAI21_X1 U8826 ( .B1(n7848), .B2(n7847), .A(n7846), .ZN(n7849) );
  AOI21_X1 U8827 ( .B1(n7851), .B2(n7850), .A(n7849), .ZN(n7921) );
  NOR2_X1 U8828 ( .A1(data_addr_o_23_), .A2(n2529), .ZN(n7854) );
  NOR2_X1 U8829 ( .A1(n10738), .A2(n2490), .ZN(n7891) );
  NOR2_X1 U8830 ( .A1(n7854), .A2(n7891), .ZN(n7858) );
  NOR2_X1 U8831 ( .A1(n11320), .A2(n2532), .ZN(n7857) );
  NOR2_X1 U8832 ( .A1(data_addr_o_26_), .A2(n2482), .ZN(n7894) );
  NOR2_X1 U8833 ( .A1(n7857), .A2(n7894), .ZN(n7897) );
  NAND2_X1 U8834 ( .A1(n7858), .A2(n7897), .ZN(n7899) );
  NOR2_X1 U8835 ( .A1(n11312), .A2(n2520), .ZN(n7861) );
  NOR2_X1 U8836 ( .A1(n11313), .A2(n3289), .ZN(n7885) );
  NOR2_X1 U8837 ( .A1(n7861), .A2(n7885), .ZN(n7888) );
  NOR2_X1 U8838 ( .A1(n11283), .A2(n2517), .ZN(n7864) );
  NOR2_X1 U8839 ( .A1(n11285), .A2(n3291), .ZN(n7882) );
  NOR2_X1 U8840 ( .A1(n7864), .A2(n7882), .ZN(n7865) );
  NAND2_X1 U8841 ( .A1(n7888), .A2(n7865), .ZN(n7866) );
  NOR2_X1 U8842 ( .A1(n7899), .A2(n7866), .ZN(n7879) );
  NOR2_X1 U8843 ( .A1(n11322), .A2(n2545), .ZN(n7869) );
  INV_X1 U8844 ( .A(n7868), .ZN(n7901) );
  NOR2_X1 U8845 ( .A1(n10635), .A2(n7901), .ZN(n7904) );
  NOR2_X1 U8846 ( .A1(n7869), .A2(n7904), .ZN(n7873) );
  NOR2_X1 U8847 ( .A1(n11303), .A2(n2548), .ZN(n7872) );
  NOR2_X1 U8848 ( .A1(data_addr_o_30_), .A2(n2550), .ZN(n7907) );
  NOR2_X1 U8849 ( .A1(n7872), .A2(n7907), .ZN(n7910) );
  NOR2_X1 U8851 ( .A1(n10662), .A2(n2549), .ZN(n7875) );
  NOR2_X1 U8852 ( .A1(n7875), .A2(pmp_addr_i[446]), .ZN(n7877) );
  INV_X1 U8853 ( .A(pmp_addr_i[447]), .ZN(n7876) );
  NAND2_X1 U8854 ( .A1(n7877), .A2(n7876), .ZN(n7914) );
  NAND2_X1 U8856 ( .A1(n7879), .A2(n7917), .ZN(n7920) );
  NAND2_X1 U8857 ( .A1(n11283), .A2(n2517), .ZN(n7881) );
  NAND2_X1 U8858 ( .A1(n11285), .A2(n3291), .ZN(n7880) );
  OAI21_X1 U8859 ( .B1(n7882), .B2(n7881), .A(n7880), .ZN(n7887) );
  NAND2_X1 U8860 ( .A1(n11312), .A2(n2520), .ZN(n7884) );
  NAND2_X1 U8861 ( .A1(n11313), .A2(n3289), .ZN(n7883) );
  OAI21_X1 U8862 ( .B1(n7885), .B2(n7884), .A(n7883), .ZN(n7886) );
  AOI21_X1 U8863 ( .B1(n7888), .B2(n7887), .A(n7886), .ZN(n7900) );
  NAND2_X1 U8864 ( .A1(data_addr_o_23_), .A2(n2529), .ZN(n7890) );
  NAND2_X1 U8865 ( .A1(n10899), .A2(n2490), .ZN(n7889) );
  OAI21_X1 U8866 ( .B1(n7891), .B2(n7890), .A(n7889), .ZN(n7896) );
  NAND2_X1 U8867 ( .A1(n11320), .A2(n2532), .ZN(n7893) );
  NAND2_X1 U8868 ( .A1(data_addr_o_26_), .A2(n2482), .ZN(n7892) );
  OAI21_X1 U8869 ( .B1(n7894), .B2(n7893), .A(n7892), .ZN(n7895) );
  AOI21_X1 U8870 ( .B1(n7897), .B2(n7896), .A(n7895), .ZN(n7898) );
  OAI21_X1 U8871 ( .B1(n7900), .B2(n7899), .A(n7898), .ZN(n7918) );
  NAND2_X1 U8872 ( .A1(n11322), .A2(n2545), .ZN(n7903) );
  NAND2_X1 U8873 ( .A1(n10747), .A2(n7901), .ZN(n7902) );
  OAI21_X1 U8874 ( .B1(n7904), .B2(n7903), .A(n7902), .ZN(n7909) );
  NAND2_X1 U8875 ( .A1(n11303), .A2(n2548), .ZN(n7906) );
  NAND2_X1 U8876 ( .A1(data_addr_o_30_), .A2(n2550), .ZN(n7905) );
  OAI21_X1 U8877 ( .B1(n7907), .B2(n7906), .A(n7905), .ZN(n7908) );
  AOI21_X1 U8878 ( .B1(n7910), .B2(n7909), .A(n7908), .ZN(n7915) );
  NAND2_X1 U8879 ( .A1(n10662), .A2(n2549), .ZN(n7911) );
  NOR2_X1 U8880 ( .A1(n7911), .A2(pmp_addr_i[446]), .ZN(n7912) );
  NAND2_X1 U8881 ( .A1(n7912), .A2(n7876), .ZN(n7913) );
  OAI21_X1 U8882 ( .B1(n7915), .B2(n7914), .A(n7913), .ZN(n7916) );
  AOI21_X1 U8883 ( .B1(n7918), .B2(n7917), .A(n7916), .ZN(n7919) );
  OAI21_X1 U8884 ( .B1(n7921), .B2(n7920), .A(n7919), .ZN(n7922) );
  NAND3_X1 U8885 ( .A1(n7924), .A2(n7923), .A3(n7922), .ZN(n7925) );
  OAI21_X1 U8886 ( .B1(n11083), .B2(n7926), .A(n7925), .ZN(n7929) );
  MUX2_X1 U8887 ( .A(pmp_cfg_i[112]), .B(pmp_cfg_i[113]), .S(n11019), .Z(n7928) );
  AND2_X1 U8888 ( .A1(n7927), .A2(n7928), .ZN(n11085) );
  NAND2_X1 U8889 ( .A1(n7929), .A2(n11085), .ZN(n8084) );
  INV_X1 U8890 ( .A(n11014), .ZN(n7990) );
  NOR2_X1 U8891 ( .A1(n7990), .A2(n7989), .ZN(n7993) );
  NOR2_X1 U8892 ( .A1(n10721), .A2(n7988), .ZN(n7930) );
  NOR2_X1 U8893 ( .A1(n7993), .A2(n7930), .ZN(n7931) );
  NOR2_X1 U8894 ( .A1(n12184), .A2(n7996), .ZN(n7998) );
  INV_X1 U8895 ( .A(data_addr_i[17]), .ZN(n7995) );
  NOR2_X1 U8896 ( .A1(n7995), .A2(n7994), .ZN(n11225) );
  NOR2_X1 U8897 ( .A1(n7998), .A2(n11225), .ZN(n8000) );
  NAND2_X1 U8898 ( .A1(n7931), .A2(n8000), .ZN(n8004) );
  NOR2_X1 U8899 ( .A1(n10711), .A2(n7974), .ZN(n7932) );
  INV_X1 U8900 ( .A(data_addr_o_12_), .ZN(n7976) );
  NOR2_X1 U8901 ( .A1(n7976), .A2(n7975), .ZN(n7979) );
  NOR2_X1 U8902 ( .A1(n7932), .A2(n7979), .ZN(n7934) );
  NOR2_X1 U8903 ( .A1(n10342), .A2(n7980), .ZN(n7933) );
  NOR2_X1 U8904 ( .A1(n6154), .A2(n7981), .ZN(n7984) );
  NOR2_X1 U8905 ( .A1(n7933), .A2(n7984), .ZN(n7987) );
  NAND2_X1 U8906 ( .A1(n7934), .A2(n7987), .ZN(n7935) );
  NOR2_X1 U8907 ( .A1(n8004), .A2(n7935), .ZN(n8007) );
  NOR2_X1 U8908 ( .A1(n6127), .A2(n7946), .ZN(n7936) );
  NOR2_X1 U8909 ( .A1(n8410), .A2(n7947), .ZN(n7950) );
  NOR2_X1 U8910 ( .A1(n7936), .A2(n7950), .ZN(n7953) );
  OR2_X1 U8911 ( .A1(n10010), .A2(n7938), .ZN(n7941) );
  AND2_X1 U8912 ( .A1(n10651), .A2(n7937), .ZN(n7940) );
  AND2_X1 U8913 ( .A1(n10010), .A2(n7938), .ZN(n7939) );
  AOI21_X1 U8914 ( .B1(n7941), .B2(n7940), .A(n7939), .ZN(n7945) );
  NOR2_X1 U8915 ( .A1(n6123), .A2(n7942), .ZN(n7944) );
  NAND2_X1 U8916 ( .A1(n6123), .A2(n7942), .ZN(n7943) );
  OAI21_X1 U8917 ( .B1(n7945), .B2(n7944), .A(n7943), .ZN(n7952) );
  NAND2_X1 U8918 ( .A1(n6127), .A2(n7946), .ZN(n7949) );
  NAND2_X1 U8919 ( .A1(n9363), .A2(n7947), .ZN(n7948) );
  OAI21_X1 U8920 ( .B1(n7950), .B2(n7949), .A(n7948), .ZN(n7951) );
  AOI21_X1 U8921 ( .B1(n7953), .B2(n7952), .A(n7951), .ZN(n7973) );
  NOR2_X1 U8922 ( .A1(n29), .A2(n7958), .ZN(n7961) );
  NOR2_X1 U8923 ( .A1(n10697), .A2(n7957), .ZN(n7954) );
  NOR2_X1 U8924 ( .A1(n7961), .A2(n7954), .ZN(n7956) );
  NOR2_X1 U8925 ( .A1(n6140), .A2(n7962), .ZN(n7955) );
  INV_X1 U8926 ( .A(n8238), .ZN(n7964) );
  NOR2_X1 U8927 ( .A1(n7964), .A2(n7963), .ZN(n7967) );
  NOR2_X1 U8928 ( .A1(n7955), .A2(n7967), .ZN(n7970) );
  NAND2_X1 U8929 ( .A1(n7956), .A2(n7970), .ZN(n7972) );
  NAND2_X1 U8930 ( .A1(n10697), .A2(n7957), .ZN(n7960) );
  NAND2_X1 U8931 ( .A1(n29), .A2(n7958), .ZN(n7959) );
  OAI21_X1 U8932 ( .B1(n7961), .B2(n7960), .A(n7959), .ZN(n7969) );
  NAND2_X1 U8933 ( .A1(n10501), .A2(n7962), .ZN(n7966) );
  NAND2_X1 U8934 ( .A1(n7964), .A2(n7963), .ZN(n7965) );
  OAI21_X1 U8935 ( .B1(n7967), .B2(n7966), .A(n7965), .ZN(n7968) );
  AOI21_X1 U8936 ( .B1(n7970), .B2(n7969), .A(n7968), .ZN(n7971) );
  OAI21_X1 U8937 ( .B1(n7973), .B2(n7972), .A(n7971), .ZN(n8006) );
  NAND2_X1 U8938 ( .A1(n7324), .A2(n7974), .ZN(n7978) );
  NAND2_X1 U8939 ( .A1(n7976), .A2(n7975), .ZN(n7977) );
  OAI21_X1 U8940 ( .B1(n7979), .B2(n7978), .A(n7977), .ZN(n7986) );
  NAND2_X1 U8941 ( .A1(n10342), .A2(n7980), .ZN(n7983) );
  NAND2_X1 U8942 ( .A1(n6154), .A2(n7981), .ZN(n7982) );
  OAI21_X1 U8943 ( .B1(n7984), .B2(n7983), .A(n7982), .ZN(n7985) );
  AOI21_X1 U8944 ( .B1(n7987), .B2(n7986), .A(n7985), .ZN(n8003) );
  NAND2_X1 U8945 ( .A1(n10338), .A2(n7988), .ZN(n7992) );
  NAND2_X1 U8946 ( .A1(n7990), .A2(n7989), .ZN(n7991) );
  OAI21_X1 U8947 ( .B1(n7993), .B2(n7992), .A(n7991), .ZN(n8001) );
  NAND2_X1 U8948 ( .A1(n7995), .A2(n7994), .ZN(n11308) );
  NAND2_X1 U8949 ( .A1(n10403), .A2(n7996), .ZN(n7997) );
  OAI21_X1 U8950 ( .B1(n7998), .B2(n11308), .A(n7997), .ZN(n7999) );
  AOI21_X1 U8951 ( .B1(n8001), .B2(n8000), .A(n7999), .ZN(n8002) );
  OAI21_X1 U8952 ( .B1(n8004), .B2(n8003), .A(n8002), .ZN(n8005) );
  AOI21_X1 U8953 ( .B1(n8007), .B2(n8006), .A(n8005), .ZN(n8076) );
  NOR2_X1 U8954 ( .A1(n10424), .A2(n8033), .ZN(n8008) );
  NOR2_X1 U8955 ( .A1(n9163), .A2(n8034), .ZN(n8037) );
  NOR2_X1 U8956 ( .A1(n8008), .A2(n8037), .ZN(n8010) );
  NOR2_X1 U8957 ( .A1(n6462), .A2(n8038), .ZN(n8009) );
  NOR2_X1 U8958 ( .A1(n10439), .A2(n8039), .ZN(n8042) );
  NOR2_X1 U8959 ( .A1(n8009), .A2(n8042), .ZN(n8045) );
  NAND2_X1 U8960 ( .A1(n8010), .A2(n8045), .ZN(n8047) );
  NOR2_X1 U8961 ( .A1(n9418), .A2(n8025), .ZN(n8011) );
  NOR2_X1 U8962 ( .A1(n9425), .A2(n8026), .ZN(n8029) );
  NOR2_X1 U8963 ( .A1(n8011), .A2(n8029), .ZN(n8032) );
  NOR2_X1 U8964 ( .A1(n9414), .A2(n8020), .ZN(n8012) );
  NOR2_X1 U8965 ( .A1(n10295), .A2(n8021), .ZN(n8024) );
  NOR2_X1 U8966 ( .A1(n8012), .A2(n8024), .ZN(n8013) );
  NAND2_X1 U8967 ( .A1(n8032), .A2(n8013), .ZN(n8014) );
  NOR2_X1 U8968 ( .A1(n8047), .A2(n8014), .ZN(n8019) );
  NOR2_X1 U8969 ( .A1(n9438), .A2(n8049), .ZN(n8015) );
  NOR2_X1 U8970 ( .A1(n10778), .A2(n8050), .ZN(n8053) );
  NOR2_X1 U8971 ( .A1(n8015), .A2(n8053), .ZN(n8017) );
  NOR2_X1 U8972 ( .A1(n10782), .A2(n8054), .ZN(n8016) );
  NOR2_X1 U8973 ( .A1(n8494), .A2(n8055), .ZN(n8058) );
  NOR2_X1 U8974 ( .A1(n8016), .A2(n8058), .ZN(n8061) );
  NAND2_X1 U8975 ( .A1(n8017), .A2(n8061), .ZN(n8018) );
  NOR2_X1 U8976 ( .A1(data_addr_o_31__BAR), .A2(n8062), .ZN(n8069) );
  NOR2_X1 U8977 ( .A1(n8018), .A2(n8069), .ZN(n8072) );
  NAND2_X1 U8978 ( .A1(n8019), .A2(n8072), .ZN(n8075) );
  NAND2_X1 U8979 ( .A1(n9414), .A2(n8020), .ZN(n8023) );
  NAND2_X1 U8980 ( .A1(n6188), .A2(n8021), .ZN(n8022) );
  OAI21_X1 U8981 ( .B1(n8024), .B2(n8023), .A(n8022), .ZN(n8031) );
  NAND2_X1 U8982 ( .A1(n6192), .A2(n8025), .ZN(n8028) );
  NAND2_X1 U8983 ( .A1(n9425), .A2(n8026), .ZN(n8027) );
  OAI21_X1 U8984 ( .B1(n8029), .B2(n8028), .A(n8027), .ZN(n8030) );
  AOI21_X1 U8985 ( .B1(n8032), .B2(n8031), .A(n8030), .ZN(n8048) );
  NAND2_X1 U8986 ( .A1(n10424), .A2(n8033), .ZN(n8036) );
  NAND2_X1 U8987 ( .A1(n10428), .A2(n8034), .ZN(n8035) );
  OAI21_X1 U8988 ( .B1(n8037), .B2(n8036), .A(n8035), .ZN(n8044) );
  NAND2_X1 U8989 ( .A1(n10429), .A2(n8038), .ZN(n8041) );
  NAND2_X1 U8990 ( .A1(n10439), .A2(n8039), .ZN(n8040) );
  OAI21_X1 U8991 ( .B1(n8042), .B2(n8041), .A(n8040), .ZN(n8043) );
  AOI21_X1 U8992 ( .B1(n8045), .B2(n8044), .A(n8043), .ZN(n8046) );
  OAI21_X1 U8993 ( .B1(n8048), .B2(n8047), .A(n8046), .ZN(n8073) );
  NAND2_X1 U8994 ( .A1(n6212), .A2(n8049), .ZN(n8052) );
  NAND2_X1 U8995 ( .A1(n8807), .A2(n8050), .ZN(n8051) );
  OAI21_X1 U8996 ( .B1(n8053), .B2(n8052), .A(n8051), .ZN(n8060) );
  NAND2_X1 U8997 ( .A1(n6216), .A2(n8054), .ZN(n8057) );
  NAND2_X1 U8998 ( .A1(n8494), .A2(n8055), .ZN(n8056) );
  OAI21_X1 U8999 ( .B1(n8058), .B2(n8057), .A(n8056), .ZN(n8059) );
  AOI21_X1 U9000 ( .B1(n8061), .B2(n8060), .A(n8059), .ZN(n8070) );
  NAND2_X1 U9001 ( .A1(data_addr_o_31__BAR), .A2(n8062), .ZN(n8065) );
  INV_X1 U9002 ( .A(n8063), .ZN(n8064) );
  NAND2_X1 U9003 ( .A1(n8065), .A2(n8064), .ZN(n8067) );
  NOR2_X1 U9004 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  OAI21_X1 U9005 ( .B1(n8070), .B2(n8069), .A(n8068), .ZN(n8071) );
  AOI21_X1 U9006 ( .B1(n8073), .B2(n8072), .A(n8071), .ZN(n8074) );
  OAI21_X1 U9007 ( .B1(n8076), .B2(n8075), .A(n8074), .ZN(n8080) );
  INV_X1 U9008 ( .A(pmp_cfg_i[0]), .ZN(n8078) );
  NAND2_X1 U9009 ( .A1(n11019), .A2(pmp_cfg_i[1]), .ZN(n8077) );
  OAI21_X1 U9010 ( .B1(n8078), .B2(n11019), .A(n8077), .ZN(n11330) );
  NAND3_X1 U9011 ( .A1(n8080), .A2(n11330), .A3(n8079), .ZN(n8082) );
  AND2_X1 U9012 ( .A1(n8082), .A2(n8081), .ZN(n8083) );
  NAND4_X1 U9013 ( .A1(n8086), .A2(n8085), .A3(n8084), .A4(n8083), .ZN(n8087)
         );
  NOR2_X1 U9014 ( .A1(n8088), .A2(n8087), .ZN(n9340) );
  NOR2_X1 U9015 ( .A1(n10047), .A2(pmp_addr_i[46]), .ZN(n8090) );
  NOR2_X1 U9016 ( .A1(n8757), .A2(pmp_addr_i[47]), .ZN(n8136) );
  NOR2_X1 U9017 ( .A1(n8090), .A2(n8136), .ZN(n8139) );
  NOR2_X1 U9018 ( .A1(pmp_addr_i[44]), .A2(n10000), .ZN(n8091) );
  NOR2_X1 U9019 ( .A1(pmp_addr_i[45]), .A2(n10721), .ZN(n8133) );
  NOR2_X1 U9020 ( .A1(n8091), .A2(n8133), .ZN(n8092) );
  NAND2_X1 U9021 ( .A1(n8139), .A2(n8092), .ZN(n8142) );
  NOR2_X1 U9022 ( .A1(pmp_addr_i[41]), .A2(n10711), .ZN(n8124) );
  NOR2_X1 U9023 ( .A1(pmp_addr_i[40]), .A2(n6141), .ZN(n8093) );
  NOR2_X1 U9024 ( .A1(n8124), .A2(n8093), .ZN(n8095) );
  NOR2_X1 U9025 ( .A1(pmp_addr_i[42]), .A2(n10005), .ZN(n8094) );
  NOR2_X1 U9026 ( .A1(pmp_addr_i[43]), .A2(n10342), .ZN(n8127) );
  NOR2_X1 U9027 ( .A1(n8094), .A2(n8127), .ZN(n8130) );
  NAND2_X1 U9028 ( .A1(n8095), .A2(n8130), .ZN(n8096) );
  NOR2_X1 U9029 ( .A1(n8142), .A2(n8096), .ZN(n8145) );
  NOR2_X1 U9030 ( .A1(pmp_addr_i[34]), .A2(n10351), .ZN(n8097) );
  NOR2_X1 U9031 ( .A1(pmp_addr_i[35]), .A2(n10346), .ZN(n8103) );
  NOR2_X1 U9032 ( .A1(n8097), .A2(n8103), .ZN(n8106) );
  NOR2_X1 U9033 ( .A1(pmp_addr_i[33]), .A2(n9350), .ZN(n8100) );
  NAND2_X1 U9034 ( .A1(pmp_addr_i[32]), .A2(n10651), .ZN(n8099) );
  NAND2_X1 U9035 ( .A1(pmp_addr_i[33]), .A2(n9350), .ZN(n8098) );
  OAI21_X1 U9036 ( .B1(n8100), .B2(n8099), .A(n8098), .ZN(n8105) );
  NAND2_X1 U9037 ( .A1(pmp_addr_i[34]), .A2(n10351), .ZN(n8102) );
  NAND2_X1 U9038 ( .A1(pmp_addr_i[35]), .A2(n6127), .ZN(n8101) );
  OAI21_X1 U9039 ( .B1(n8103), .B2(n8102), .A(n8101), .ZN(n8104) );
  AOI21_X1 U9040 ( .B1(n8106), .B2(n8105), .A(n8104), .ZN(n8121) );
  NOR2_X1 U9041 ( .A1(n8735), .A2(pmp_addr_i[38]), .ZN(n8107) );
  NOR2_X1 U9042 ( .A1(pmp_addr_i[39]), .A2(n9367), .ZN(n8115) );
  NOR2_X1 U9043 ( .A1(n8107), .A2(n8115), .ZN(n8118) );
  NOR2_X1 U9044 ( .A1(pmp_addr_i[36]), .A2(n9363), .ZN(n8108) );
  NOR2_X1 U9045 ( .A1(pmp_addr_i[37]), .A2(n10697), .ZN(n8112) );
  NOR2_X1 U9046 ( .A1(n8108), .A2(n8112), .ZN(n8109) );
  NAND2_X1 U9047 ( .A1(n8118), .A2(n8109), .ZN(n8120) );
  NAND2_X1 U9048 ( .A1(pmp_addr_i[36]), .A2(n9363), .ZN(n8111) );
  NAND2_X1 U9049 ( .A1(pmp_addr_i[37]), .A2(n10697), .ZN(n8110) );
  OAI21_X1 U9050 ( .B1(n8112), .B2(n8111), .A(n8110), .ZN(n8117) );
  NAND2_X1 U9051 ( .A1(n8735), .A2(pmp_addr_i[38]), .ZN(n8114) );
  NAND2_X1 U9052 ( .A1(pmp_addr_i[39]), .A2(n10501), .ZN(n8113) );
  OAI21_X1 U9053 ( .B1(n8115), .B2(n8114), .A(n8113), .ZN(n8116) );
  AOI21_X1 U9054 ( .B1(n8118), .B2(n8117), .A(n8116), .ZN(n8119) );
  OAI21_X1 U9055 ( .B1(n8121), .B2(n8120), .A(n8119), .ZN(n8144) );
  NAND2_X1 U9056 ( .A1(pmp_addr_i[40]), .A2(n10701), .ZN(n8123) );
  NAND2_X1 U9057 ( .A1(pmp_addr_i[41]), .A2(n9508), .ZN(n8122) );
  OAI21_X1 U9058 ( .B1(n8124), .B2(n8123), .A(n8122), .ZN(n8129) );
  NAND2_X1 U9059 ( .A1(pmp_addr_i[42]), .A2(n10005), .ZN(n8126) );
  NAND2_X1 U9060 ( .A1(pmp_addr_i[43]), .A2(n11006), .ZN(n8125) );
  OAI21_X1 U9061 ( .B1(n8127), .B2(n8126), .A(n8125), .ZN(n8128) );
  AOI21_X1 U9062 ( .B1(n8130), .B2(n8129), .A(n8128), .ZN(n8141) );
  NAND2_X1 U9063 ( .A1(pmp_addr_i[44]), .A2(n6154), .ZN(n8132) );
  NAND2_X1 U9064 ( .A1(pmp_addr_i[45]), .A2(n10338), .ZN(n8131) );
  OAI21_X1 U9065 ( .B1(n8133), .B2(n8132), .A(n8131), .ZN(n8138) );
  NAND2_X1 U9066 ( .A1(n7057), .A2(pmp_addr_i[46]), .ZN(n8135) );
  NAND2_X1 U9067 ( .A1(n8757), .A2(pmp_addr_i[47]), .ZN(n8134) );
  OAI21_X1 U9068 ( .B1(n8136), .B2(n8135), .A(n8134), .ZN(n8137) );
  AOI21_X1 U9069 ( .B1(n8139), .B2(n8138), .A(n8137), .ZN(n8140) );
  OAI21_X1 U9070 ( .B1(n8142), .B2(n8141), .A(n8140), .ZN(n8143) );
  AOI21_X1 U9071 ( .B1(n8145), .B2(n8144), .A(n8143), .ZN(n8203) );
  NOR2_X1 U9072 ( .A1(n9425), .A2(pmp_addr_i[52]), .ZN(n8146) );
  NOR2_X1 U9073 ( .A1(n10424), .A2(pmp_addr_i[53]), .ZN(n8170) );
  NOR2_X1 U9074 ( .A1(n8146), .A2(n8170), .ZN(n8148) );
  NOR2_X1 U9075 ( .A1(n10428), .A2(pmp_addr_i[54]), .ZN(n8147) );
  NOR2_X1 U9076 ( .A1(n10429), .A2(pmp_addr_i[55]), .ZN(n8173) );
  NOR2_X1 U9077 ( .A1(n8147), .A2(n8173), .ZN(n8176) );
  NAND2_X1 U9078 ( .A1(n8148), .A2(n8176), .ZN(n8178) );
  NOR2_X1 U9079 ( .A1(n9418), .A2(pmp_addr_i[51]), .ZN(n8164) );
  NOR2_X1 U9080 ( .A1(n10754), .A2(pmp_addr_i[50]), .ZN(n8149) );
  NOR2_X1 U9081 ( .A1(n8164), .A2(n8149), .ZN(n8167) );
  NOR2_X1 U9082 ( .A1(n9414), .A2(pmp_addr_i[49]), .ZN(n8161) );
  NOR2_X1 U9083 ( .A1(n10060), .A2(pmp_addr_i[48]), .ZN(n8150) );
  NOR2_X1 U9084 ( .A1(n8161), .A2(n8150), .ZN(n8151) );
  NAND2_X1 U9085 ( .A1(n8167), .A2(n8151), .ZN(n8152) );
  NOR2_X1 U9086 ( .A1(n8178), .A2(n8152), .ZN(n8158) );
  NOR2_X1 U9087 ( .A1(n10439), .A2(pmp_addr_i[56]), .ZN(n8153) );
  NOR2_X1 U9088 ( .A1(n9438), .A2(pmp_addr_i[57]), .ZN(n8182) );
  NOR2_X1 U9089 ( .A1(n8153), .A2(n8182), .ZN(n8155) );
  NOR2_X1 U9090 ( .A1(n10778), .A2(pmp_addr_i[58]), .ZN(n8154) );
  NOR2_X1 U9091 ( .A1(n10782), .A2(pmp_addr_i[59]), .ZN(n8185) );
  NOR2_X1 U9092 ( .A1(n8154), .A2(n8185), .ZN(n8188) );
  NAND2_X1 U9093 ( .A1(n8155), .A2(n8188), .ZN(n8157) );
  NOR2_X1 U9095 ( .A1(n8494), .A2(pmp_addr_i[60]), .ZN(n8156) );
  NOR2_X1 U9096 ( .A1(n10107), .A2(pmp_addr_i[61]), .ZN(n8192) );
  OR2_X1 U9097 ( .A1(n8156), .A2(n8192), .ZN(n8196) );
  NOR2_X1 U9098 ( .A1(n8157), .A2(n8196), .ZN(n8199) );
  NAND2_X1 U9099 ( .A1(n8158), .A2(n8199), .ZN(n8202) );
  NAND2_X1 U9100 ( .A1(n10060), .A2(pmp_addr_i[48]), .ZN(n8160) );
  NAND2_X1 U9101 ( .A1(n10414), .A2(pmp_addr_i[49]), .ZN(n8159) );
  OAI21_X1 U9102 ( .B1(n8161), .B2(n8160), .A(n8159), .ZN(n8166) );
  NAND2_X1 U9103 ( .A1(n10754), .A2(pmp_addr_i[50]), .ZN(n8163) );
  NAND2_X1 U9104 ( .A1(n6192), .A2(pmp_addr_i[51]), .ZN(n8162) );
  OAI21_X1 U9105 ( .B1(n8164), .B2(n8163), .A(n8162), .ZN(n8165) );
  AOI21_X1 U9106 ( .B1(n8167), .B2(n8166), .A(n8165), .ZN(n8179) );
  NAND2_X1 U9107 ( .A1(n9425), .A2(pmp_addr_i[52]), .ZN(n8169) );
  NAND2_X1 U9108 ( .A1(n10424), .A2(pmp_addr_i[53]), .ZN(n8168) );
  OAI21_X1 U9109 ( .B1(n8170), .B2(n8169), .A(n8168), .ZN(n8175) );
  NAND2_X1 U9110 ( .A1(n10428), .A2(pmp_addr_i[54]), .ZN(n8172) );
  NAND2_X1 U9111 ( .A1(n6462), .A2(pmp_addr_i[55]), .ZN(n8171) );
  OAI21_X1 U9112 ( .B1(n8173), .B2(n8172), .A(n8171), .ZN(n8174) );
  AOI21_X1 U9113 ( .B1(n8176), .B2(n8175), .A(n8174), .ZN(n8177) );
  OAI21_X1 U9114 ( .B1(n8179), .B2(n8178), .A(n8177), .ZN(n8200) );
  NAND2_X1 U9115 ( .A1(n10439), .A2(pmp_addr_i[56]), .ZN(n8181) );
  NAND2_X1 U9116 ( .A1(n9438), .A2(pmp_addr_i[57]), .ZN(n8180) );
  OAI21_X1 U9117 ( .B1(n8182), .B2(n8181), .A(n8180), .ZN(n8187) );
  NAND2_X1 U9118 ( .A1(n10778), .A2(pmp_addr_i[58]), .ZN(n8184) );
  NAND2_X1 U9119 ( .A1(n6216), .A2(pmp_addr_i[59]), .ZN(n8183) );
  OAI21_X1 U9120 ( .B1(n8185), .B2(n8184), .A(n8183), .ZN(n8186) );
  AOI21_X1 U9121 ( .B1(n8188), .B2(n8187), .A(n8186), .ZN(n8197) );
  NAND2_X1 U9122 ( .A1(n8494), .A2(pmp_addr_i[60]), .ZN(n8191) );
  NAND2_X1 U9123 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[61]), .ZN(n8190)
         );
  OAI21_X1 U9124 ( .B1(n8192), .B2(n8191), .A(n8190), .ZN(n8194) );
  NOR2_X1 U9125 ( .A1(n8194), .A2(n2028), .ZN(n8195) );
  OAI21_X1 U9126 ( .B1(n8197), .B2(n8196), .A(n8195), .ZN(n8198) );
  AOI21_X1 U9127 ( .B1(n8200), .B2(n8199), .A(n8198), .ZN(n8201) );
  OAI21_X1 U9128 ( .B1(n8203), .B2(n8202), .A(n8201), .ZN(n8324) );
  NOR2_X1 U9129 ( .A1(n10335), .A2(n325), .ZN(n8253) );
  NOR2_X1 U9130 ( .A1(data_addr_o_15_), .A2(n8326), .ZN(n8205) );
  NOR2_X1 U9131 ( .A1(n8253), .A2(n8205), .ZN(n8207) );
  NOR2_X1 U9132 ( .A1(n10857), .A2(n2719), .ZN(n8256) );
  NAND2_X1 U9133 ( .A1(n7995), .A2(n8254), .ZN(n8344) );
  INV_X1 U9134 ( .A(n8344), .ZN(n8206) );
  NOR2_X1 U9135 ( .A1(n8256), .A2(n8206), .ZN(n8259) );
  NAND2_X1 U9136 ( .A1(n8207), .A2(n8259), .ZN(n8262) );
  NOR2_X1 U9137 ( .A1(n8246), .A2(n326), .ZN(n8209) );
  NOR2_X1 U9138 ( .A1(data_addr_o_12_), .A2(n8341), .ZN(n8247) );
  NOR2_X1 U9139 ( .A1(n8209), .A2(n8247), .ZN(n8213) );
  NOR2_X1 U9140 ( .A1(n10847), .A2(n8340), .ZN(n8212) );
  NOR2_X1 U9141 ( .A1(n10848), .A2(n8325), .ZN(n8248) );
  NOR2_X1 U9142 ( .A1(n8212), .A2(n8248), .ZN(n8251) );
  NAND2_X1 U9143 ( .A1(n8213), .A2(n8251), .ZN(n8214) );
  NOR2_X1 U9144 ( .A1(n8262), .A2(n8214), .ZN(n8265) );
  OAI22_X1 U9145 ( .A1(n8379), .A2(data_addr_o_5_), .B1(n10358), .B2(n327), 
        .ZN(n8337) );
  INV_X1 U9146 ( .A(n8337), .ZN(n8227) );
  INV_X1 U9147 ( .A(n8381), .ZN(n8215) );
  OR2_X1 U9148 ( .A1(data_addr_o_2_), .A2(n8215), .ZN(n8218) );
  NAND2_X1 U9149 ( .A1(n10473), .A2(n8380), .ZN(n8333) );
  INV_X1 U9150 ( .A(n8380), .ZN(n8216) );
  AND2_X1 U9151 ( .A1(n22), .A2(n8216), .ZN(n8217) );
  AOI21_X1 U9152 ( .B1(n8218), .B2(n8333), .A(n8217), .ZN(n8221) );
  NOR2_X1 U9153 ( .A1(n10135), .A2(n8334), .ZN(n8220) );
  NAND2_X1 U9154 ( .A1(n10479), .A2(n8334), .ZN(n11485) );
  OAI21_X1 U9155 ( .B1(n8221), .B2(n8220), .A(n11485), .ZN(n8226) );
  NOR2_X1 U9156 ( .A1(data_addr_o_6_), .A2(n327), .ZN(n8224) );
  NAND2_X1 U9157 ( .A1(n10486), .A2(n8379), .ZN(n8223) );
  NAND2_X1 U9158 ( .A1(data_addr_o_6_), .A2(n327), .ZN(n11475) );
  OAI21_X1 U9159 ( .B1(n8224), .B2(n8223), .A(n11475), .ZN(n8225) );
  AOI21_X1 U9160 ( .B1(n8227), .B2(n8226), .A(n8225), .ZN(n8245) );
  OAI22_X1 U9161 ( .A1(n8229), .A2(n11343), .B1(data_addr_o_9_), .B2(n8228), 
        .ZN(n8328) );
  INV_X1 U9162 ( .A(n8328), .ZN(n8242) );
  NOR2_X1 U9163 ( .A1(n10494), .A2(n8339), .ZN(n8234) );
  NOR2_X1 U9164 ( .A1(data_addr_o_7_), .A2(n4989), .ZN(n8336) );
  NOR2_X1 U9165 ( .A1(n8234), .A2(n8336), .ZN(n8232) );
  NAND2_X1 U9166 ( .A1(n8242), .A2(n8232), .ZN(n8244) );
  NAND2_X1 U9167 ( .A1(data_addr_o_7_), .A2(n4989), .ZN(n11474) );
  NAND2_X1 U9168 ( .A1(n9805), .A2(n8339), .ZN(n8378) );
  OAI21_X1 U9169 ( .B1(n8234), .B2(n11474), .A(n8378), .ZN(n8241) );
  NOR2_X1 U9170 ( .A1(n8238), .A2(n8229), .ZN(n8239) );
  NAND2_X1 U9171 ( .A1(n8237), .A2(n8228), .ZN(n11494) );
  NAND2_X1 U9172 ( .A1(n8238), .A2(n8229), .ZN(n11495) );
  OAI21_X1 U9173 ( .B1(n8239), .B2(n11494), .A(n11495), .ZN(n8240) );
  AOI21_X1 U9174 ( .B1(n8242), .B2(n8241), .A(n8240), .ZN(n8243) );
  OAI21_X1 U9175 ( .B1(n8245), .B2(n8244), .A(n8243), .ZN(n8264) );
  NAND2_X1 U9176 ( .A1(n8246), .A2(n326), .ZN(n11507) );
  NAND2_X1 U9177 ( .A1(data_addr_o_12_), .A2(n8341), .ZN(n11464) );
  OAI21_X1 U9178 ( .B1(n8247), .B2(n11507), .A(n11464), .ZN(n8250) );
  NAND2_X1 U9179 ( .A1(n10847), .A2(n8340), .ZN(n11501) );
  NAND2_X1 U9180 ( .A1(n10848), .A2(n8325), .ZN(n11491) );
  OAI21_X1 U9181 ( .B1(n8248), .B2(n11501), .A(n11491), .ZN(n8249) );
  AOI21_X1 U9182 ( .B1(n8251), .B2(n8250), .A(n8249), .ZN(n8261) );
  NAND2_X1 U9183 ( .A1(data_addr_o_15_), .A2(n8326), .ZN(n11468) );
  NAND2_X1 U9184 ( .A1(n10335), .A2(n325), .ZN(n8252) );
  OAI21_X1 U9185 ( .B1(n8253), .B2(n11468), .A(n8252), .ZN(n8258) );
  NAND2_X1 U9186 ( .A1(n6813), .A2(n5000), .ZN(n11500) );
  NAND2_X1 U9187 ( .A1(n10857), .A2(n2719), .ZN(n8255) );
  OAI21_X1 U9188 ( .B1(n8256), .B2(n11500), .A(n8255), .ZN(n8257) );
  AOI21_X1 U9189 ( .B1(n8259), .B2(n8258), .A(n8257), .ZN(n8260) );
  OAI21_X1 U9190 ( .B1(n8262), .B2(n8261), .A(n8260), .ZN(n8263) );
  AOI21_X1 U9191 ( .B1(n8265), .B2(n8264), .A(n8263), .ZN(n8322) );
  NOR2_X1 U9192 ( .A1(n10898), .A2(n2810), .ZN(n8266) );
  NOR2_X1 U9193 ( .A1(n10738), .A2(n2795), .ZN(n8292) );
  NOR2_X1 U9194 ( .A1(n8266), .A2(n8292), .ZN(n8268) );
  NOR2_X1 U9195 ( .A1(n10903), .A2(n2813), .ZN(n8267) );
  NOR2_X1 U9196 ( .A1(n10267), .A2(n2787), .ZN(n8295) );
  NOR2_X1 U9197 ( .A1(n8267), .A2(n8295), .ZN(n8298) );
  NAND2_X1 U9198 ( .A1(n8268), .A2(n8298), .ZN(n8300) );
  NOR2_X1 U9199 ( .A1(n11312), .A2(n2801), .ZN(n8269) );
  NOR2_X1 U9200 ( .A1(n9529), .A2(n2779), .ZN(n8286) );
  NOR2_X1 U9201 ( .A1(n8269), .A2(n8286), .ZN(n8289) );
  NOR2_X1 U9202 ( .A1(n9846), .A2(n2798), .ZN(n8270) );
  NOR2_X1 U9203 ( .A1(data_addr_o_20_), .A2(n2776), .ZN(n8283) );
  NOR2_X1 U9204 ( .A1(n8270), .A2(n8283), .ZN(n8271) );
  NAND2_X1 U9205 ( .A1(n8289), .A2(n8271), .ZN(n8272) );
  NOR2_X1 U9206 ( .A1(n8300), .A2(n8272), .ZN(n8280) );
  NOR2_X1 U9207 ( .A1(n9886), .A2(n2826), .ZN(n8273) );
  INV_X1 U9208 ( .A(n8360), .ZN(n8302) );
  NOR2_X1 U9209 ( .A1(n10635), .A2(n8302), .ZN(n8305) );
  NOR2_X1 U9210 ( .A1(n8273), .A2(n8305), .ZN(n8275) );
  NOR2_X1 U9211 ( .A1(n10918), .A2(n2829), .ZN(n8274) );
  NOR2_X1 U9212 ( .A1(data_addr_o_30_), .A2(n2830), .ZN(n8308) );
  NOR2_X1 U9213 ( .A1(n8274), .A2(n8308), .ZN(n8311) );
  NAND2_X1 U9214 ( .A1(n8275), .A2(n8311), .ZN(n8279) );
  NOR2_X1 U9215 ( .A1(n24), .A2(n8385), .ZN(n8277) );
  NOR2_X1 U9216 ( .A1(n8277), .A2(pmp_addr_i[30]), .ZN(n8278) );
  NAND2_X1 U9217 ( .A1(n8278), .A2(n2760), .ZN(n8315) );
  NOR2_X1 U9218 ( .A1(n8279), .A2(n8315), .ZN(n8318) );
  NAND2_X1 U9219 ( .A1(n8280), .A2(n8318), .ZN(n8321) );
  NAND2_X1 U9220 ( .A1(n9846), .A2(n2798), .ZN(n8282) );
  NAND2_X1 U9221 ( .A1(n10887), .A2(n2776), .ZN(n8281) );
  OAI21_X1 U9222 ( .B1(n8283), .B2(n8282), .A(n8281), .ZN(n8288) );
  NAND2_X1 U9223 ( .A1(n11312), .A2(n2801), .ZN(n8285) );
  NAND2_X1 U9224 ( .A1(n9529), .A2(n2779), .ZN(n8284) );
  OAI21_X1 U9225 ( .B1(n8286), .B2(n8285), .A(n8284), .ZN(n8287) );
  AOI21_X1 U9226 ( .B1(n8289), .B2(n8288), .A(n8287), .ZN(n8301) );
  NAND2_X1 U9227 ( .A1(data_addr_o_23_), .A2(n2810), .ZN(n8291) );
  NAND2_X1 U9228 ( .A1(n10899), .A2(n2795), .ZN(n8290) );
  OAI21_X1 U9229 ( .B1(n8292), .B2(n8291), .A(n8290), .ZN(n8297) );
  NAND2_X1 U9230 ( .A1(n10903), .A2(n2813), .ZN(n8294) );
  NAND2_X1 U9231 ( .A1(n10267), .A2(n2787), .ZN(n8293) );
  OAI21_X1 U9232 ( .B1(n8295), .B2(n8294), .A(n8293), .ZN(n8296) );
  AOI21_X1 U9233 ( .B1(n8298), .B2(n8297), .A(n8296), .ZN(n8299) );
  OAI21_X1 U9234 ( .B1(n8301), .B2(n8300), .A(n8299), .ZN(n8319) );
  NAND2_X1 U9235 ( .A1(n9886), .A2(n2826), .ZN(n8304) );
  NAND2_X1 U9236 ( .A1(n10635), .A2(n8302), .ZN(n8303) );
  OAI21_X1 U9237 ( .B1(n8305), .B2(n8304), .A(n8303), .ZN(n8310) );
  NAND2_X1 U9238 ( .A1(n10918), .A2(n2829), .ZN(n8307) );
  NAND2_X1 U9239 ( .A1(data_addr_o_30_), .A2(n2830), .ZN(n8306) );
  OAI21_X1 U9240 ( .B1(n8308), .B2(n8307), .A(n8306), .ZN(n8309) );
  AOI21_X1 U9241 ( .B1(n8311), .B2(n8310), .A(n8309), .ZN(n8316) );
  NAND2_X1 U9242 ( .A1(n24), .A2(n8385), .ZN(n8312) );
  NOR2_X1 U9243 ( .A1(n8312), .A2(pmp_addr_i[30]), .ZN(n8313) );
  NAND2_X1 U9244 ( .A1(n8313), .A2(n2760), .ZN(n8314) );
  OAI21_X1 U9245 ( .B1(n8316), .B2(n8315), .A(n8314), .ZN(n8317) );
  AOI21_X1 U9246 ( .B1(n8319), .B2(n8318), .A(n8317), .ZN(n8320) );
  OAI21_X1 U9247 ( .B1(n8322), .B2(n8321), .A(n8320), .ZN(n8323) );
  NAND3_X1 U9248 ( .A1(n8324), .A2(n36), .A3(n8323), .ZN(n8394) );
  OAI22_X1 U9249 ( .A1(n9987), .A2(n325), .B1(n326), .B2(data_addr_o_11_), 
        .ZN(n8329) );
  OAI22_X1 U9250 ( .A1(n8326), .A2(data_addr_o_15_), .B1(data_addr_o_14_), 
        .B2(n8325), .ZN(n8327) );
  NOR3_X1 U9251 ( .A1(n8329), .A2(n8328), .A3(n8327), .ZN(n8347) );
  XNOR2_X1 U9252 ( .A(n11303), .B(n8330), .ZN(n8346) );
  INV_X1 U9253 ( .A(pmp_cfg_i[12]), .ZN(n8331) );
  AOI21_X1 U9254 ( .B1(n8695), .B2(n8381), .A(n8331), .ZN(n8332) );
  OAI211_X1 U9255 ( .C1(n8334), .C2(n11288), .A(n8333), .B(n8332), .ZN(n8335)
         );
  NOR2_X1 U9256 ( .A1(n8336), .A2(n8335), .ZN(n8338) );
  OAI211_X1 U9257 ( .C1(n8339), .C2(n10281), .A(n8338), .B(n8227), .ZN(n8343)
         );
  OAI22_X1 U9258 ( .A1(n8341), .A2(n31), .B1(data_addr_o_13_), .B2(n8340), 
        .ZN(n8342) );
  NOR2_X1 U9259 ( .A1(n8343), .A2(n8342), .ZN(n8345) );
  NAND4_X1 U9260 ( .A1(n8347), .A2(n8346), .A3(n8345), .A4(n8344), .ZN(n8357)
         );
  XNOR2_X1 U9261 ( .A(n10627), .B(n8348), .ZN(n8355) );
  XNOR2_X1 U9262 ( .A(n11285), .B(n8349), .ZN(n8354) );
  XNOR2_X1 U9263 ( .A(n10638), .B(n8350), .ZN(n8353) );
  XNOR2_X1 U9264 ( .A(n10898), .B(n8351), .ZN(n8352) );
  NAND4_X1 U9265 ( .A1(n8355), .A2(n8354), .A3(n8353), .A4(n8352), .ZN(n8356)
         );
  NOR2_X1 U9266 ( .A1(n8357), .A2(n8356), .ZN(n8377) );
  XNOR2_X1 U9267 ( .A(n10614), .B(n8358), .ZN(n8365) );
  XNOR2_X1 U9268 ( .A(n10606), .B(n8359), .ZN(n8364) );
  XNOR2_X1 U9269 ( .A(n10635), .B(n8360), .ZN(n8363) );
  XNOR2_X1 U9270 ( .A(data_addr_o_30_), .B(n8361), .ZN(n8362) );
  NAND4_X1 U9271 ( .A1(n8365), .A2(n8364), .A3(n8363), .A4(n8362), .ZN(n8375)
         );
  XNOR2_X1 U9272 ( .A(n10967), .B(n8366), .ZN(n8373) );
  XNOR2_X1 U9273 ( .A(n10612), .B(n8367), .ZN(n8372) );
  XNOR2_X1 U9274 ( .A(n10629), .B(n8368), .ZN(n8371) );
  XNOR2_X1 U9275 ( .A(n10616), .B(n8369), .ZN(n8370) );
  NAND4_X1 U9276 ( .A1(n8373), .A2(n8372), .A3(n8371), .A4(n8370), .ZN(n8374)
         );
  NOR2_X1 U9277 ( .A1(n8375), .A2(n8374), .ZN(n8376) );
  AND2_X1 U9278 ( .A1(n8377), .A2(n8376), .ZN(n11517) );
  NAND4_X1 U9279 ( .A1(n11468), .A2(n11494), .A3(n11495), .A4(n8378), .ZN(
        n11513) );
  INV_X1 U9280 ( .A(n11513), .ZN(n8390) );
  AND2_X1 U9281 ( .A1(n10335), .A2(n325), .ZN(n11463) );
  AND2_X1 U9282 ( .A1(n10824), .A2(n8379), .ZN(n11488) );
  NAND2_X1 U9283 ( .A1(n22), .A2(n8216), .ZN(n11481) );
  OAI211_X1 U9284 ( .C1(n8381), .C2(n8695), .A(n11485), .B(n11481), .ZN(n8382)
         );
  NOR2_X1 U9285 ( .A1(n11488), .A2(n8382), .ZN(n8383) );
  NAND4_X1 U9286 ( .A1(n11491), .A2(n8383), .A3(n11475), .A4(n11474), .ZN(
        n8384) );
  NOR2_X1 U9287 ( .A1(n11463), .A2(n8384), .ZN(n8389) );
  NAND4_X1 U9288 ( .A1(n11500), .A2(n11464), .A3(n11507), .A4(n11501), .ZN(
        n8387) );
  XNOR2_X1 U9289 ( .A(n12123), .B(n8385), .ZN(n8386) );
  NOR2_X1 U9290 ( .A1(n8387), .A2(n8386), .ZN(n8388) );
  NAND4_X1 U9291 ( .A1(n11517), .A2(n8390), .A3(n8389), .A4(n8388), .ZN(n8393)
         );
  MUX2_X1 U9292 ( .A(pmp_cfg_i[8]), .B(pmp_cfg_i[9]), .S(n11019), .Z(n8392) );
  NAND2_X1 U9293 ( .A1(n8391), .A2(n8392), .ZN(n11504) );
  AOI21_X1 U9294 ( .B1(n8394), .B2(n8393), .A(n11504), .ZN(n8711) );
  NOR2_X1 U9295 ( .A1(n7990), .A2(pmp_addr_i[398]), .ZN(n8443) );
  NOR2_X1 U9296 ( .A1(n10721), .A2(pmp_addr_i[397]), .ZN(n8395) );
  NOR2_X1 U9297 ( .A1(n8443), .A2(n8395), .ZN(n8397) );
  NOR2_X1 U9299 ( .A1(n12184), .A2(pmp_addr_i[400]), .ZN(n8448) );
  INV_X1 U9300 ( .A(data_addr_i[17]), .ZN(n8444) );
  NOR2_X1 U9301 ( .A1(n8444), .A2(pmp_addr_i[399]), .ZN(n8396) );
  NOR2_X1 U9302 ( .A1(n8448), .A2(n8396), .ZN(n8450) );
  NAND2_X1 U9303 ( .A1(n8397), .A2(n8450), .ZN(n8454) );
  NOR2_X1 U9304 ( .A1(n9508), .A2(pmp_addr_i[393]), .ZN(n8398) );
  NOR2_X1 U9305 ( .A1(n9947), .A2(pmp_addr_i[394]), .ZN(n8434) );
  NOR2_X1 U9306 ( .A1(n8398), .A2(n8434), .ZN(n8400) );
  NOR2_X1 U9307 ( .A1(n11006), .A2(pmp_addr_i[395]), .ZN(n8399) );
  NOR2_X1 U9308 ( .A1(n6154), .A2(pmp_addr_i[396]), .ZN(n8437) );
  NOR2_X1 U9309 ( .A1(n8399), .A2(n8437), .ZN(n8440) );
  NAND2_X1 U9310 ( .A1(n8400), .A2(n8440), .ZN(n8401) );
  NOR2_X1 U9311 ( .A1(n8454), .A2(n8401), .ZN(n8457) );
  NOR2_X1 U9312 ( .A1(n6127), .A2(pmp_addr_i[387]), .ZN(n8402) );
  INV_X1 U9313 ( .A(n10655), .ZN(n8410) );
  NOR2_X1 U9314 ( .A1(n8410), .A2(pmp_addr_i[388]), .ZN(n8413) );
  NOR2_X1 U9315 ( .A1(n8402), .A2(n8413), .ZN(n8416) );
  OR2_X1 U9316 ( .A1(n10010), .A2(pmp_addr_i[385]), .ZN(n8405) );
  AND2_X1 U9317 ( .A1(n10651), .A2(pmp_addr_i[384]), .ZN(n8404) );
  AND2_X1 U9318 ( .A1(n10010), .A2(pmp_addr_i[385]), .ZN(n8403) );
  AOI21_X1 U9319 ( .B1(n8405), .B2(n8404), .A(n8403), .ZN(n8409) );
  INV_X1 U9320 ( .A(n10479), .ZN(n8406) );
  NOR2_X1 U9321 ( .A1(n8406), .A2(pmp_addr_i[386]), .ZN(n8408) );
  NAND2_X1 U9322 ( .A1(n8406), .A2(pmp_addr_i[386]), .ZN(n8407) );
  OAI21_X1 U9323 ( .B1(n8409), .B2(n8408), .A(n8407), .ZN(n8415) );
  NAND2_X1 U9324 ( .A1(n6127), .A2(pmp_addr_i[387]), .ZN(n8412) );
  NAND2_X1 U9325 ( .A1(n8410), .A2(pmp_addr_i[388]), .ZN(n8411) );
  OAI21_X1 U9326 ( .B1(n8413), .B2(n8412), .A(n8411), .ZN(n8414) );
  AOI21_X1 U9327 ( .B1(n8416), .B2(n8415), .A(n8414), .ZN(n8431) );
  NOR2_X1 U9328 ( .A1(n8735), .A2(pmp_addr_i[390]), .ZN(n8422) );
  NOR2_X1 U9329 ( .A1(n6400), .A2(pmp_addr_i[389]), .ZN(n8417) );
  NOR2_X1 U9330 ( .A1(n8422), .A2(n8417), .ZN(n8419) );
  NOR2_X1 U9331 ( .A1(n6140), .A2(pmp_addr_i[391]), .ZN(n8418) );
  NOR2_X1 U9332 ( .A1(n6141), .A2(pmp_addr_i[392]), .ZN(n8425) );
  NOR2_X1 U9333 ( .A1(n8418), .A2(n8425), .ZN(n8428) );
  NAND2_X1 U9334 ( .A1(n8419), .A2(n8428), .ZN(n8430) );
  NAND2_X1 U9335 ( .A1(n6400), .A2(pmp_addr_i[389]), .ZN(n8421) );
  NAND2_X1 U9336 ( .A1(n8735), .A2(pmp_addr_i[390]), .ZN(n8420) );
  OAI21_X1 U9337 ( .B1(n8422), .B2(n8421), .A(n8420), .ZN(n8427) );
  NAND2_X1 U9338 ( .A1(n10501), .A2(pmp_addr_i[391]), .ZN(n8424) );
  NAND2_X1 U9339 ( .A1(n10701), .A2(pmp_addr_i[392]), .ZN(n8423) );
  OAI21_X1 U9340 ( .B1(n8425), .B2(n8424), .A(n8423), .ZN(n8426) );
  AOI21_X1 U9341 ( .B1(n8428), .B2(n8427), .A(n8426), .ZN(n8429) );
  OAI21_X1 U9342 ( .B1(n8431), .B2(n8430), .A(n8429), .ZN(n8456) );
  NAND2_X1 U9343 ( .A1(n9508), .A2(pmp_addr_i[393]), .ZN(n8433) );
  NAND2_X1 U9344 ( .A1(n9947), .A2(pmp_addr_i[394]), .ZN(n8432) );
  OAI21_X1 U9345 ( .B1(n8434), .B2(n8433), .A(n8432), .ZN(n8439) );
  NAND2_X1 U9346 ( .A1(n11006), .A2(pmp_addr_i[395]), .ZN(n8436) );
  NAND2_X1 U9347 ( .A1(n6154), .A2(pmp_addr_i[396]), .ZN(n8435) );
  OAI21_X1 U9348 ( .B1(n8437), .B2(n8436), .A(n8435), .ZN(n8438) );
  AOI21_X1 U9349 ( .B1(n8440), .B2(n8439), .A(n8438), .ZN(n8453) );
  NAND2_X1 U9350 ( .A1(n9125), .A2(pmp_addr_i[397]), .ZN(n8442) );
  NAND2_X1 U9351 ( .A1(n10047), .A2(pmp_addr_i[398]), .ZN(n8441) );
  OAI21_X1 U9352 ( .B1(n8443), .B2(n8442), .A(n8441), .ZN(n8451) );
  NAND2_X1 U9353 ( .A1(n8444), .A2(pmp_addr_i[399]), .ZN(n8447) );
  NAND2_X1 U9354 ( .A1(n12184), .A2(pmp_addr_i[400]), .ZN(n8446) );
  OAI21_X1 U9355 ( .B1(n8448), .B2(n8447), .A(n8446), .ZN(n8449) );
  AOI21_X1 U9356 ( .B1(n8451), .B2(n8450), .A(n8449), .ZN(n8452) );
  OAI21_X1 U9357 ( .B1(n8454), .B2(n8453), .A(n8452), .ZN(n8455) );
  AOI21_X1 U9358 ( .B1(n8457), .B2(n8456), .A(n8455), .ZN(n8511) );
  NOR2_X1 U9359 ( .A1(n10424), .A2(pmp_addr_i[405]), .ZN(n8458) );
  NOR2_X1 U9360 ( .A1(n9163), .A2(pmp_addr_i[406]), .ZN(n8481) );
  NOR2_X1 U9361 ( .A1(n8458), .A2(n8481), .ZN(n8460) );
  NOR2_X1 U9362 ( .A1(n10429), .A2(pmp_addr_i[407]), .ZN(n8459) );
  NOR2_X1 U9363 ( .A1(n6202), .A2(pmp_addr_i[408]), .ZN(n8484) );
  NOR2_X1 U9364 ( .A1(n8459), .A2(n8484), .ZN(n8487) );
  NAND2_X1 U9365 ( .A1(n8460), .A2(n8487), .ZN(n8489) );
  NOR2_X1 U9366 ( .A1(n9418), .A2(pmp_addr_i[403]), .ZN(n8461) );
  NOR2_X1 U9367 ( .A1(n9156), .A2(pmp_addr_i[404]), .ZN(n8475) );
  NOR2_X1 U9368 ( .A1(n8461), .A2(n8475), .ZN(n8478) );
  NOR2_X1 U9369 ( .A1(n9414), .A2(pmp_addr_i[401]), .ZN(n8462) );
  NOR2_X1 U9370 ( .A1(n6188), .A2(pmp_addr_i[402]), .ZN(n8472) );
  NOR2_X1 U9371 ( .A1(n8462), .A2(n8472), .ZN(n8463) );
  NAND2_X1 U9372 ( .A1(n8478), .A2(n8463), .ZN(n8464) );
  NOR2_X1 U9373 ( .A1(n8489), .A2(n8464), .ZN(n8469) );
  NOR2_X1 U9374 ( .A1(n6212), .A2(pmp_addr_i[409]), .ZN(n8465) );
  NOR2_X1 U9375 ( .A1(n8807), .A2(pmp_addr_i[410]), .ZN(n8493) );
  NOR2_X1 U9376 ( .A1(n8465), .A2(n8493), .ZN(n8467) );
  NOR2_X1 U9377 ( .A1(n6216), .A2(pmp_addr_i[411]), .ZN(n8466) );
  INV_X1 U9378 ( .A(data_addr_i[30]), .ZN(n8494) );
  NOR2_X1 U9379 ( .A1(n8494), .A2(pmp_addr_i[412]), .ZN(n8497) );
  NOR2_X1 U9380 ( .A1(n8466), .A2(n8497), .ZN(n8500) );
  NAND2_X1 U9381 ( .A1(n8467), .A2(n8500), .ZN(n8468) );
  NOR2_X1 U9382 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[413]), .ZN(n8504)
         );
  NOR2_X1 U9383 ( .A1(n8468), .A2(n8504), .ZN(n8507) );
  NAND2_X1 U9384 ( .A1(n8469), .A2(n8507), .ZN(n8510) );
  NAND2_X1 U9385 ( .A1(n9414), .A2(pmp_addr_i[401]), .ZN(n8471) );
  NAND2_X1 U9386 ( .A1(n6188), .A2(pmp_addr_i[402]), .ZN(n8470) );
  OAI21_X1 U9387 ( .B1(n8472), .B2(n8471), .A(n8470), .ZN(n8477) );
  NAND2_X1 U9388 ( .A1(n6192), .A2(pmp_addr_i[403]), .ZN(n8474) );
  NAND2_X1 U9389 ( .A1(n9425), .A2(pmp_addr_i[404]), .ZN(n8473) );
  OAI21_X1 U9390 ( .B1(n8475), .B2(n8474), .A(n8473), .ZN(n8476) );
  AOI21_X1 U9391 ( .B1(n8478), .B2(n8477), .A(n8476), .ZN(n8490) );
  NAND2_X1 U9392 ( .A1(n10424), .A2(pmp_addr_i[405]), .ZN(n8480) );
  NAND2_X1 U9393 ( .A1(n10428), .A2(pmp_addr_i[406]), .ZN(n8479) );
  OAI21_X1 U9394 ( .B1(n8481), .B2(n8480), .A(n8479), .ZN(n8486) );
  NAND2_X1 U9395 ( .A1(n6462), .A2(pmp_addr_i[407]), .ZN(n8483) );
  NAND2_X1 U9396 ( .A1(n6202), .A2(pmp_addr_i[408]), .ZN(n8482) );
  OAI21_X1 U9397 ( .B1(n8484), .B2(n8483), .A(n8482), .ZN(n8485) );
  AOI21_X1 U9398 ( .B1(n8487), .B2(n8486), .A(n8485), .ZN(n8488) );
  OAI21_X1 U9399 ( .B1(n8490), .B2(n8489), .A(n8488), .ZN(n8508) );
  NAND2_X1 U9400 ( .A1(n6212), .A2(pmp_addr_i[409]), .ZN(n8492) );
  NAND2_X1 U9401 ( .A1(n10443), .A2(pmp_addr_i[410]), .ZN(n8491) );
  OAI21_X1 U9402 ( .B1(n8493), .B2(n8492), .A(n8491), .ZN(n8499) );
  NAND2_X1 U9403 ( .A1(n10782), .A2(pmp_addr_i[411]), .ZN(n8496) );
  NAND2_X1 U9404 ( .A1(n8494), .A2(pmp_addr_i[412]), .ZN(n8495) );
  OAI21_X1 U9405 ( .B1(n8497), .B2(n8496), .A(n8495), .ZN(n8498) );
  AOI21_X1 U9406 ( .B1(n8500), .B2(n8499), .A(n8498), .ZN(n8505) );
  NAND2_X1 U9407 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[413]), .ZN(n8501)
         );
  NAND2_X1 U9408 ( .A1(n8501), .A2(n4457), .ZN(n8502) );
  NOR2_X1 U9409 ( .A1(n8502), .A2(pmp_addr_i[415]), .ZN(n8503) );
  OAI21_X1 U9410 ( .B1(n8505), .B2(n8504), .A(n8503), .ZN(n8506) );
  AOI21_X1 U9411 ( .B1(n8508), .B2(n8507), .A(n8506), .ZN(n8509) );
  OAI21_X1 U9412 ( .B1(n8511), .B2(n8510), .A(n8509), .ZN(n8632) );
  NOR2_X1 U9413 ( .A1(data_addr_o_16_), .A2(n11409), .ZN(n8561) );
  NOR2_X1 U9414 ( .A1(n10657), .A2(n8678), .ZN(n8513) );
  NOR2_X1 U9415 ( .A1(n8561), .A2(n8513), .ZN(n8516) );
  NOR2_X1 U9417 ( .A1(n6813), .A2(n8691), .ZN(n8515) );
  NOR2_X1 U9418 ( .A1(n8564), .A2(n8515), .ZN(n8566) );
  NAND2_X1 U9419 ( .A1(n8516), .A2(n8566), .ZN(n8570) );
  NOR2_X1 U9420 ( .A1(data_addr_o_11_), .A2(n8671), .ZN(n8519) );
  INV_X1 U9421 ( .A(n9947), .ZN(n10499) );
  NOR2_X1 U9422 ( .A1(n10499), .A2(n8677), .ZN(n8555) );
  NOR2_X1 U9423 ( .A1(n8519), .A2(n8555), .ZN(n8522) );
  NOR2_X1 U9424 ( .A1(n10847), .A2(n8676), .ZN(n8521) );
  NOR2_X1 U9425 ( .A1(n10848), .A2(n8679), .ZN(n8557) );
  NOR2_X1 U9426 ( .A1(n8521), .A2(n8557), .ZN(n8560) );
  NAND2_X1 U9427 ( .A1(n8522), .A2(n8560), .ZN(n8523) );
  NOR2_X1 U9428 ( .A1(n8570), .A2(n8523), .ZN(n8573) );
  OAI22_X1 U9429 ( .A1(n8694), .A2(n10486), .B1(data_addr_o_6_), .B2(n8524), 
        .ZN(n8667) );
  INV_X1 U9430 ( .A(n8667), .ZN(n8539) );
  INV_X1 U9431 ( .A(n8696), .ZN(n8525) );
  OR2_X1 U9432 ( .A1(n10129), .A2(n8525), .ZN(n8529) );
  INV_X1 U9433 ( .A(n8660), .ZN(n8526) );
  OR2_X1 U9434 ( .A1(n10818), .A2(n8526), .ZN(n8528) );
  AND2_X1 U9435 ( .A1(n10130), .A2(n8526), .ZN(n8527) );
  AOI21_X1 U9436 ( .B1(n8529), .B2(n8528), .A(n8527), .ZN(n8532) );
  NOR2_X1 U9437 ( .A1(n10135), .A2(n8661), .ZN(n8531) );
  NAND2_X1 U9438 ( .A1(n10135), .A2(n8661), .ZN(n11426) );
  OAI21_X1 U9439 ( .B1(n8532), .B2(n8531), .A(n11426), .ZN(n8538) );
  NOR2_X1 U9440 ( .A1(n10358), .A2(n8524), .ZN(n8536) );
  NAND2_X1 U9441 ( .A1(data_addr_o_5_), .A2(n8694), .ZN(n8535) );
  NAND2_X1 U9442 ( .A1(n10358), .A2(n8524), .ZN(n11419) );
  OAI21_X1 U9443 ( .B1(n8536), .B2(n8535), .A(n11419), .ZN(n8537) );
  AOI21_X1 U9444 ( .B1(n8539), .B2(n8538), .A(n8537), .ZN(n8554) );
  NOR2_X1 U9445 ( .A1(n9805), .A2(n8672), .ZN(n8547) );
  NOR2_X1 U9446 ( .A1(n7816), .A2(n8665), .ZN(n8542) );
  NOR2_X1 U9447 ( .A1(n8547), .A2(n8542), .ZN(n8546) );
  NOR2_X1 U9448 ( .A1(n8237), .A2(n8673), .ZN(n8545) );
  NOR2_X1 U9449 ( .A1(data_addr_o_10_), .A2(n8670), .ZN(n8548) );
  NOR2_X1 U9450 ( .A1(n8545), .A2(n8548), .ZN(n8551) );
  NAND2_X1 U9451 ( .A1(n8546), .A2(n8551), .ZN(n8553) );
  NAND2_X1 U9452 ( .A1(n7816), .A2(n8665), .ZN(n11418) );
  NAND2_X1 U9453 ( .A1(n9805), .A2(n8672), .ZN(n11408) );
  OAI21_X1 U9454 ( .B1(n8547), .B2(n11418), .A(n11408), .ZN(n8550) );
  NAND2_X1 U9455 ( .A1(data_addr_o_9_), .A2(n8673), .ZN(n11412) );
  NAND2_X1 U9456 ( .A1(data_addr_o_10_), .A2(n8670), .ZN(n11413) );
  OAI21_X1 U9457 ( .B1(n8548), .B2(n11412), .A(n11413), .ZN(n8549) );
  AOI21_X1 U9458 ( .B1(n8551), .B2(n8550), .A(n8549), .ZN(n8552) );
  OAI21_X1 U9459 ( .B1(n8554), .B2(n8553), .A(n8552), .ZN(n8572) );
  NAND2_X1 U9460 ( .A1(data_addr_o_11_), .A2(n8671), .ZN(n11436) );
  NAND2_X1 U9461 ( .A1(n10499), .A2(n8677), .ZN(n11437) );
  OAI21_X1 U9462 ( .B1(n8555), .B2(n11436), .A(n11437), .ZN(n8559) );
  NAND2_X1 U9463 ( .A1(n10847), .A2(n8676), .ZN(n8556) );
  NAND2_X1 U9464 ( .A1(n10848), .A2(n8679), .ZN(n11451) );
  OAI21_X1 U9465 ( .B1(n8557), .B2(n8556), .A(n11451), .ZN(n8558) );
  AOI21_X1 U9466 ( .B1(n8560), .B2(n8559), .A(n8558), .ZN(n8569) );
  NAND2_X1 U9467 ( .A1(n10657), .A2(n8678), .ZN(n11444) );
  NAND2_X1 U9468 ( .A1(data_addr_o_16_), .A2(n11409), .ZN(n11443) );
  OAI21_X1 U9469 ( .B1(n8561), .B2(n11444), .A(n11443), .ZN(n8567) );
  NAND2_X1 U9470 ( .A1(n6813), .A2(n8691), .ZN(n8563) );
  NAND2_X1 U9471 ( .A1(n10857), .A2(n1417), .ZN(n8562) );
  OAI21_X1 U9472 ( .B1(n8564), .B2(n8563), .A(n8562), .ZN(n8565) );
  AOI21_X1 U9473 ( .B1(n8567), .B2(n8566), .A(n8565), .ZN(n8568) );
  OAI21_X1 U9474 ( .B1(n8570), .B2(n8569), .A(n8568), .ZN(n8571) );
  AOI21_X1 U9475 ( .B1(n8573), .B2(n8572), .A(n8571), .ZN(n8630) );
  NOR2_X1 U9476 ( .A1(n10898), .A2(n1539), .ZN(n8574) );
  NOR2_X1 U9477 ( .A1(n10738), .A2(n1485), .ZN(n8601) );
  NOR2_X1 U9478 ( .A1(n8574), .A2(n8601), .ZN(n8576) );
  NOR2_X1 U9479 ( .A1(n9923), .A2(n1542), .ZN(n8575) );
  NOR2_X1 U9480 ( .A1(n10606), .A2(n1480), .ZN(n8604) );
  NOR2_X1 U9481 ( .A1(n8575), .A2(n8604), .ZN(n8607) );
  NAND2_X1 U9482 ( .A1(n8576), .A2(n8607), .ZN(n8609) );
  NOR2_X1 U9483 ( .A1(n10202), .A2(n1516), .ZN(n8577) );
  NOR2_X1 U9484 ( .A1(n9915), .A2(n1489), .ZN(n8595) );
  NOR2_X1 U9485 ( .A1(n8577), .A2(n8595), .ZN(n8598) );
  NOR2_X1 U9486 ( .A1(n9846), .A2(n1512), .ZN(n8578) );
  NOR2_X1 U9487 ( .A1(n10530), .A2(n1492), .ZN(n8592) );
  NOR2_X1 U9488 ( .A1(n8578), .A2(n8592), .ZN(n8579) );
  NAND2_X1 U9489 ( .A1(n8598), .A2(n8579), .ZN(n8580) );
  NOR2_X1 U9490 ( .A1(n8609), .A2(n8580), .ZN(n8589) );
  NOR2_X1 U9491 ( .A1(n9886), .A2(n1523), .ZN(n8581) );
  NOR2_X1 U9492 ( .A1(n10914), .A2(n1501), .ZN(n8613) );
  NOR2_X1 U9493 ( .A1(n8581), .A2(n8613), .ZN(n8583) );
  NOR2_X1 U9494 ( .A1(n9955), .A2(n1526), .ZN(n8582) );
  NOR2_X1 U9495 ( .A1(data_addr_o_30_), .A2(n1496), .ZN(n8616) );
  NOR2_X1 U9496 ( .A1(n8582), .A2(n8616), .ZN(n8619) );
  NAND2_X1 U9497 ( .A1(n8583), .A2(n8619), .ZN(n8588) );
  NOR2_X1 U9498 ( .A1(n10662), .A2(n8693), .ZN(n8585) );
  NOR2_X1 U9499 ( .A1(n8585), .A2(pmp_addr_i[382]), .ZN(n8587) );
  INV_X1 U9500 ( .A(pmp_addr_i[383]), .ZN(n8586) );
  NAND2_X1 U9501 ( .A1(n8587), .A2(n8586), .ZN(n8623) );
  NOR2_X1 U9502 ( .A1(n8588), .A2(n8623), .ZN(n8626) );
  NAND2_X1 U9503 ( .A1(n8589), .A2(n8626), .ZN(n8629) );
  NAND2_X1 U9504 ( .A1(n9846), .A2(n1512), .ZN(n8591) );
  NAND2_X1 U9505 ( .A1(n10530), .A2(n1492), .ZN(n8590) );
  OAI21_X1 U9506 ( .B1(n8592), .B2(n8591), .A(n8590), .ZN(n8597) );
  NAND2_X1 U9507 ( .A1(n10202), .A2(n1516), .ZN(n8594) );
  NAND2_X1 U9508 ( .A1(n9915), .A2(n1489), .ZN(n8593) );
  OAI21_X1 U9509 ( .B1(n8595), .B2(n8594), .A(n8593), .ZN(n8596) );
  AOI21_X1 U9510 ( .B1(n8598), .B2(n8597), .A(n8596), .ZN(n8610) );
  NAND2_X1 U9511 ( .A1(n10898), .A2(n1539), .ZN(n8600) );
  NAND2_X1 U9512 ( .A1(n10738), .A2(n1485), .ZN(n8599) );
  OAI21_X1 U9513 ( .B1(n8601), .B2(n8600), .A(n8599), .ZN(n8606) );
  NAND2_X1 U9514 ( .A1(n9923), .A2(n1542), .ZN(n8603) );
  NAND2_X1 U9515 ( .A1(n10606), .A2(n1480), .ZN(n8602) );
  OAI21_X1 U9516 ( .B1(n8604), .B2(n8603), .A(n8602), .ZN(n8605) );
  AOI21_X1 U9517 ( .B1(n8607), .B2(n8606), .A(n8605), .ZN(n8608) );
  OAI21_X1 U9518 ( .B1(n8610), .B2(n8609), .A(n8608), .ZN(n8627) );
  NAND2_X1 U9519 ( .A1(n9886), .A2(n1523), .ZN(n8612) );
  NAND2_X1 U9520 ( .A1(n10914), .A2(n1501), .ZN(n8611) );
  OAI21_X1 U9521 ( .B1(n8613), .B2(n8612), .A(n8611), .ZN(n8618) );
  NAND2_X1 U9522 ( .A1(n9955), .A2(n1526), .ZN(n8615) );
  NAND2_X1 U9523 ( .A1(n10919), .A2(n1496), .ZN(n8614) );
  OAI21_X1 U9524 ( .B1(n8616), .B2(n8615), .A(n8614), .ZN(n8617) );
  AOI21_X1 U9525 ( .B1(n8619), .B2(n8618), .A(n8617), .ZN(n8624) );
  NAND2_X1 U9526 ( .A1(n10662), .A2(n8693), .ZN(n8620) );
  NOR2_X1 U9527 ( .A1(n8620), .A2(pmp_addr_i[382]), .ZN(n8621) );
  NAND2_X1 U9528 ( .A1(n8621), .A2(n8586), .ZN(n8622) );
  OAI21_X1 U9529 ( .B1(n8624), .B2(n8623), .A(n8622), .ZN(n8625) );
  AOI21_X1 U9530 ( .B1(n8627), .B2(n8626), .A(n8625), .ZN(n8628) );
  OAI21_X1 U9531 ( .B1(n8630), .B2(n8629), .A(n8628), .ZN(n8631) );
  NAND3_X1 U9532 ( .A1(n8632), .A2(n1644), .A3(n8631), .ZN(n8709) );
  XNOR2_X1 U9533 ( .A(n10627), .B(n8633), .ZN(n8640) );
  XNOR2_X1 U9534 ( .A(n10638), .B(n8634), .ZN(n8639) );
  XNOR2_X1 U9535 ( .A(n10629), .B(n8635), .ZN(n8638) );
  XNOR2_X1 U9536 ( .A(n10606), .B(n8636), .ZN(n8637) );
  NAND4_X1 U9537 ( .A1(n8640), .A2(n8639), .A3(n8638), .A4(n8637), .ZN(n8650)
         );
  XNOR2_X1 U9538 ( .A(n11285), .B(n8641), .ZN(n8648) );
  XNOR2_X1 U9539 ( .A(n10612), .B(n8642), .ZN(n8647) );
  XNOR2_X1 U9540 ( .A(data_addr_o_23_), .B(n8643), .ZN(n8646) );
  XNOR2_X1 U9541 ( .A(n10616), .B(n8644), .ZN(n8645) );
  NAND4_X1 U9542 ( .A1(n8648), .A2(n8647), .A3(n8646), .A4(n8645), .ZN(n8649)
         );
  NOR2_X1 U9543 ( .A1(n8650), .A2(n8649), .ZN(n8689) );
  XNOR2_X1 U9544 ( .A(data_addr_o_30_), .B(n8651), .ZN(n8658) );
  XNOR2_X1 U9545 ( .A(n10967), .B(n8652), .ZN(n8657) );
  XNOR2_X1 U9546 ( .A(n10614), .B(n8653), .ZN(n8656) );
  XNOR2_X1 U9547 ( .A(n10635), .B(n8654), .ZN(n8655) );
  NAND4_X1 U9548 ( .A1(n8658), .A2(n8657), .A3(n8656), .A4(n8655), .ZN(n8687)
         );
  XNOR2_X1 U9549 ( .A(n9955), .B(n8659), .ZN(n8685) );
  OAI22_X1 U9550 ( .A1(n11288), .A2(n8661), .B1(n22), .B2(n8526), .ZN(n8662)
         );
  INV_X1 U9551 ( .A(n8662), .ZN(n8664) );
  AOI21_X1 U9552 ( .B1(n8695), .B2(n8696), .A(n220), .ZN(n8663) );
  OAI211_X1 U9553 ( .C1(n7816), .C2(n8665), .A(n8664), .B(n8663), .ZN(n8666)
         );
  NOR2_X1 U9554 ( .A1(n8667), .A2(n8666), .ZN(n8668) );
  OAI21_X1 U9555 ( .B1(n6813), .B2(n8691), .A(n8668), .ZN(n8669) );
  INV_X1 U9556 ( .A(n8669), .ZN(n8684) );
  OAI22_X1 U9557 ( .A1(n8671), .A2(data_addr_o_11_), .B1(n11343), .B2(n8670), 
        .ZN(n8675) );
  OAI22_X1 U9558 ( .A1(data_addr_o_9_), .A2(n8673), .B1(n10281), .B2(n8672), 
        .ZN(n8674) );
  NOR2_X1 U9559 ( .A1(n8675), .A2(n8674), .ZN(n8683) );
  OAI22_X1 U9560 ( .A1(n8677), .A2(n31), .B1(data_addr_o_13_), .B2(n8676), 
        .ZN(n8681) );
  OAI22_X1 U9561 ( .A1(n8679), .A2(n9066), .B1(n10657), .B2(n8678), .ZN(n8680)
         );
  NOR2_X1 U9562 ( .A1(n8681), .A2(n8680), .ZN(n8682) );
  NAND4_X1 U9563 ( .A1(n8685), .A2(n8684), .A3(n8683), .A4(n8682), .ZN(n8686)
         );
  NOR2_X1 U9564 ( .A1(n8687), .A2(n8686), .ZN(n8688) );
  AND2_X1 U9565 ( .A1(n8689), .A2(n8688), .ZN(n11458) );
  XNOR2_X1 U9566 ( .A(n11014), .B(n8690), .ZN(n8705) );
  AND2_X1 U9567 ( .A1(data_addr_o_17_), .A2(n8691), .ZN(n11449) );
  OAI21_X1 U9568 ( .B1(n11006), .B2(n8692), .A(n11451), .ZN(n11454) );
  NOR2_X1 U9569 ( .A1(n11449), .A2(n11454), .ZN(n8704) );
  XNOR2_X1 U9570 ( .A(n12123), .B(n8693), .ZN(n8702) );
  AND2_X1 U9571 ( .A1(n11418), .A2(n11419), .ZN(n8699) );
  AND2_X1 U9572 ( .A1(n10486), .A2(n8694), .ZN(n11417) );
  NAND2_X1 U9573 ( .A1(data_addr_o_3_), .A2(n8526), .ZN(n11429) );
  OAI211_X1 U9574 ( .C1(n8696), .C2(n8695), .A(n11426), .B(n11429), .ZN(n8697)
         );
  NOR2_X1 U9575 ( .A1(n11417), .A2(n8697), .ZN(n8698) );
  NAND4_X1 U9576 ( .A1(n8699), .A2(n11437), .A3(n11444), .A4(n8698), .ZN(n8701) );
  NAND4_X1 U9577 ( .A1(n11413), .A2(n11412), .A3(n11436), .A4(n11408), .ZN(
        n8700) );
  NOR3_X1 U9578 ( .A1(n8702), .A2(n8701), .A3(n8700), .ZN(n8703) );
  NAND4_X1 U9579 ( .A1(n11458), .A2(n8705), .A3(n8704), .A4(n8703), .ZN(n8708)
         );
  MUX2_X1 U9580 ( .A(pmp_cfg_i[96]), .B(pmp_cfg_i[97]), .S(n11019), .Z(n8707)
         );
  NAND2_X1 U9581 ( .A1(n8706), .A2(n8707), .ZN(n11427) );
  AOI21_X1 U9582 ( .B1(n8709), .B2(n8708), .A(n11427), .ZN(n8710) );
  NOR2_X1 U9583 ( .A1(n8711), .A2(n8710), .ZN(n9338) );
  NOR2_X1 U9584 ( .A1(n10047), .A2(pmp_addr_i[270]), .ZN(n8712) );
  INV_X1 U9585 ( .A(data_addr_i[17]), .ZN(n8757) );
  NOR2_X1 U9586 ( .A1(n8757), .A2(pmp_addr_i[271]), .ZN(n8760) );
  NOR2_X1 U9587 ( .A1(n8712), .A2(n8760), .ZN(n8763) );
  NOR2_X1 U9588 ( .A1(pmp_addr_i[268]), .A2(n10000), .ZN(n8713) );
  NOR2_X1 U9589 ( .A1(pmp_addr_i[269]), .A2(n10721), .ZN(n8756) );
  NOR2_X1 U9590 ( .A1(n8713), .A2(n8756), .ZN(n8714) );
  NAND2_X1 U9591 ( .A1(n8763), .A2(n8714), .ZN(n8766) );
  NOR2_X1 U9592 ( .A1(pmp_addr_i[264]), .A2(n10701), .ZN(n8715) );
  NOR2_X1 U9593 ( .A1(pmp_addr_i[265]), .A2(n10711), .ZN(n8747) );
  NOR2_X1 U9594 ( .A1(n8715), .A2(n8747), .ZN(n8717) );
  NOR2_X1 U9595 ( .A1(pmp_addr_i[266]), .A2(n10005), .ZN(n8716) );
  NOR2_X1 U9596 ( .A1(pmp_addr_i[267]), .A2(n11006), .ZN(n8750) );
  NOR2_X1 U9597 ( .A1(n8716), .A2(n8750), .ZN(n8753) );
  NAND2_X1 U9598 ( .A1(n8717), .A2(n8753), .ZN(n8718) );
  NOR2_X1 U9599 ( .A1(n8766), .A2(n8718), .ZN(n8769) );
  NOR2_X1 U9600 ( .A1(pmp_addr_i[258]), .A2(n6123), .ZN(n8719) );
  NOR2_X1 U9601 ( .A1(pmp_addr_i[259]), .A2(n10346), .ZN(n8725) );
  NOR2_X1 U9602 ( .A1(n8719), .A2(n8725), .ZN(n8728) );
  NOR2_X1 U9603 ( .A1(pmp_addr_i[257]), .A2(n9350), .ZN(n8722) );
  NAND2_X1 U9604 ( .A1(pmp_addr_i[256]), .A2(n10651), .ZN(n8721) );
  NAND2_X1 U9605 ( .A1(pmp_addr_i[257]), .A2(n9350), .ZN(n8720) );
  OAI21_X1 U9606 ( .B1(n8722), .B2(n8721), .A(n8720), .ZN(n8727) );
  NAND2_X1 U9607 ( .A1(pmp_addr_i[258]), .A2(n8406), .ZN(n8724) );
  NAND2_X1 U9608 ( .A1(pmp_addr_i[259]), .A2(n10346), .ZN(n8723) );
  OAI21_X1 U9609 ( .B1(n8725), .B2(n8724), .A(n8723), .ZN(n8726) );
  AOI21_X1 U9610 ( .B1(n8728), .B2(n8727), .A(n8726), .ZN(n8744) );
  NOR2_X1 U9611 ( .A1(pmp_addr_i[260]), .A2(n9363), .ZN(n8729) );
  NOR2_X1 U9612 ( .A1(pmp_addr_i[261]), .A2(n10697), .ZN(n8734) );
  NOR2_X1 U9613 ( .A1(n8729), .A2(n8734), .ZN(n8731) );
  INV_X1 U9614 ( .A(data_addr_i[8]), .ZN(n8735) );
  NOR2_X1 U9615 ( .A1(pmp_addr_i[262]), .A2(n8735), .ZN(n8730) );
  NOR2_X1 U9616 ( .A1(pmp_addr_i[263]), .A2(n6140), .ZN(n8738) );
  NOR2_X1 U9617 ( .A1(n8730), .A2(n8738), .ZN(n8741) );
  NAND2_X1 U9618 ( .A1(n8731), .A2(n8741), .ZN(n8743) );
  NAND2_X1 U9619 ( .A1(pmp_addr_i[260]), .A2(n10362), .ZN(n8733) );
  NAND2_X1 U9620 ( .A1(pmp_addr_i[261]), .A2(n6400), .ZN(n8732) );
  OAI21_X1 U9621 ( .B1(n8734), .B2(n8733), .A(n8732), .ZN(n8740) );
  NAND2_X1 U9622 ( .A1(pmp_addr_i[262]), .A2(n8735), .ZN(n8737) );
  NAND2_X1 U9623 ( .A1(pmp_addr_i[263]), .A2(n6140), .ZN(n8736) );
  OAI21_X1 U9624 ( .B1(n8738), .B2(n8737), .A(n8736), .ZN(n8739) );
  AOI21_X1 U9625 ( .B1(n8741), .B2(n8740), .A(n8739), .ZN(n8742) );
  OAI21_X1 U9626 ( .B1(n8744), .B2(n8743), .A(n8742), .ZN(n8768) );
  NAND2_X1 U9627 ( .A1(pmp_addr_i[264]), .A2(n6141), .ZN(n8746) );
  NAND2_X1 U9628 ( .A1(pmp_addr_i[265]), .A2(n9508), .ZN(n8745) );
  OAI21_X1 U9629 ( .B1(n8747), .B2(n8746), .A(n8745), .ZN(n8752) );
  NAND2_X1 U9630 ( .A1(pmp_addr_i[266]), .A2(n10005), .ZN(n8749) );
  NAND2_X1 U9631 ( .A1(pmp_addr_i[267]), .A2(n11006), .ZN(n8748) );
  OAI21_X1 U9632 ( .B1(n8750), .B2(n8749), .A(n8748), .ZN(n8751) );
  AOI21_X1 U9633 ( .B1(n8753), .B2(n8752), .A(n8751), .ZN(n8765) );
  NAND2_X1 U9634 ( .A1(pmp_addr_i[268]), .A2(n10000), .ZN(n8755) );
  NAND2_X1 U9635 ( .A1(pmp_addr_i[269]), .A2(n10338), .ZN(n8754) );
  OAI21_X1 U9636 ( .B1(n8756), .B2(n8755), .A(n8754), .ZN(n8762) );
  NAND2_X1 U9637 ( .A1(n10047), .A2(pmp_addr_i[270]), .ZN(n8759) );
  NAND2_X1 U9638 ( .A1(n8757), .A2(pmp_addr_i[271]), .ZN(n8758) );
  OAI21_X1 U9639 ( .B1(n8760), .B2(n8759), .A(n8758), .ZN(n8761) );
  AOI21_X1 U9640 ( .B1(n8763), .B2(n8762), .A(n8761), .ZN(n8764) );
  OAI21_X1 U9641 ( .B1(n8766), .B2(n8765), .A(n8764), .ZN(n8767) );
  AOI21_X1 U9642 ( .B1(n8769), .B2(n8768), .A(n8767), .ZN(n8829) );
  NOR2_X1 U9643 ( .A1(n9425), .A2(pmp_addr_i[276]), .ZN(n8770) );
  NOR2_X1 U9644 ( .A1(n10764), .A2(pmp_addr_i[277]), .ZN(n8794) );
  NOR2_X1 U9645 ( .A1(n8770), .A2(n8794), .ZN(n8772) );
  NOR2_X1 U9646 ( .A1(n10428), .A2(pmp_addr_i[278]), .ZN(n8771) );
  NOR2_X1 U9647 ( .A1(n10429), .A2(pmp_addr_i[279]), .ZN(n8797) );
  NOR2_X1 U9648 ( .A1(n8771), .A2(n8797), .ZN(n8800) );
  NAND2_X1 U9649 ( .A1(n8772), .A2(n8800), .ZN(n8802) );
  NOR2_X1 U9650 ( .A1(n6192), .A2(pmp_addr_i[275]), .ZN(n8788) );
  NOR2_X1 U9651 ( .A1(n6188), .A2(pmp_addr_i[274]), .ZN(n8773) );
  NOR2_X1 U9652 ( .A1(n8788), .A2(n8773), .ZN(n8791) );
  NOR2_X1 U9653 ( .A1(n10414), .A2(pmp_addr_i[273]), .ZN(n8785) );
  NOR2_X1 U9654 ( .A1(n10060), .A2(pmp_addr_i[272]), .ZN(n8774) );
  NOR2_X1 U9655 ( .A1(n8785), .A2(n8774), .ZN(n8775) );
  NAND2_X1 U9656 ( .A1(n8791), .A2(n8775), .ZN(n8776) );
  NOR2_X1 U9657 ( .A1(n8802), .A2(n8776), .ZN(n8782) );
  NOR2_X1 U9658 ( .A1(n10439), .A2(pmp_addr_i[280]), .ZN(n8777) );
  NOR2_X1 U9659 ( .A1(n9438), .A2(pmp_addr_i[281]), .ZN(n8806) );
  NOR2_X1 U9660 ( .A1(n8777), .A2(n8806), .ZN(n8779) );
  INV_X1 U9661 ( .A(data_addr_i[28]), .ZN(n8807) );
  NOR2_X1 U9662 ( .A1(n8807), .A2(pmp_addr_i[282]), .ZN(n8778) );
  NOR2_X1 U9663 ( .A1(n6216), .A2(pmp_addr_i[283]), .ZN(n8810) );
  NOR2_X1 U9664 ( .A1(n8778), .A2(n8810), .ZN(n8813) );
  NAND2_X1 U9665 ( .A1(n8779), .A2(n8813), .ZN(n8781) );
  INV_X1 U9666 ( .A(data_addr_i[30]), .ZN(n8814) );
  NOR2_X1 U9667 ( .A1(n8814), .A2(pmp_addr_i[284]), .ZN(n8780) );
  NOR2_X1 U9668 ( .A1(n10107), .A2(pmp_addr_i[285]), .ZN(n8817) );
  OR2_X1 U9669 ( .A1(n8780), .A2(n8817), .ZN(n8822) );
  NOR2_X1 U9670 ( .A1(n8781), .A2(n8822), .ZN(n8825) );
  NAND2_X1 U9671 ( .A1(n8782), .A2(n8825), .ZN(n8828) );
  NAND2_X1 U9672 ( .A1(n10403), .A2(pmp_addr_i[272]), .ZN(n8784) );
  NAND2_X1 U9673 ( .A1(n10414), .A2(pmp_addr_i[273]), .ZN(n8783) );
  OAI21_X1 U9674 ( .B1(n8785), .B2(n8784), .A(n8783), .ZN(n8790) );
  NAND2_X1 U9675 ( .A1(n6188), .A2(pmp_addr_i[274]), .ZN(n8787) );
  NAND2_X1 U9676 ( .A1(n9418), .A2(pmp_addr_i[275]), .ZN(n8786) );
  OAI21_X1 U9677 ( .B1(n8788), .B2(n8787), .A(n8786), .ZN(n8789) );
  AOI21_X1 U9678 ( .B1(n8791), .B2(n8790), .A(n8789), .ZN(n8803) );
  NAND2_X1 U9679 ( .A1(n9425), .A2(pmp_addr_i[276]), .ZN(n8793) );
  NAND2_X1 U9680 ( .A1(n10764), .A2(pmp_addr_i[277]), .ZN(n8792) );
  OAI21_X1 U9681 ( .B1(n8794), .B2(n8793), .A(n8792), .ZN(n8799) );
  NAND2_X1 U9682 ( .A1(n10428), .A2(pmp_addr_i[278]), .ZN(n8796) );
  NAND2_X1 U9683 ( .A1(n10429), .A2(pmp_addr_i[279]), .ZN(n8795) );
  OAI21_X1 U9684 ( .B1(n8797), .B2(n8796), .A(n8795), .ZN(n8798) );
  AOI21_X1 U9685 ( .B1(n8800), .B2(n8799), .A(n8798), .ZN(n8801) );
  OAI21_X1 U9686 ( .B1(n8803), .B2(n8802), .A(n8801), .ZN(n8826) );
  NAND2_X1 U9687 ( .A1(n6202), .A2(pmp_addr_i[280]), .ZN(n8805) );
  NAND2_X1 U9688 ( .A1(n6212), .A2(pmp_addr_i[281]), .ZN(n8804) );
  OAI21_X1 U9689 ( .B1(n8806), .B2(n8805), .A(n8804), .ZN(n8812) );
  NAND2_X1 U9690 ( .A1(n8807), .A2(pmp_addr_i[282]), .ZN(n8809) );
  NAND2_X1 U9691 ( .A1(n10782), .A2(pmp_addr_i[283]), .ZN(n8808) );
  OAI21_X1 U9692 ( .B1(n8810), .B2(n8809), .A(n8808), .ZN(n8811) );
  AOI21_X1 U9693 ( .B1(n8813), .B2(n8812), .A(n8811), .ZN(n8823) );
  NAND2_X1 U9694 ( .A1(n8814), .A2(pmp_addr_i[284]), .ZN(n8816) );
  NAND2_X1 U9695 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[285]), .ZN(n8815)
         );
  OAI21_X1 U9696 ( .B1(n8817), .B2(n8816), .A(n8815), .ZN(n8820) );
  INV_X1 U9697 ( .A(n8818), .ZN(n8819) );
  NOR2_X1 U9698 ( .A1(n8820), .A2(n8819), .ZN(n8821) );
  OAI21_X1 U9699 ( .B1(n8823), .B2(n8822), .A(n8821), .ZN(n8824) );
  AOI21_X1 U9700 ( .B1(n8826), .B2(n8825), .A(n8824), .ZN(n8827) );
  OAI21_X1 U9701 ( .B1(n8829), .B2(n8828), .A(n8827), .ZN(n8949) );
  NOR2_X1 U9702 ( .A1(n9987), .A2(n11609), .ZN(n8878) );
  NOR2_X1 U9703 ( .A1(n11309), .A2(n9008), .ZN(n8831) );
  NOR2_X1 U9704 ( .A1(n8878), .A2(n8831), .ZN(n8833) );
  NOR2_X1 U9705 ( .A1(n10857), .A2(n1722), .ZN(n8881) );
  NAND2_X1 U9706 ( .A1(n8757), .A2(n8879), .ZN(n8991) );
  INV_X1 U9707 ( .A(n8991), .ZN(n8832) );
  NOR2_X1 U9708 ( .A1(n8881), .A2(n8832), .ZN(n8884) );
  NAND2_X1 U9709 ( .A1(n8833), .A2(n8884), .ZN(n8887) );
  NOR2_X1 U9710 ( .A1(n10508), .A2(n8979), .ZN(n8836) );
  NOR2_X1 U9711 ( .A1(n31), .A2(n8987), .ZN(n8871) );
  NOR2_X1 U9712 ( .A1(n8836), .A2(n8871), .ZN(n8840) );
  NOR2_X1 U9713 ( .A1(n10847), .A2(n8986), .ZN(n8839) );
  NOR2_X1 U9714 ( .A1(n10848), .A2(n8988), .ZN(n8872) );
  NOR2_X1 U9715 ( .A1(n8839), .A2(n8872), .ZN(n8875) );
  NAND2_X1 U9716 ( .A1(n8840), .A2(n8875), .ZN(n8841) );
  NOR2_X1 U9717 ( .A1(n8887), .A2(n8841), .ZN(n8890) );
  NOR2_X1 U9718 ( .A1(n10486), .A2(n8968), .ZN(n8843) );
  NOR2_X1 U9719 ( .A1(n11331), .A2(n8977), .ZN(n8852) );
  NOR2_X1 U9720 ( .A1(n8843), .A2(n8852), .ZN(n8855) );
  INV_X1 U9721 ( .A(n8972), .ZN(n8844) );
  OR2_X1 U9722 ( .A1(n10129), .A2(n8844), .ZN(n8848) );
  INV_X1 U9723 ( .A(n8971), .ZN(n8845) );
  OR2_X1 U9724 ( .A1(n22), .A2(n8845), .ZN(n8847) );
  AND2_X1 U9725 ( .A1(n22), .A2(n8845), .ZN(n8846) );
  AOI21_X1 U9726 ( .B1(n8848), .B2(n8847), .A(n8846), .ZN(n8850) );
  NOR2_X1 U9727 ( .A1(n10479), .A2(n5786), .ZN(n8849) );
  NAND2_X1 U9728 ( .A1(n10479), .A2(n5786), .ZN(n11624) );
  OAI21_X1 U9729 ( .B1(n8850), .B2(n8849), .A(n11624), .ZN(n8854) );
  NAND2_X1 U9730 ( .A1(n10486), .A2(n8968), .ZN(n8851) );
  NAND2_X1 U9731 ( .A1(n11331), .A2(n8977), .ZN(n11601) );
  OAI21_X1 U9732 ( .B1(n8852), .B2(n8851), .A(n11601), .ZN(n8853) );
  AOI21_X1 U9733 ( .B1(n8855), .B2(n8854), .A(n8853), .ZN(n8870) );
  NOR2_X1 U9734 ( .A1(n10494), .A2(n8980), .ZN(n8863) );
  NOR2_X1 U9735 ( .A1(n10493), .A2(n8969), .ZN(n8858) );
  NOR2_X1 U9736 ( .A1(n8863), .A2(n8858), .ZN(n8862) );
  NOR2_X1 U9737 ( .A1(n10504), .A2(n8981), .ZN(n8861) );
  NOR2_X1 U9738 ( .A1(n10838), .A2(n8978), .ZN(n8864) );
  NOR2_X1 U9739 ( .A1(n8861), .A2(n8864), .ZN(n8867) );
  NAND2_X1 U9740 ( .A1(n8862), .A2(n8867), .ZN(n8869) );
  NAND2_X1 U9741 ( .A1(n10493), .A2(n8969), .ZN(n11631) );
  NAND2_X1 U9742 ( .A1(n10494), .A2(n8980), .ZN(n11634) );
  OAI21_X1 U9743 ( .B1(n8863), .B2(n11631), .A(n11634), .ZN(n8866) );
  NAND2_X1 U9744 ( .A1(n10504), .A2(n8981), .ZN(n11615) );
  NAND2_X1 U9745 ( .A1(n10838), .A2(n8978), .ZN(n11614) );
  OAI21_X1 U9746 ( .B1(n8864), .B2(n11615), .A(n11614), .ZN(n8865) );
  AOI21_X1 U9747 ( .B1(n8867), .B2(n8866), .A(n8865), .ZN(n8868) );
  OAI21_X1 U9748 ( .B1(n8870), .B2(n8869), .A(n8868), .ZN(n8889) );
  NAND2_X1 U9749 ( .A1(n10508), .A2(n8979), .ZN(n11590) );
  NAND2_X1 U9750 ( .A1(n31), .A2(n8987), .ZN(n11584) );
  OAI21_X1 U9751 ( .B1(n8871), .B2(n11590), .A(n11584), .ZN(n8874) );
  NAND2_X1 U9752 ( .A1(n10847), .A2(n8986), .ZN(n11594) );
  NAND2_X1 U9753 ( .A1(n10848), .A2(n8988), .ZN(n11589) );
  OAI21_X1 U9754 ( .B1(n8872), .B2(n11594), .A(n11589), .ZN(n8873) );
  AOI21_X1 U9755 ( .B1(n8875), .B2(n8874), .A(n8873), .ZN(n8886) );
  NAND2_X1 U9756 ( .A1(n11309), .A2(n9008), .ZN(n8877) );
  NAND2_X1 U9757 ( .A1(n10335), .A2(n11609), .ZN(n8876) );
  OAI21_X1 U9758 ( .B1(n8878), .B2(n8877), .A(n8876), .ZN(n8883) );
  NAND2_X1 U9759 ( .A1(data_addr_o_17_), .A2(n1776), .ZN(n11627) );
  NAND2_X1 U9760 ( .A1(n10857), .A2(n1722), .ZN(n8880) );
  OAI21_X1 U9761 ( .B1(n8881), .B2(n11627), .A(n8880), .ZN(n8882) );
  AOI21_X1 U9762 ( .B1(n8884), .B2(n8883), .A(n8882), .ZN(n8885) );
  OAI21_X1 U9763 ( .B1(n8887), .B2(n8886), .A(n8885), .ZN(n8888) );
  AOI21_X1 U9764 ( .B1(n8890), .B2(n8889), .A(n8888), .ZN(n8947) );
  NOR2_X1 U9765 ( .A1(n10898), .A2(n1695), .ZN(n8891) );
  NOR2_X1 U9766 ( .A1(n10738), .A2(n1664), .ZN(n8918) );
  NOR2_X1 U9767 ( .A1(n8891), .A2(n8918), .ZN(n8893) );
  NOR2_X1 U9768 ( .A1(n10903), .A2(n1698), .ZN(n8892) );
  NOR2_X1 U9769 ( .A1(n10267), .A2(n1660), .ZN(n8921) );
  NOR2_X1 U9770 ( .A1(n8892), .A2(n8921), .ZN(n8924) );
  NAND2_X1 U9771 ( .A1(n8893), .A2(n8924), .ZN(n8926) );
  INV_X1 U9772 ( .A(n8985), .ZN(n8909) );
  NOR2_X1 U9773 ( .A1(n11312), .A2(n8909), .ZN(n8894) );
  NOR2_X1 U9774 ( .A1(n9529), .A2(n1667), .ZN(n8912) );
  NOR2_X1 U9775 ( .A1(n8894), .A2(n8912), .ZN(n8915) );
  NOR2_X1 U9776 ( .A1(n9846), .A2(n1713), .ZN(n8895) );
  NOR2_X1 U9777 ( .A1(n10530), .A2(n1670), .ZN(n8908) );
  NOR2_X1 U9778 ( .A1(n8895), .A2(n8908), .ZN(n8896) );
  NAND2_X1 U9779 ( .A1(n8915), .A2(n8896), .ZN(n8897) );
  NOR2_X1 U9780 ( .A1(n8926), .A2(n8897), .ZN(n8905) );
  NOR2_X1 U9781 ( .A1(n9886), .A2(n1679), .ZN(n8898) );
  NOR2_X1 U9782 ( .A1(n10635), .A2(n1654), .ZN(n8930) );
  NOR2_X1 U9783 ( .A1(n8898), .A2(n8930), .ZN(n8900) );
  NOR2_X1 U9784 ( .A1(n10918), .A2(n1682), .ZN(n8899) );
  NOR2_X1 U9785 ( .A1(n10919), .A2(n1650), .ZN(n8933) );
  NOR2_X1 U9786 ( .A1(n8899), .A2(n8933), .ZN(n8936) );
  NAND2_X1 U9787 ( .A1(n8900), .A2(n8936), .ZN(n8904) );
  NOR2_X1 U9788 ( .A1(n10662), .A2(n1704), .ZN(n8901) );
  NOR2_X1 U9789 ( .A1(n8901), .A2(pmp_addr_i[254]), .ZN(n8903) );
  INV_X1 U9790 ( .A(pmp_addr_i[255]), .ZN(n8902) );
  NAND2_X1 U9791 ( .A1(n8903), .A2(n8902), .ZN(n8940) );
  NOR2_X1 U9792 ( .A1(n8904), .A2(n8940), .ZN(n8943) );
  NAND2_X1 U9793 ( .A1(n8905), .A2(n8943), .ZN(n8946) );
  NAND2_X1 U9794 ( .A1(n9846), .A2(n1713), .ZN(n8907) );
  NAND2_X1 U9795 ( .A1(n10530), .A2(n1670), .ZN(n8906) );
  OAI21_X1 U9796 ( .B1(n8908), .B2(n8907), .A(n8906), .ZN(n8914) );
  NAND2_X1 U9797 ( .A1(n10202), .A2(n8909), .ZN(n8911) );
  NAND2_X1 U9798 ( .A1(n9529), .A2(n1667), .ZN(n8910) );
  OAI21_X1 U9799 ( .B1(n8912), .B2(n8911), .A(n8910), .ZN(n8913) );
  AOI21_X1 U9800 ( .B1(n8915), .B2(n8914), .A(n8913), .ZN(n8927) );
  NAND2_X1 U9801 ( .A1(data_addr_o_23_), .A2(n1695), .ZN(n8917) );
  NAND2_X1 U9802 ( .A1(n10738), .A2(n1664), .ZN(n8916) );
  OAI21_X1 U9803 ( .B1(n8918), .B2(n8917), .A(n8916), .ZN(n8923) );
  NAND2_X1 U9804 ( .A1(n10903), .A2(n1698), .ZN(n8920) );
  NAND2_X1 U9805 ( .A1(n10267), .A2(n1660), .ZN(n8919) );
  OAI21_X1 U9806 ( .B1(n8921), .B2(n8920), .A(n8919), .ZN(n8922) );
  AOI21_X1 U9807 ( .B1(n8924), .B2(n8923), .A(n8922), .ZN(n8925) );
  OAI21_X1 U9808 ( .B1(n8927), .B2(n8926), .A(n8925), .ZN(n8944) );
  NAND2_X1 U9809 ( .A1(n9886), .A2(n1679), .ZN(n8929) );
  NAND2_X1 U9810 ( .A1(n10635), .A2(n1654), .ZN(n8928) );
  OAI21_X1 U9811 ( .B1(n8930), .B2(n8929), .A(n8928), .ZN(n8935) );
  NAND2_X1 U9812 ( .A1(n10918), .A2(n1682), .ZN(n8932) );
  NAND2_X1 U9813 ( .A1(n10919), .A2(n1650), .ZN(n8931) );
  OAI21_X1 U9814 ( .B1(n8933), .B2(n8932), .A(n8931), .ZN(n8934) );
  AOI21_X1 U9815 ( .B1(n8936), .B2(n8935), .A(n8934), .ZN(n8941) );
  NAND2_X1 U9816 ( .A1(n10662), .A2(n1704), .ZN(n8937) );
  NOR2_X1 U9817 ( .A1(n8937), .A2(pmp_addr_i[254]), .ZN(n8938) );
  NAND2_X1 U9818 ( .A1(n8938), .A2(n8902), .ZN(n8939) );
  OAI21_X1 U9819 ( .B1(n8941), .B2(n8940), .A(n8939), .ZN(n8942) );
  AOI21_X1 U9820 ( .B1(n8944), .B2(n8943), .A(n8942), .ZN(n8945) );
  OAI21_X1 U9821 ( .B1(n8947), .B2(n8946), .A(n8945), .ZN(n8948) );
  XNOR2_X1 U9822 ( .A(data_addr_o_26_), .B(n8950), .ZN(n8957) );
  XNOR2_X1 U9823 ( .A(n10635), .B(n8951), .ZN(n8956) );
  XNOR2_X1 U9824 ( .A(data_addr_o_30_), .B(n8952), .ZN(n8955) );
  XNOR2_X1 U9825 ( .A(n11283), .B(n8953), .ZN(n8954) );
  NAND4_X1 U9826 ( .A1(n8957), .A2(n8956), .A3(n8955), .A4(n8954), .ZN(n8967)
         );
  XNOR2_X1 U9827 ( .A(data_addr_o_23_), .B(n8958), .ZN(n8965) );
  XNOR2_X1 U9828 ( .A(n11313), .B(n8959), .ZN(n8964) );
  XNOR2_X1 U9829 ( .A(n11322), .B(n8960), .ZN(n8963) );
  XNOR2_X1 U9830 ( .A(n11298), .B(n8961), .ZN(n8962) );
  NAND4_X1 U9831 ( .A1(n8965), .A2(n8964), .A3(n8963), .A4(n8962), .ZN(n8966)
         );
  NOR2_X1 U9832 ( .A1(n8967), .A2(n8966), .ZN(n9006) );
  OAI22_X1 U9833 ( .A1(n8969), .A2(n7816), .B1(n11255), .B2(n8968), .ZN(n8970)
         );
  INV_X1 U9834 ( .A(n8970), .ZN(n8976) );
  OAI22_X1 U9835 ( .A1(n10130), .A2(n8845), .B1(n11259), .B2(n8844), .ZN(n8973) );
  AOI21_X1 U9836 ( .B1(n8974), .B2(n12058), .A(n8973), .ZN(n8975) );
  OAI211_X1 U9837 ( .C1(n8977), .C2(n10953), .A(n8976), .B(n8975), .ZN(n8984)
         );
  OAI22_X1 U9838 ( .A1(n8979), .A2(data_addr_o_11_), .B1(n11343), .B2(n8978), 
        .ZN(n8983) );
  OAI22_X1 U9839 ( .A1(n8237), .A2(n8981), .B1(n10836), .B2(n8980), .ZN(n8982)
         );
  NOR3_X1 U9840 ( .A1(n8984), .A2(n8983), .A3(n8982), .ZN(n8994) );
  XNOR2_X1 U9841 ( .A(n11312), .B(n8985), .ZN(n8993) );
  OAI22_X1 U9842 ( .A1(n8987), .A2(data_addr_o_12_), .B1(n6649), .B2(n8986), 
        .ZN(n8990) );
  OAI22_X1 U9843 ( .A1(n8988), .A2(data_addr_o_14_), .B1(n10657), .B2(n9008), 
        .ZN(n8989) );
  NOR2_X1 U9844 ( .A1(n8990), .A2(n8989), .ZN(n8992) );
  NAND4_X1 U9845 ( .A1(n8994), .A2(n8993), .A3(n8992), .A4(n8991), .ZN(n9000)
         );
  XNOR2_X1 U9846 ( .A(n10899), .B(n8995), .ZN(n8998) );
  XNOR2_X1 U9847 ( .A(n11320), .B(n8996), .ZN(n8997) );
  NAND2_X1 U9848 ( .A1(n8998), .A2(n8997), .ZN(n8999) );
  NOR2_X1 U9849 ( .A1(n9000), .A2(n8999), .ZN(n9005) );
  XNOR2_X1 U9850 ( .A(n11285), .B(n9001), .ZN(n9004) );
  XNOR2_X1 U9851 ( .A(n11303), .B(n9002), .ZN(n9003) );
  AND4_X1 U9852 ( .A1(n9006), .A2(n9005), .A3(n9004), .A4(n9003), .ZN(n11639)
         );
  XNOR2_X1 U9853 ( .A(n9007), .B(n12123), .ZN(n9018) );
  XNOR2_X1 U9854 ( .A(n9987), .B(n11607), .ZN(n9013) );
  AND2_X1 U9855 ( .A1(data_addr_o_15_), .A2(n9008), .ZN(n11582) );
  AOI21_X1 U9856 ( .B1(n11259), .B2(n8844), .A(n9009), .ZN(n9010) );
  NAND2_X1 U9857 ( .A1(n22), .A2(n8845), .ZN(n11598) );
  NAND4_X1 U9858 ( .A1(n11631), .A2(n9010), .A3(n11624), .A4(n11598), .ZN(
        n9011) );
  NOR2_X1 U9859 ( .A1(n11582), .A2(n9011), .ZN(n9012) );
  NAND4_X1 U9860 ( .A1(n9013), .A2(n9012), .A3(n11589), .A4(n11594), .ZN(n9016) );
  OAI211_X1 U9861 ( .C1(n11291), .C2(n9014), .A(n11615), .B(n11601), .ZN(
        n11621) );
  NAND4_X1 U9862 ( .A1(n11614), .A2(n11584), .A3(n11590), .A4(n11634), .ZN(
        n9015) );
  NOR3_X1 U9863 ( .A1(n9016), .A2(n11621), .A3(n9015), .ZN(n9017) );
  NAND4_X1 U9864 ( .A1(n11639), .A2(n9018), .A3(n9017), .A4(n11627), .ZN(n9019) );
  INV_X1 U9865 ( .A(pmp_cfg_i[64]), .ZN(n9022) );
  NAND2_X1 U9866 ( .A1(data_we_i), .A2(pmp_cfg_i[65]), .ZN(n9021) );
  OAI21_X1 U9867 ( .B1(n9022), .B2(n11019), .A(n9021), .ZN(n11596) );
  NAND2_X1 U9868 ( .A1(n9023), .A2(n11596), .ZN(n9337) );
  XNOR2_X1 U9869 ( .A(n10747), .B(n9276), .ZN(n9027) );
  XNOR2_X1 U9870 ( .A(data_addr_o_30_), .B(n9279), .ZN(n9026) );
  XNOR2_X1 U9871 ( .A(n11313), .B(n9268), .ZN(n9025) );
  XNOR2_X1 U9872 ( .A(n10629), .B(n9261), .ZN(n9024) );
  NAND4_X1 U9873 ( .A1(n9027), .A2(n9026), .A3(n9025), .A4(n9024), .ZN(n9033)
         );
  XNOR2_X1 U9874 ( .A(n11283), .B(n9270), .ZN(n9031) );
  XNOR2_X1 U9875 ( .A(n11320), .B(n9263), .ZN(n9030) );
  XNOR2_X1 U9876 ( .A(n10967), .B(n9199), .ZN(n9029) );
  XNOR2_X1 U9877 ( .A(data_addr_o_23_), .B(n9260), .ZN(n9028) );
  NAND4_X1 U9878 ( .A1(n9031), .A2(n9030), .A3(n9029), .A4(n9028), .ZN(n9032)
         );
  NOR2_X1 U9879 ( .A1(n9033), .A2(n9032), .ZN(n9056) );
  OAI22_X1 U9880 ( .A1(n9034), .A2(data_addr_o_5_), .B1(n10953), .B2(n9071), 
        .ZN(n9211) );
  INV_X1 U9881 ( .A(n9211), .ZN(n9039) );
  INV_X1 U9882 ( .A(n9213), .ZN(n9060) );
  OAI22_X1 U9883 ( .A1(n10135), .A2(n9059), .B1(n10130), .B2(n9060), .ZN(n9037) );
  INV_X1 U9884 ( .A(n9212), .ZN(n9035) );
  OAI21_X1 U9885 ( .B1(n10129), .B2(n9035), .A(pmp_cfg_i[84]), .ZN(n9036) );
  NOR2_X1 U9886 ( .A1(n9037), .A2(n9036), .ZN(n9038) );
  OAI211_X1 U9887 ( .C1(n9058), .C2(n7816), .A(n9039), .B(n9038), .ZN(n9042)
         );
  OAI22_X1 U9888 ( .A1(n9073), .A2(data_addr_o_11_), .B1(n11343), .B2(n9074), 
        .ZN(n9041) );
  OAI22_X1 U9889 ( .A1(data_addr_o_9_), .A2(n9070), .B1(n9805), .B2(n9075), 
        .ZN(n9040) );
  NOR3_X1 U9890 ( .A1(n9042), .A2(n9041), .A3(n9040), .ZN(n9048) );
  XNOR2_X1 U9891 ( .A(n9935), .B(n9271), .ZN(n9047) );
  OAI22_X1 U9892 ( .A1(n9072), .A2(data_addr_o_12_), .B1(data_addr_o_13_), 
        .B2(n9063), .ZN(n9044) );
  OAI22_X1 U9893 ( .A1(n9065), .A2(data_addr_o_14_), .B1(data_addr_o_15_), 
        .B2(n9062), .ZN(n9043) );
  NOR2_X1 U9894 ( .A1(n9044), .A2(n9043), .ZN(n9046) );
  NAND2_X1 U9895 ( .A1(n8444), .A2(n9045), .ZN(n9200) );
  NAND4_X1 U9896 ( .A1(n9048), .A2(n9047), .A3(n9046), .A4(n9200), .ZN(n9052)
         );
  XNOR2_X1 U9897 ( .A(n11312), .B(n9267), .ZN(n9050) );
  XNOR2_X1 U9898 ( .A(data_addr_o_26_), .B(n9264), .ZN(n9049) );
  NAND2_X1 U9899 ( .A1(n9050), .A2(n9049), .ZN(n9051) );
  NOR2_X1 U9900 ( .A1(n9052), .A2(n9051), .ZN(n9055) );
  XNOR2_X1 U9901 ( .A(n11322), .B(n9275), .ZN(n9054) );
  XNOR2_X1 U9902 ( .A(n11303), .B(n9278), .ZN(n9053) );
  NAND4_X1 U9903 ( .A1(n9056), .A2(n9055), .A3(n9054), .A4(n9053), .ZN(n11696)
         );
  XNOR2_X1 U9904 ( .A(n9987), .B(n9057), .ZN(n9069) );
  AND2_X1 U9905 ( .A1(n10493), .A2(n9058), .ZN(n11654) );
  NAND2_X1 U9906 ( .A1(data_addr_o_4_), .A2(n9059), .ZN(n11661) );
  NAND2_X1 U9907 ( .A1(n22), .A2(n9060), .ZN(n11658) );
  OAI211_X1 U9908 ( .C1(n9212), .C2(n10651), .A(n11661), .B(n11658), .ZN(n9061) );
  NOR2_X1 U9909 ( .A1(n11654), .A2(n9061), .ZN(n9067) );
  NAND2_X1 U9910 ( .A1(n11309), .A2(n9062), .ZN(n11647) );
  NAND2_X1 U9911 ( .A1(data_addr_o_13_), .A2(n9063), .ZN(n11646) );
  NAND2_X1 U9912 ( .A1(n9066), .A2(n9065), .ZN(n11657) );
  NAND4_X1 U9913 ( .A1(n9067), .A2(n11647), .A3(n11646), .A4(n11657), .ZN(
        n9068) );
  NOR2_X1 U9914 ( .A1(n9069), .A2(n9068), .ZN(n9080) );
  XNOR2_X1 U9915 ( .A(n12123), .B(n9282), .ZN(n9079) );
  NAND2_X1 U9916 ( .A1(data_addr_o_9_), .A2(n9070), .ZN(n11641) );
  NAND2_X1 U9917 ( .A1(n11331), .A2(n9071), .ZN(n11666) );
  OAI211_X1 U9918 ( .C1(n11291), .C2(n9221), .A(n11641), .B(n11666), .ZN(
        n11687) );
  NAND2_X1 U9919 ( .A1(data_addr_o_12_), .A2(n9072), .ZN(n11678) );
  NAND2_X1 U9920 ( .A1(n8246), .A2(n9073), .ZN(n11674) );
  NAND2_X1 U9921 ( .A1(data_addr_o_10_), .A2(n9074), .ZN(n11640) );
  NAND2_X1 U9922 ( .A1(n10836), .A2(n9075), .ZN(n11652) );
  NAND4_X1 U9923 ( .A1(n11678), .A2(n11674), .A3(n11640), .A4(n11652), .ZN(
        n9076) );
  NOR2_X1 U9924 ( .A1(n11687), .A2(n9076), .ZN(n9078) );
  NAND2_X1 U9925 ( .A1(data_addr_o_17_), .A2(n9077), .ZN(n11688) );
  NAND4_X1 U9926 ( .A1(n9080), .A2(n9079), .A3(n9078), .A4(n11688), .ZN(n9332)
         );
  NOR2_X1 U9927 ( .A1(n7990), .A2(pmp_addr_i[334]), .ZN(n9128) );
  INV_X1 U9928 ( .A(n11227), .ZN(n9125) );
  NOR2_X1 U9929 ( .A1(n9125), .A2(pmp_addr_i[333]), .ZN(n9081) );
  NOR2_X1 U9930 ( .A1(n9128), .A2(n9081), .ZN(n9083) );
  NOR2_X1 U9931 ( .A1(n12184), .A2(pmp_addr_i[336]), .ZN(n9131) );
  NOR2_X1 U9932 ( .A1(n8757), .A2(pmp_addr_i[335]), .ZN(n9082) );
  NOR2_X1 U9933 ( .A1(n9131), .A2(n9082), .ZN(n9133) );
  NAND2_X1 U9934 ( .A1(n9083), .A2(n9133), .ZN(n9137) );
  NOR2_X1 U9935 ( .A1(n10711), .A2(pmp_addr_i[329]), .ZN(n9084) );
  NOR2_X1 U9936 ( .A1(n7472), .A2(pmp_addr_i[330]), .ZN(n9118) );
  NOR2_X1 U9937 ( .A1(n9084), .A2(n9118), .ZN(n9086) );
  NOR2_X1 U9938 ( .A1(n11006), .A2(pmp_addr_i[331]), .ZN(n9085) );
  NOR2_X1 U9939 ( .A1(n10000), .A2(pmp_addr_i[332]), .ZN(n9121) );
  NOR2_X1 U9940 ( .A1(n9085), .A2(n9121), .ZN(n9124) );
  NAND2_X1 U9941 ( .A1(n9086), .A2(n9124), .ZN(n9087) );
  NOR2_X1 U9942 ( .A1(n9137), .A2(n9087), .ZN(n9140) );
  OR2_X1 U9943 ( .A1(pmp_addr_i[321]), .A2(n10010), .ZN(n9090) );
  AND2_X1 U9944 ( .A1(pmp_addr_i[320]), .A2(n10651), .ZN(n9089) );
  AND2_X1 U9945 ( .A1(pmp_addr_i[321]), .A2(n10010), .ZN(n9088) );
  AOI21_X1 U9946 ( .B1(n9090), .B2(n9089), .A(n9088), .ZN(n9093) );
  NOR2_X1 U9947 ( .A1(pmp_addr_i[322]), .A2(n8406), .ZN(n9092) );
  NAND2_X1 U9948 ( .A1(pmp_addr_i[322]), .A2(n6123), .ZN(n9091) );
  OAI21_X1 U9949 ( .B1(n9093), .B2(n9092), .A(n9091), .ZN(n9100) );
  NOR2_X1 U9950 ( .A1(n6127), .A2(pmp_addr_i[323]), .ZN(n9094) );
  NOR2_X1 U9951 ( .A1(n9363), .A2(pmp_addr_i[324]), .ZN(n9097) );
  NOR2_X1 U9952 ( .A1(n9094), .A2(n9097), .ZN(n9099) );
  NAND2_X1 U9953 ( .A1(n6127), .A2(pmp_addr_i[323]), .ZN(n9096) );
  NAND2_X1 U9954 ( .A1(n9363), .A2(pmp_addr_i[324]), .ZN(n9095) );
  OAI21_X1 U9955 ( .B1(n9097), .B2(n9096), .A(n9095), .ZN(n9098) );
  AOI21_X1 U9956 ( .B1(n9100), .B2(n9099), .A(n9098), .ZN(n9115) );
  NOR2_X1 U9957 ( .A1(n8735), .A2(pmp_addr_i[326]), .ZN(n9106) );
  NOR2_X1 U9958 ( .A1(n7152), .A2(pmp_addr_i[325]), .ZN(n9101) );
  NOR2_X1 U9959 ( .A1(n9106), .A2(n9101), .ZN(n9103) );
  NOR2_X1 U9960 ( .A1(n6140), .A2(pmp_addr_i[327]), .ZN(n9102) );
  NOR2_X1 U9961 ( .A1(n7964), .A2(pmp_addr_i[328]), .ZN(n9109) );
  NOR2_X1 U9962 ( .A1(n9102), .A2(n9109), .ZN(n9112) );
  NAND2_X1 U9963 ( .A1(n9103), .A2(n9112), .ZN(n9114) );
  NAND2_X1 U9964 ( .A1(n10697), .A2(pmp_addr_i[325]), .ZN(n9105) );
  NAND2_X1 U9965 ( .A1(n8735), .A2(pmp_addr_i[326]), .ZN(n9104) );
  OAI21_X1 U9966 ( .B1(n9106), .B2(n9105), .A(n9104), .ZN(n9111) );
  NAND2_X1 U9967 ( .A1(n10501), .A2(pmp_addr_i[327]), .ZN(n9108) );
  NAND2_X1 U9968 ( .A1(n7820), .A2(pmp_addr_i[328]), .ZN(n9107) );
  OAI21_X1 U9969 ( .B1(n9109), .B2(n9108), .A(n9107), .ZN(n9110) );
  AOI21_X1 U9970 ( .B1(n9112), .B2(n9111), .A(n9110), .ZN(n9113) );
  OAI21_X1 U9971 ( .B1(n9115), .B2(n9114), .A(n9113), .ZN(n9139) );
  NAND2_X1 U9972 ( .A1(n7324), .A2(pmp_addr_i[329]), .ZN(n9117) );
  NAND2_X1 U9973 ( .A1(n7976), .A2(pmp_addr_i[330]), .ZN(n9116) );
  OAI21_X1 U9974 ( .B1(n9118), .B2(n9117), .A(n9116), .ZN(n9123) );
  NAND2_X1 U9975 ( .A1(n10342), .A2(pmp_addr_i[331]), .ZN(n9120) );
  NAND2_X1 U9976 ( .A1(n10000), .A2(pmp_addr_i[332]), .ZN(n9119) );
  OAI21_X1 U9977 ( .B1(n9121), .B2(n9120), .A(n9119), .ZN(n9122) );
  AOI21_X1 U9978 ( .B1(n9124), .B2(n9123), .A(n9122), .ZN(n9136) );
  NAND2_X1 U9979 ( .A1(n9125), .A2(pmp_addr_i[333]), .ZN(n9127) );
  NAND2_X1 U9980 ( .A1(n10047), .A2(pmp_addr_i[334]), .ZN(n9126) );
  OAI21_X1 U9981 ( .B1(n9128), .B2(n9127), .A(n9126), .ZN(n9134) );
  NAND2_X1 U9982 ( .A1(n8757), .A2(pmp_addr_i[335]), .ZN(n9130) );
  NAND2_X1 U9983 ( .A1(n12184), .A2(pmp_addr_i[336]), .ZN(n9129) );
  OAI21_X1 U9984 ( .B1(n9131), .B2(n9130), .A(n9129), .ZN(n9132) );
  AOI21_X1 U9985 ( .B1(n9134), .B2(n9133), .A(n9132), .ZN(n9135) );
  OAI21_X1 U9986 ( .B1(n9137), .B2(n9136), .A(n9135), .ZN(n9138) );
  AOI21_X1 U9987 ( .B1(n9140), .B2(n9139), .A(n9138), .ZN(n9196) );
  NOR2_X1 U9988 ( .A1(n10764), .A2(pmp_addr_i[341]), .ZN(n9141) );
  INV_X1 U9989 ( .A(data_addr_i[24]), .ZN(n9163) );
  NOR2_X1 U9990 ( .A1(n9163), .A2(pmp_addr_i[342]), .ZN(n9166) );
  NOR2_X1 U9991 ( .A1(n9141), .A2(n9166), .ZN(n9143) );
  NOR2_X1 U9992 ( .A1(n10429), .A2(pmp_addr_i[343]), .ZN(n9142) );
  NOR2_X1 U9993 ( .A1(n6202), .A2(pmp_addr_i[344]), .ZN(n9169) );
  NOR2_X1 U9994 ( .A1(n9142), .A2(n9169), .ZN(n9172) );
  NAND2_X1 U9995 ( .A1(n9143), .A2(n9172), .ZN(n9174) );
  NOR2_X1 U9996 ( .A1(n6192), .A2(pmp_addr_i[339]), .ZN(n9144) );
  INV_X1 U9997 ( .A(data_addr_i[22]), .ZN(n9156) );
  NOR2_X1 U9998 ( .A1(n9156), .A2(pmp_addr_i[340]), .ZN(n9159) );
  NOR2_X1 U9999 ( .A1(n9144), .A2(n9159), .ZN(n9162) );
  NOR2_X1 U10000 ( .A1(n9414), .A2(pmp_addr_i[337]), .ZN(n9145) );
  NOR2_X1 U10001 ( .A1(n10754), .A2(pmp_addr_i[338]), .ZN(n9155) );
  NOR2_X1 U10002 ( .A1(n9145), .A2(n9155), .ZN(n9146) );
  NAND2_X1 U10003 ( .A1(n9162), .A2(n9146), .ZN(n9147) );
  NOR2_X1 U10004 ( .A1(n9174), .A2(n9147), .ZN(n9152) );
  NOR2_X1 U10005 ( .A1(n9438), .A2(pmp_addr_i[345]), .ZN(n9148) );
  NOR2_X1 U10006 ( .A1(n10443), .A2(pmp_addr_i[346]), .ZN(n9178) );
  NOR2_X1 U10007 ( .A1(n9148), .A2(n9178), .ZN(n9150) );
  NOR2_X1 U10008 ( .A1(n10782), .A2(pmp_addr_i[347]), .ZN(n9149) );
  NOR2_X1 U10009 ( .A1(n8494), .A2(pmp_addr_i[348]), .ZN(n9181) );
  NOR2_X1 U10010 ( .A1(n9149), .A2(n9181), .ZN(n9184) );
  NAND2_X1 U10011 ( .A1(n9150), .A2(n9184), .ZN(n9151) );
  NOR2_X1 U10012 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[349]), .ZN(n9189)
         );
  NOR2_X1 U10013 ( .A1(n9151), .A2(n9189), .ZN(n9192) );
  NAND2_X1 U10014 ( .A1(n9152), .A2(n9192), .ZN(n9195) );
  NAND2_X1 U10015 ( .A1(n9414), .A2(pmp_addr_i[337]), .ZN(n9154) );
  NAND2_X1 U10016 ( .A1(n10754), .A2(pmp_addr_i[338]), .ZN(n9153) );
  OAI21_X1 U10017 ( .B1(n9155), .B2(n9154), .A(n9153), .ZN(n9161) );
  NAND2_X1 U10018 ( .A1(n9418), .A2(pmp_addr_i[339]), .ZN(n9158) );
  NAND2_X1 U10019 ( .A1(n9156), .A2(pmp_addr_i[340]), .ZN(n9157) );
  OAI21_X1 U10020 ( .B1(n9159), .B2(n9158), .A(n9157), .ZN(n9160) );
  AOI21_X1 U10021 ( .B1(n9162), .B2(n9161), .A(n9160), .ZN(n9175) );
  NAND2_X1 U10022 ( .A1(n10764), .A2(pmp_addr_i[341]), .ZN(n9165) );
  NAND2_X1 U10023 ( .A1(n9163), .A2(pmp_addr_i[342]), .ZN(n9164) );
  OAI21_X1 U10024 ( .B1(n9166), .B2(n9165), .A(n9164), .ZN(n9171) );
  NAND2_X1 U10025 ( .A1(n6462), .A2(pmp_addr_i[343]), .ZN(n9168) );
  NAND2_X1 U10026 ( .A1(n6202), .A2(pmp_addr_i[344]), .ZN(n9167) );
  OAI21_X1 U10027 ( .B1(n9169), .B2(n9168), .A(n9167), .ZN(n9170) );
  AOI21_X1 U10028 ( .B1(n9172), .B2(n9171), .A(n9170), .ZN(n9173) );
  OAI21_X1 U10029 ( .B1(n9175), .B2(n9174), .A(n9173), .ZN(n9193) );
  NAND2_X1 U10030 ( .A1(n9438), .A2(pmp_addr_i[345]), .ZN(n9177) );
  NAND2_X1 U10031 ( .A1(n8807), .A2(pmp_addr_i[346]), .ZN(n9176) );
  OAI21_X1 U10032 ( .B1(n9178), .B2(n9177), .A(n9176), .ZN(n9183) );
  NAND2_X1 U10033 ( .A1(n10782), .A2(pmp_addr_i[347]), .ZN(n9180) );
  NAND2_X1 U10034 ( .A1(n8814), .A2(pmp_addr_i[348]), .ZN(n9179) );
  OAI21_X1 U10035 ( .B1(n9181), .B2(n9180), .A(n9179), .ZN(n9182) );
  AOI21_X1 U10036 ( .B1(n9184), .B2(n9183), .A(n9182), .ZN(n9190) );
  NAND2_X1 U10037 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[349]), .ZN(n9186)
         );
  INV_X1 U10038 ( .A(pmp_addr_i[350]), .ZN(n9185) );
  NAND2_X1 U10039 ( .A1(n9186), .A2(n9185), .ZN(n9187) );
  NOR2_X1 U10040 ( .A1(n9187), .A2(pmp_addr_i[351]), .ZN(n9188) );
  OAI21_X1 U10041 ( .B1(n9190), .B2(n9189), .A(n9188), .ZN(n9191) );
  AOI21_X1 U10042 ( .B1(n9193), .B2(n9192), .A(n9191), .ZN(n9194) );
  OAI21_X1 U10043 ( .B1(n9196), .B2(n9195), .A(n9194), .ZN(n9330) );
  NOR2_X1 U10044 ( .A1(n9987), .A2(n9057), .ZN(n9248) );
  NOR2_X1 U10045 ( .A1(data_addr_o_15_), .A2(n9062), .ZN(n9198) );
  NOR2_X1 U10046 ( .A1(n9248), .A2(n9198), .ZN(n9202) );
  NOR2_X1 U10047 ( .A1(n10857), .A2(n884), .ZN(n9250) );
  INV_X1 U10048 ( .A(n9200), .ZN(n9201) );
  NOR2_X1 U10049 ( .A1(n9250), .A2(n9201), .ZN(n9253) );
  NAND2_X1 U10050 ( .A1(n9202), .A2(n9253), .ZN(n9256) );
  NOR2_X1 U10051 ( .A1(n10508), .A2(n9073), .ZN(n9205) );
  NOR2_X1 U10052 ( .A1(n31), .A2(n9072), .ZN(n9242) );
  NOR2_X1 U10053 ( .A1(n9205), .A2(n9242), .ZN(n9209) );
  NOR2_X1 U10054 ( .A1(n10847), .A2(n9063), .ZN(n9208) );
  NOR2_X1 U10055 ( .A1(n10848), .A2(n9065), .ZN(n9243) );
  NOR2_X1 U10056 ( .A1(n9208), .A2(n9243), .ZN(n9246) );
  NAND2_X1 U10057 ( .A1(n9209), .A2(n9246), .ZN(n9210) );
  NOR2_X1 U10058 ( .A1(n9256), .A2(n9210), .ZN(n9259) );
  OR2_X1 U10059 ( .A1(n10129), .A2(n9035), .ZN(n9216) );
  OR2_X1 U10060 ( .A1(n10130), .A2(n9060), .ZN(n9215) );
  AND2_X1 U10061 ( .A1(n10130), .A2(n9060), .ZN(n9214) );
  AOI21_X1 U10062 ( .B1(n9216), .B2(n9215), .A(n9214), .ZN(n9219) );
  NOR2_X1 U10063 ( .A1(n10135), .A2(n9059), .ZN(n9218) );
  OAI21_X1 U10064 ( .B1(n9219), .B2(n9218), .A(n11661), .ZN(n9225) );
  NOR2_X1 U10065 ( .A1(n10655), .A2(n9071), .ZN(n9223) );
  NAND2_X1 U10066 ( .A1(n10824), .A2(n9034), .ZN(n9222) );
  OAI21_X1 U10067 ( .B1(n9223), .B2(n9222), .A(n11666), .ZN(n9224) );
  AOI21_X1 U10068 ( .B1(n9039), .B2(n9225), .A(n9224), .ZN(n9241) );
  NOR2_X1 U10069 ( .A1(n10836), .A2(n9075), .ZN(n9234) );
  NOR2_X1 U10070 ( .A1(n10493), .A2(n9058), .ZN(n9228) );
  NOR2_X1 U10071 ( .A1(n9234), .A2(n9228), .ZN(n9232) );
  NOR2_X1 U10072 ( .A1(data_addr_o_9_), .A2(n9070), .ZN(n9231) );
  NOR2_X1 U10073 ( .A1(data_addr_o_10_), .A2(n9074), .ZN(n9235) );
  NOR2_X1 U10074 ( .A1(n9231), .A2(n9235), .ZN(n9238) );
  NAND2_X1 U10075 ( .A1(n9232), .A2(n9238), .ZN(n9240) );
  NAND2_X1 U10076 ( .A1(data_addr_o_7_), .A2(n9058), .ZN(n9233) );
  OAI21_X1 U10077 ( .B1(n9234), .B2(n9233), .A(n11652), .ZN(n9237) );
  OAI21_X1 U10078 ( .B1(n9235), .B2(n11641), .A(n11640), .ZN(n9236) );
  AOI21_X1 U10079 ( .B1(n9238), .B2(n9237), .A(n9236), .ZN(n9239) );
  OAI21_X1 U10080 ( .B1(n9241), .B2(n9240), .A(n9239), .ZN(n9258) );
  OAI21_X1 U10081 ( .B1(n9242), .B2(n11674), .A(n11678), .ZN(n9245) );
  OAI21_X1 U10082 ( .B1(n9243), .B2(n11646), .A(n11657), .ZN(n9244) );
  AOI21_X1 U10083 ( .B1(n9246), .B2(n9245), .A(n9244), .ZN(n9255) );
  NAND2_X1 U10084 ( .A1(n9987), .A2(n9057), .ZN(n9247) );
  OAI21_X1 U10085 ( .B1(n9248), .B2(n11647), .A(n9247), .ZN(n9252) );
  NAND2_X1 U10086 ( .A1(n10857), .A2(n884), .ZN(n9249) );
  OAI21_X1 U10087 ( .B1(n9250), .B2(n11688), .A(n9249), .ZN(n9251) );
  AOI21_X1 U10088 ( .B1(n9253), .B2(n9252), .A(n9251), .ZN(n9254) );
  OAI21_X1 U10089 ( .B1(n9256), .B2(n9255), .A(n9254), .ZN(n9257) );
  AOI21_X1 U10090 ( .B1(n9259), .B2(n9258), .A(n9257), .ZN(n9327) );
  NOR2_X1 U10091 ( .A1(n10898), .A2(n1022), .ZN(n9262) );
  NOR2_X1 U10092 ( .A1(n10738), .A2(n958), .ZN(n9298) );
  NOR2_X1 U10093 ( .A1(n9262), .A2(n9298), .ZN(n9266) );
  NOR2_X1 U10094 ( .A1(n9923), .A2(n1025), .ZN(n9265) );
  NOR2_X1 U10095 ( .A1(n10267), .A2(n951), .ZN(n9301) );
  NOR2_X1 U10096 ( .A1(n9265), .A2(n9301), .ZN(n9304) );
  NAND2_X1 U10097 ( .A1(n9266), .A2(n9304), .ZN(n9306) );
  NOR2_X1 U10098 ( .A1(n10202), .A2(n998), .ZN(n9269) );
  NOR2_X1 U10099 ( .A1(n9915), .A2(n964), .ZN(n9292) );
  NOR2_X1 U10100 ( .A1(n9269), .A2(n9292), .ZN(n9295) );
  NOR2_X1 U10101 ( .A1(n11283), .A2(n994), .ZN(n9272) );
  NOR2_X1 U10102 ( .A1(data_addr_o_20_), .A2(n969), .ZN(n9289) );
  NOR2_X1 U10103 ( .A1(n9272), .A2(n9289), .ZN(n9273) );
  NAND2_X1 U10104 ( .A1(n9295), .A2(n9273), .ZN(n9274) );
  NOR2_X1 U10105 ( .A1(n9306), .A2(n9274), .ZN(n9286) );
  NOR2_X1 U10106 ( .A1(n10746), .A2(n1006), .ZN(n9277) );
  NOR2_X1 U10107 ( .A1(n10914), .A2(n980), .ZN(n9310) );
  NOR2_X1 U10108 ( .A1(n9277), .A2(n9310), .ZN(n9281) );
  NOR2_X1 U10109 ( .A1(n9955), .A2(n1009), .ZN(n9280) );
  NOR2_X1 U10110 ( .A1(n10919), .A2(n974), .ZN(n9313) );
  NOR2_X1 U10111 ( .A1(n9280), .A2(n9313), .ZN(n9316) );
  NAND2_X1 U10112 ( .A1(n9281), .A2(n9316), .ZN(n9285) );
  NOR2_X1 U10113 ( .A1(n24), .A2(n1034), .ZN(n9283) );
  NOR2_X1 U10114 ( .A1(n9283), .A2(pmp_addr_i[318]), .ZN(n9284) );
  NAND2_X1 U10115 ( .A1(n9284), .A2(n985), .ZN(n9320) );
  NOR2_X1 U10116 ( .A1(n9285), .A2(n9320), .ZN(n9323) );
  NAND2_X1 U10117 ( .A1(n9286), .A2(n9323), .ZN(n9326) );
  NAND2_X1 U10118 ( .A1(n10886), .A2(n994), .ZN(n9288) );
  NAND2_X1 U10119 ( .A1(data_addr_o_20_), .A2(n969), .ZN(n9287) );
  OAI21_X1 U10120 ( .B1(n9289), .B2(n9288), .A(n9287), .ZN(n9294) );
  NAND2_X1 U10121 ( .A1(n10202), .A2(n998), .ZN(n9291) );
  NAND2_X1 U10122 ( .A1(n9915), .A2(n964), .ZN(n9290) );
  OAI21_X1 U10123 ( .B1(n9292), .B2(n9291), .A(n9290), .ZN(n9293) );
  AOI21_X1 U10124 ( .B1(n9295), .B2(n9294), .A(n9293), .ZN(n9307) );
  NAND2_X1 U10125 ( .A1(n10898), .A2(n1022), .ZN(n9297) );
  NAND2_X1 U10126 ( .A1(n10738), .A2(n958), .ZN(n9296) );
  OAI21_X1 U10127 ( .B1(n9298), .B2(n9297), .A(n9296), .ZN(n9303) );
  NAND2_X1 U10128 ( .A1(n9923), .A2(n1025), .ZN(n9300) );
  NAND2_X1 U10129 ( .A1(n10267), .A2(n951), .ZN(n9299) );
  OAI21_X1 U10130 ( .B1(n9301), .B2(n9300), .A(n9299), .ZN(n9302) );
  AOI21_X1 U10131 ( .B1(n9304), .B2(n9303), .A(n9302), .ZN(n9305) );
  OAI21_X1 U10132 ( .B1(n9307), .B2(n9306), .A(n9305), .ZN(n9324) );
  NAND2_X1 U10133 ( .A1(n10746), .A2(n1006), .ZN(n9309) );
  NAND2_X1 U10134 ( .A1(n10914), .A2(n980), .ZN(n9308) );
  OAI21_X1 U10135 ( .B1(n9310), .B2(n9309), .A(n9308), .ZN(n9315) );
  NAND2_X1 U10136 ( .A1(n9955), .A2(n1009), .ZN(n9312) );
  NAND2_X1 U10137 ( .A1(n10919), .A2(n974), .ZN(n9311) );
  OAI21_X1 U10138 ( .B1(n9313), .B2(n9312), .A(n9311), .ZN(n9314) );
  AOI21_X1 U10139 ( .B1(n9316), .B2(n9315), .A(n9314), .ZN(n9321) );
  NAND2_X1 U10140 ( .A1(n24), .A2(n1034), .ZN(n9317) );
  NOR2_X1 U10141 ( .A1(n9317), .A2(pmp_addr_i[318]), .ZN(n9318) );
  NAND2_X1 U10142 ( .A1(n9318), .A2(n985), .ZN(n9319) );
  OAI21_X1 U10143 ( .B1(n9321), .B2(n9320), .A(n9319), .ZN(n9322) );
  AOI21_X1 U10144 ( .B1(n9324), .B2(n9323), .A(n9322), .ZN(n9325) );
  OAI21_X1 U10145 ( .B1(n9327), .B2(n9326), .A(n9325), .ZN(n9328) );
  NAND3_X1 U10146 ( .A1(n9330), .A2(n9329), .A3(n9328), .ZN(n9331) );
  OAI21_X1 U10147 ( .B1(n11696), .B2(n9332), .A(n9331), .ZN(n9335) );
  MUX2_X1 U10148 ( .A(pmp_cfg_i[80]), .B(pmp_cfg_i[81]), .S(n11019), .Z(n9334)
         );
  AND2_X1 U10149 ( .A1(n9333), .A2(n9334), .ZN(n11684) );
  NAND2_X1 U10150 ( .A1(n9335), .A2(n11684), .ZN(n9336) );
  NOR2_X1 U10152 ( .A1(pmp_addr_i[140]), .A2(n6154), .ZN(n9342) );
  INV_X1 U10153 ( .A(n11227), .ZN(n10338) );
  NOR2_X1 U10154 ( .A1(pmp_addr_i[141]), .A2(n10338), .ZN(n9388) );
  NOR2_X1 U10155 ( .A1(n9342), .A2(n9388), .ZN(n9344) );
  NOR2_X1 U10156 ( .A1(pmp_addr_i[142]), .A2(n7057), .ZN(n9343) );
  NOR2_X1 U10157 ( .A1(pmp_addr_i[143]), .A2(n8444), .ZN(n9391) );
  NOR2_X1 U10158 ( .A1(n9343), .A2(n9391), .ZN(n9394) );
  NAND2_X1 U10159 ( .A1(n9344), .A2(n9394), .ZN(n9396) );
  NOR2_X1 U10160 ( .A1(pmp_addr_i[137]), .A2(n7324), .ZN(n9379) );
  NOR2_X1 U10161 ( .A1(pmp_addr_i[136]), .A2(n10701), .ZN(n9345) );
  NOR2_X1 U10162 ( .A1(n9379), .A2(n9345), .ZN(n9347) );
  NOR2_X1 U10163 ( .A1(pmp_addr_i[138]), .A2(n10005), .ZN(n9346) );
  NOR2_X1 U10164 ( .A1(pmp_addr_i[139]), .A2(n10342), .ZN(n9382) );
  NOR2_X1 U10165 ( .A1(n9346), .A2(n9382), .ZN(n9385) );
  NAND2_X1 U10166 ( .A1(n9347), .A2(n9385), .ZN(n9348) );
  NOR2_X1 U10167 ( .A1(n9396), .A2(n9348), .ZN(n9400) );
  NOR2_X1 U10168 ( .A1(pmp_addr_i[131]), .A2(n10346), .ZN(n9356) );
  NOR2_X1 U10169 ( .A1(pmp_addr_i[130]), .A2(n6123), .ZN(n9349) );
  NOR2_X1 U10170 ( .A1(n9356), .A2(n9349), .ZN(n9359) );
  NOR2_X1 U10171 ( .A1(pmp_addr_i[129]), .A2(n9350), .ZN(n9353) );
  NAND2_X1 U10172 ( .A1(pmp_addr_i[128]), .A2(n10651), .ZN(n9352) );
  NAND2_X1 U10173 ( .A1(pmp_addr_i[129]), .A2(n9350), .ZN(n9351) );
  OAI21_X1 U10174 ( .B1(n9353), .B2(n9352), .A(n9351), .ZN(n9358) );
  NAND2_X1 U10175 ( .A1(pmp_addr_i[130]), .A2(n6123), .ZN(n9355) );
  NAND2_X1 U10176 ( .A1(pmp_addr_i[131]), .A2(n10346), .ZN(n9354) );
  OAI21_X1 U10177 ( .B1(n9356), .B2(n9355), .A(n9354), .ZN(n9357) );
  AOI21_X1 U10178 ( .B1(n9359), .B2(n9358), .A(n9357), .ZN(n9376) );
  INV_X1 U10179 ( .A(n10655), .ZN(n9363) );
  NOR2_X1 U10180 ( .A1(pmp_addr_i[132]), .A2(n9363), .ZN(n9360) );
  NOR2_X1 U10181 ( .A1(pmp_addr_i[133]), .A2(n6400), .ZN(n9366) );
  NOR2_X1 U10182 ( .A1(n9360), .A2(n9366), .ZN(n9362) );
  NOR2_X1 U10183 ( .A1(pmp_addr_i[134]), .A2(n8735), .ZN(n9361) );
  NOR2_X1 U10184 ( .A1(pmp_addr_i[135]), .A2(n9367), .ZN(n9370) );
  NOR2_X1 U10185 ( .A1(n9361), .A2(n9370), .ZN(n9373) );
  NAND2_X1 U10186 ( .A1(n9362), .A2(n9373), .ZN(n9375) );
  NAND2_X1 U10187 ( .A1(pmp_addr_i[132]), .A2(n9363), .ZN(n9365) );
  NAND2_X1 U10188 ( .A1(pmp_addr_i[133]), .A2(n7152), .ZN(n9364) );
  OAI21_X1 U10189 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(n9372) );
  NAND2_X1 U10190 ( .A1(pmp_addr_i[134]), .A2(n8735), .ZN(n9369) );
  NAND2_X1 U10191 ( .A1(pmp_addr_i[135]), .A2(n9367), .ZN(n9368) );
  OAI21_X1 U10192 ( .B1(n9370), .B2(n9369), .A(n9368), .ZN(n9371) );
  AOI21_X1 U10193 ( .B1(n9373), .B2(n9372), .A(n9371), .ZN(n9374) );
  OAI21_X1 U10194 ( .B1(n9376), .B2(n9375), .A(n9374), .ZN(n9399) );
  NAND2_X1 U10195 ( .A1(pmp_addr_i[136]), .A2(n10701), .ZN(n9378) );
  NAND2_X1 U10196 ( .A1(pmp_addr_i[137]), .A2(n9508), .ZN(n9377) );
  OAI21_X1 U10197 ( .B1(n9379), .B2(n9378), .A(n9377), .ZN(n9384) );
  NAND2_X1 U10198 ( .A1(pmp_addr_i[138]), .A2(n7976), .ZN(n9381) );
  NAND2_X1 U10199 ( .A1(pmp_addr_i[139]), .A2(n11006), .ZN(n9380) );
  OAI21_X1 U10200 ( .B1(n9382), .B2(n9381), .A(n9380), .ZN(n9383) );
  AOI21_X1 U10201 ( .B1(n9385), .B2(n9384), .A(n9383), .ZN(n9397) );
  NAND2_X1 U10202 ( .A1(pmp_addr_i[140]), .A2(n10000), .ZN(n9387) );
  NAND2_X1 U10203 ( .A1(pmp_addr_i[141]), .A2(n10338), .ZN(n9386) );
  OAI21_X1 U10204 ( .B1(n9388), .B2(n9387), .A(n9386), .ZN(n9393) );
  NAND2_X1 U10205 ( .A1(pmp_addr_i[142]), .A2(n10047), .ZN(n9390) );
  NAND2_X1 U10206 ( .A1(pmp_addr_i[143]), .A2(n8444), .ZN(n9389) );
  OAI21_X1 U10207 ( .B1(n9391), .B2(n9390), .A(n9389), .ZN(n9392) );
  AOI21_X1 U10208 ( .B1(n9394), .B2(n9393), .A(n9392), .ZN(n9395) );
  OAI21_X1 U10209 ( .B1(n9397), .B2(n9396), .A(n9395), .ZN(n9398) );
  AOI21_X1 U10210 ( .B1(n9400), .B2(n9399), .A(n9398), .ZN(n9462) );
  NOR2_X1 U10211 ( .A1(pmp_addr_i[144]), .A2(n10403), .ZN(n9401) );
  INV_X1 U10212 ( .A(data_addr_i[19]), .ZN(n9414) );
  NOR2_X1 U10213 ( .A1(pmp_addr_i[145]), .A2(n9414), .ZN(n9417) );
  NOR2_X1 U10214 ( .A1(n9401), .A2(n9417), .ZN(n9403) );
  NOR2_X1 U10215 ( .A1(pmp_addr_i[146]), .A2(n6188), .ZN(n9402) );
  INV_X1 U10216 ( .A(data_addr_i[21]), .ZN(n9418) );
  NOR2_X1 U10217 ( .A1(pmp_addr_i[147]), .A2(n9418), .ZN(n9421) );
  NOR2_X1 U10218 ( .A1(n9402), .A2(n9421), .ZN(n9424) );
  NAND2_X1 U10219 ( .A1(n9403), .A2(n9424), .ZN(n9407) );
  INV_X1 U10220 ( .A(data_addr_i[22]), .ZN(n9425) );
  NOR2_X1 U10221 ( .A1(pmp_addr_i[148]), .A2(n9425), .ZN(n9404) );
  NOR2_X1 U10222 ( .A1(pmp_addr_i[149]), .A2(n10764), .ZN(n9428) );
  NOR2_X1 U10223 ( .A1(n9404), .A2(n9428), .ZN(n9406) );
  NOR2_X1 U10224 ( .A1(pmp_addr_i[150]), .A2(n9163), .ZN(n9405) );
  NOR2_X1 U10225 ( .A1(pmp_addr_i[151]), .A2(n10768), .ZN(n9431) );
  NOR2_X1 U10226 ( .A1(n9405), .A2(n9431), .ZN(n9434) );
  NAND2_X1 U10227 ( .A1(n9406), .A2(n9434), .ZN(n9436) );
  NOR2_X1 U10228 ( .A1(n9407), .A2(n9436), .ZN(n9413) );
  NOR2_X1 U10229 ( .A1(pmp_addr_i[154]), .A2(n8807), .ZN(n9408) );
  NOR2_X1 U10230 ( .A1(pmp_addr_i[155]), .A2(n6216), .ZN(n9444) );
  NOR2_X1 U10231 ( .A1(n9408), .A2(n9444), .ZN(n9447) );
  NOR2_X1 U10232 ( .A1(pmp_addr_i[152]), .A2(n10439), .ZN(n9409) );
  INV_X1 U10233 ( .A(data_addr_i[27]), .ZN(n9438) );
  NOR2_X1 U10234 ( .A1(pmp_addr_i[153]), .A2(n9438), .ZN(n9441) );
  NOR2_X1 U10235 ( .A1(n9409), .A2(n9441), .ZN(n9410) );
  NAND2_X1 U10236 ( .A1(n9447), .A2(n9410), .ZN(n9412) );
  NOR2_X1 U10237 ( .A1(pmp_addr_i[156]), .A2(n8814), .ZN(n9411) );
  NOR2_X1 U10238 ( .A1(pmp_addr_i[157]), .A2(n10107), .ZN(n9450) );
  OR2_X1 U10239 ( .A1(n9411), .A2(n9450), .ZN(n9455) );
  NOR2_X1 U10240 ( .A1(n9412), .A2(n9455), .ZN(n9458) );
  NAND2_X1 U10241 ( .A1(n9413), .A2(n9458), .ZN(n9461) );
  NAND2_X1 U10242 ( .A1(pmp_addr_i[144]), .A2(n12184), .ZN(n9416) );
  NAND2_X1 U10243 ( .A1(pmp_addr_i[145]), .A2(n9414), .ZN(n9415) );
  OAI21_X1 U10244 ( .B1(n9417), .B2(n9416), .A(n9415), .ZN(n9423) );
  NAND2_X1 U10245 ( .A1(pmp_addr_i[146]), .A2(n6188), .ZN(n9420) );
  NAND2_X1 U10246 ( .A1(pmp_addr_i[147]), .A2(n9418), .ZN(n9419) );
  OAI21_X1 U10247 ( .B1(n9421), .B2(n9420), .A(n9419), .ZN(n9422) );
  AOI21_X1 U10248 ( .B1(n9424), .B2(n9423), .A(n9422), .ZN(n9437) );
  NAND2_X1 U10249 ( .A1(pmp_addr_i[148]), .A2(n9425), .ZN(n9427) );
  NAND2_X1 U10250 ( .A1(pmp_addr_i[149]), .A2(n10764), .ZN(n9426) );
  OAI21_X1 U10251 ( .B1(n9428), .B2(n9427), .A(n9426), .ZN(n9433) );
  NAND2_X1 U10252 ( .A1(pmp_addr_i[150]), .A2(n9163), .ZN(n9430) );
  NAND2_X1 U10253 ( .A1(pmp_addr_i[151]), .A2(n6462), .ZN(n9429) );
  OAI21_X1 U10254 ( .B1(n9431), .B2(n9430), .A(n9429), .ZN(n9432) );
  AOI21_X1 U10255 ( .B1(n9434), .B2(n9433), .A(n9432), .ZN(n9435) );
  OAI21_X1 U10256 ( .B1(n9437), .B2(n9436), .A(n9435), .ZN(n9459) );
  NAND2_X1 U10257 ( .A1(pmp_addr_i[152]), .A2(n10439), .ZN(n9440) );
  NAND2_X1 U10258 ( .A1(pmp_addr_i[153]), .A2(n9438), .ZN(n9439) );
  OAI21_X1 U10259 ( .B1(n9441), .B2(n9440), .A(n9439), .ZN(n9446) );
  NAND2_X1 U10260 ( .A1(pmp_addr_i[154]), .A2(n8807), .ZN(n9443) );
  NAND2_X1 U10261 ( .A1(pmp_addr_i[155]), .A2(n6216), .ZN(n9442) );
  OAI21_X1 U10262 ( .B1(n9444), .B2(n9443), .A(n9442), .ZN(n9445) );
  AOI21_X1 U10263 ( .B1(n9447), .B2(n9446), .A(n9445), .ZN(n9456) );
  NAND2_X1 U10264 ( .A1(pmp_addr_i[156]), .A2(n8814), .ZN(n9449) );
  NAND2_X1 U10265 ( .A1(pmp_addr_i[157]), .A2(data_addr_o_31__BAR), .ZN(n9448)
         );
  OAI21_X1 U10266 ( .B1(n9450), .B2(n9449), .A(n9448), .ZN(n9453) );
  INV_X1 U10267 ( .A(n9451), .ZN(n9452) );
  NOR2_X1 U10268 ( .A1(n9453), .A2(n9452), .ZN(n9454) );
  OAI21_X1 U10269 ( .B1(n9456), .B2(n9455), .A(n9454), .ZN(n9457) );
  AOI21_X1 U10270 ( .B1(n9459), .B2(n9458), .A(n9457), .ZN(n9460) );
  OAI21_X1 U10271 ( .B1(n9462), .B2(n9461), .A(n9460), .ZN(n9585) );
  NOR2_X1 U10272 ( .A1(n1176), .A2(n10530), .ZN(n9527) );
  NOR2_X1 U10273 ( .A1(n1244), .A2(n11283), .ZN(n9463) );
  NOR2_X1 U10274 ( .A1(n9527), .A2(n9463), .ZN(n9465) );
  NOR2_X1 U10275 ( .A1(n1170), .A2(n9529), .ZN(n9532) );
  INV_X1 U10276 ( .A(n9625), .ZN(n9528) );
  NOR2_X1 U10277 ( .A1(n9528), .A2(n10891), .ZN(n9464) );
  NOR2_X1 U10278 ( .A1(n9532), .A2(n9464), .ZN(n9535) );
  NAND2_X1 U10279 ( .A1(n9465), .A2(n9535), .ZN(n9537) );
  NOR2_X1 U10280 ( .A1(n1194), .A2(n10857), .ZN(n9521) );
  NAND2_X1 U10281 ( .A1(n9519), .A2(n7995), .ZN(n9614) );
  INV_X1 U10282 ( .A(n9614), .ZN(n9466) );
  NOR2_X1 U10283 ( .A1(n9521), .A2(n9466), .ZN(n9524) );
  NOR2_X1 U10284 ( .A1(n1292), .A2(n11309), .ZN(n9467) );
  NOR2_X1 U10285 ( .A1(n1293), .A2(n11014), .ZN(n9518) );
  NOR2_X1 U10286 ( .A1(n9467), .A2(n9518), .ZN(n9468) );
  NAND2_X1 U10287 ( .A1(n9524), .A2(n9468), .ZN(n9469) );
  NOR2_X1 U10288 ( .A1(n9537), .A2(n9469), .ZN(n9541) );
  INV_X1 U10289 ( .A(n9637), .ZN(n9470) );
  NOR2_X1 U10290 ( .A1(data_addr_o_2_), .A2(n9470), .ZN(n9474) );
  INV_X1 U10291 ( .A(n9643), .ZN(n9472) );
  NOR2_X1 U10292 ( .A1(n10818), .A2(n9472), .ZN(n9473) );
  NAND2_X1 U10293 ( .A1(n10818), .A2(n9472), .ZN(n11908) );
  OAI21_X1 U10294 ( .B1(n9474), .B2(n9473), .A(n11908), .ZN(n9477) );
  NAND2_X1 U10295 ( .A1(n12058), .A2(n9475), .ZN(n9646) );
  AND2_X1 U10296 ( .A1(n10479), .A2(n9639), .ZN(n9476) );
  AOI21_X1 U10297 ( .B1(n9477), .B2(n9646), .A(n9476), .ZN(n9486) );
  OR2_X1 U10298 ( .A1(n10824), .A2(n9647), .ZN(n9480) );
  OR2_X1 U10299 ( .A1(n11331), .A2(n9642), .ZN(n9483) );
  NAND2_X1 U10300 ( .A1(n9480), .A2(n9483), .ZN(n9485) );
  AND2_X1 U10301 ( .A1(n10824), .A2(n9647), .ZN(n9482) );
  AND2_X1 U10302 ( .A1(data_addr_o_6_), .A2(n9642), .ZN(n9481) );
  AOI21_X1 U10303 ( .B1(n9483), .B2(n9482), .A(n9481), .ZN(n9484) );
  OAI21_X1 U10304 ( .B1(n9486), .B2(n9485), .A(n9484), .ZN(n9502) );
  OR2_X1 U10305 ( .A1(n10836), .A2(n9606), .ZN(n9494) );
  OR2_X1 U10306 ( .A1(n7816), .A2(n9636), .ZN(n9489) );
  NAND2_X1 U10307 ( .A1(n9494), .A2(n9489), .ZN(n9492) );
  OR2_X1 U10308 ( .A1(n8237), .A2(n9649), .ZN(n9491) );
  NAND2_X1 U10309 ( .A1(n7964), .A2(n9495), .ZN(n9609) );
  NAND2_X1 U10310 ( .A1(n9491), .A2(n9609), .ZN(n9498) );
  NOR2_X1 U10311 ( .A1(n9492), .A2(n9498), .ZN(n9501) );
  AND2_X1 U10312 ( .A1(n7816), .A2(n9636), .ZN(n9493) );
  AND2_X1 U10313 ( .A1(n10836), .A2(n9606), .ZN(n11915) );
  AOI21_X1 U10314 ( .B1(n9494), .B2(n9493), .A(n11915), .ZN(n9499) );
  AND2_X1 U10315 ( .A1(data_addr_o_9_), .A2(n9649), .ZN(n9496) );
  NOR2_X1 U10316 ( .A1(n9495), .A2(n10701), .ZN(n11922) );
  AOI21_X1 U10317 ( .B1(n9609), .B2(n9496), .A(n11922), .ZN(n9497) );
  OAI21_X1 U10318 ( .B1(n9499), .B2(n9498), .A(n9497), .ZN(n9500) );
  AOI21_X1 U10319 ( .B1(n9502), .B2(n9501), .A(n9500), .ZN(n9516) );
  NOR2_X1 U10320 ( .A1(n1288), .A2(n10848), .ZN(n9510) );
  NOR2_X1 U10321 ( .A1(n1287), .A2(n10847), .ZN(n9503) );
  NOR2_X1 U10322 ( .A1(n9510), .A2(n9503), .ZN(n9513) );
  NOR2_X1 U10323 ( .A1(n1285), .A2(n31), .ZN(n9509) );
  NAND2_X1 U10324 ( .A1(n9508), .A2(n9507), .ZN(n9612) );
  INV_X1 U10325 ( .A(n9612), .ZN(n9505) );
  NOR2_X1 U10326 ( .A1(n9509), .A2(n9505), .ZN(n9506) );
  NAND2_X1 U10327 ( .A1(n9513), .A2(n9506), .ZN(n9515) );
  OR2_X1 U10328 ( .A1(n9508), .A2(n9507), .ZN(n11928) );
  OR2_X1 U10329 ( .A1(n9605), .A2(n7472), .ZN(n11933) );
  OAI21_X1 U10330 ( .B1(n9509), .B2(n11928), .A(n11933), .ZN(n9512) );
  OR2_X1 U10331 ( .A1(n9604), .A2(n11006), .ZN(n11893) );
  OR2_X1 U10332 ( .A1(n9616), .A2(n11334), .ZN(n11887) );
  OAI21_X1 U10333 ( .B1(n9510), .B2(n11893), .A(n11887), .ZN(n9511) );
  AOI21_X1 U10334 ( .B1(n9513), .B2(n9512), .A(n9511), .ZN(n9514) );
  OAI21_X1 U10335 ( .B1(n9516), .B2(n9515), .A(n9514), .ZN(n9540) );
  OR2_X1 U10336 ( .A1(n9617), .A2(n9941), .ZN(n11879) );
  NAND2_X1 U10337 ( .A1(n1293), .A2(n11014), .ZN(n9517) );
  OAI21_X1 U10338 ( .B1(n9518), .B2(n11879), .A(n9517), .ZN(n9523) );
  OR2_X1 U10339 ( .A1(n9519), .A2(n8757), .ZN(n11888) );
  NAND2_X1 U10340 ( .A1(n1194), .A2(n10857), .ZN(n9520) );
  OAI21_X1 U10341 ( .B1(n9521), .B2(n11888), .A(n9520), .ZN(n9522) );
  AOI21_X1 U10342 ( .B1(n9524), .B2(n9523), .A(n9522), .ZN(n9538) );
  NAND2_X1 U10343 ( .A1(n1244), .A2(n10886), .ZN(n9526) );
  NAND2_X1 U10344 ( .A1(n1176), .A2(n10530), .ZN(n9525) );
  OAI21_X1 U10345 ( .B1(n9527), .B2(n9526), .A(n9525), .ZN(n9534) );
  NAND2_X1 U10346 ( .A1(n9528), .A2(n10891), .ZN(n9531) );
  NAND2_X1 U10347 ( .A1(n1170), .A2(n9529), .ZN(n9530) );
  OAI21_X1 U10348 ( .B1(n9532), .B2(n9531), .A(n9530), .ZN(n9533) );
  AOI21_X1 U10349 ( .B1(n9535), .B2(n9534), .A(n9533), .ZN(n9536) );
  OAI21_X1 U10350 ( .B1(n9538), .B2(n9537), .A(n9536), .ZN(n9539) );
  AOI21_X1 U10351 ( .B1(n9541), .B2(n9540), .A(n9539), .ZN(n9582) );
  INV_X1 U10352 ( .A(n9587), .ZN(n9553) );
  NOR2_X1 U10353 ( .A1(n9553), .A2(n10738), .ZN(n9556) );
  NOR2_X1 U10354 ( .A1(n1268), .A2(n10898), .ZN(n9542) );
  NOR2_X1 U10355 ( .A1(n9556), .A2(n9542), .ZN(n9544) );
  NOR2_X1 U10356 ( .A1(n1185), .A2(n10267), .ZN(n9559) );
  NOR2_X1 U10357 ( .A1(n1272), .A2(n9923), .ZN(n9543) );
  NOR2_X1 U10358 ( .A1(n9559), .A2(n9543), .ZN(n9562) );
  NAND2_X1 U10359 ( .A1(n9544), .A2(n9562), .ZN(n9548) );
  NOR2_X1 U10360 ( .A1(n1156), .A2(n10914), .ZN(n9565) );
  NOR2_X1 U10361 ( .A1(n1253), .A2(n10746), .ZN(n9545) );
  NOR2_X1 U10362 ( .A1(n9565), .A2(n9545), .ZN(n9547) );
  NOR2_X1 U10363 ( .A1(n1162), .A2(data_addr_o_30_), .ZN(n9568) );
  NOR2_X1 U10364 ( .A1(n1256), .A2(n10918), .ZN(n9546) );
  NOR2_X1 U10365 ( .A1(n9568), .A2(n9546), .ZN(n9571) );
  NAND2_X1 U10366 ( .A1(n9547), .A2(n9571), .ZN(n9573) );
  NOR2_X1 U10367 ( .A1(n9548), .A2(n9573), .ZN(n9552) );
  OR2_X1 U10368 ( .A1(n1278), .A2(n24), .ZN(n9550) );
  NAND2_X1 U10369 ( .A1(n9550), .A2(n7539), .ZN(n9551) );
  NOR2_X1 U10370 ( .A1(n9551), .A2(pmp_addr_i[127]), .ZN(n9578) );
  NAND2_X1 U10371 ( .A1(n9552), .A2(n9578), .ZN(n9581) );
  NAND2_X1 U10372 ( .A1(n1268), .A2(n10898), .ZN(n9555) );
  NAND2_X1 U10373 ( .A1(n9553), .A2(n10738), .ZN(n9554) );
  OAI21_X1 U10374 ( .B1(n9556), .B2(n9555), .A(n9554), .ZN(n9561) );
  NAND2_X1 U10375 ( .A1(n1272), .A2(n9923), .ZN(n9558) );
  NAND2_X1 U10376 ( .A1(n1185), .A2(n10267), .ZN(n9557) );
  OAI21_X1 U10377 ( .B1(n9559), .B2(n9558), .A(n9557), .ZN(n9560) );
  AOI21_X1 U10378 ( .B1(n9562), .B2(n9561), .A(n9560), .ZN(n9574) );
  NAND2_X1 U10379 ( .A1(n1253), .A2(n10746), .ZN(n9564) );
  NAND2_X1 U10380 ( .A1(n1156), .A2(n10914), .ZN(n9563) );
  OAI21_X1 U10381 ( .B1(n9565), .B2(n9564), .A(n9563), .ZN(n9570) );
  NAND2_X1 U10382 ( .A1(n1256), .A2(n10918), .ZN(n9567) );
  NAND2_X1 U10383 ( .A1(n1162), .A2(n10919), .ZN(n9566) );
  OAI21_X1 U10384 ( .B1(n9568), .B2(n9567), .A(n9566), .ZN(n9569) );
  AOI21_X1 U10385 ( .B1(n9571), .B2(n9570), .A(n9569), .ZN(n9572) );
  OAI21_X1 U10386 ( .B1(n9574), .B2(n9573), .A(n9572), .ZN(n9579) );
  AND2_X1 U10387 ( .A1(n1278), .A2(n24), .ZN(n9575) );
  NAND2_X1 U10388 ( .A1(n9575), .A2(n7539), .ZN(n9576) );
  NOR2_X1 U10389 ( .A1(n9576), .A2(pmp_addr_i[127]), .ZN(n9577) );
  AOI21_X1 U10390 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(n9580) );
  OAI21_X1 U10391 ( .B1(n9582), .B2(n9581), .A(n9580), .ZN(n9583) );
  NAND3_X1 U10392 ( .A1(n9585), .A2(n9584), .A3(n9583), .ZN(n9661) );
  XNOR2_X1 U10393 ( .A(n9586), .B(n11322), .ZN(n9593) );
  XNOR2_X1 U10394 ( .A(n9587), .B(n10899), .ZN(n9592) );
  XNOR2_X1 U10395 ( .A(n9588), .B(n9935), .ZN(n9591) );
  XNOR2_X1 U10396 ( .A(n9589), .B(data_addr_o_26_), .ZN(n9590) );
  NAND4_X1 U10397 ( .A1(n9593), .A2(n9592), .A3(n9591), .A4(n9590), .ZN(n9603)
         );
  XNOR2_X1 U10398 ( .A(n9594), .B(data_addr_o_23_), .ZN(n9601) );
  XNOR2_X1 U10399 ( .A(n9595), .B(n11283), .ZN(n9600) );
  XNOR2_X1 U10400 ( .A(n9596), .B(n11298), .ZN(n9599) );
  XNOR2_X1 U10401 ( .A(n9597), .B(data_addr_o_30_), .ZN(n9598) );
  NAND4_X1 U10402 ( .A1(n9601), .A2(n9600), .A3(n9599), .A4(n9598), .ZN(n9602)
         );
  NOR2_X1 U10403 ( .A1(n9603), .A2(n9602), .ZN(n9631) );
  AOI22_X1 U10404 ( .A1(n9605), .A2(n7472), .B1(n9604), .B2(n10466), .ZN(n9615) );
  NOR2_X1 U10405 ( .A1(n9606), .A2(n10281), .ZN(n9608) );
  OAI22_X1 U10406 ( .A1(n9636), .A2(n7816), .B1(n10358), .B2(n9642), .ZN(n9607) );
  NOR2_X1 U10407 ( .A1(n9608), .A2(n9607), .ZN(n9610) );
  OAI211_X1 U10408 ( .C1(n9649), .C2(data_addr_o_9_), .A(n9610), .B(n9609), 
        .ZN(n9611) );
  INV_X1 U10409 ( .A(n9611), .ZN(n9613) );
  AND4_X1 U10410 ( .A1(n9615), .A2(n9614), .A3(n9613), .A4(n9612), .ZN(n9623)
         );
  AOI22_X1 U10411 ( .A1(n9617), .A2(n9941), .B1(n9616), .B2(n11334), .ZN(n9622) );
  XNOR2_X1 U10412 ( .A(n9618), .B(n11320), .ZN(n9621) );
  XNOR2_X1 U10413 ( .A(n9619), .B(n10635), .ZN(n9620) );
  NAND4_X1 U10414 ( .A1(n9623), .A2(n9622), .A3(n9621), .A4(n9620), .ZN(n9629)
         );
  XNOR2_X1 U10415 ( .A(n9624), .B(n11313), .ZN(n9627) );
  XNOR2_X1 U10416 ( .A(n9625), .B(n11312), .ZN(n9626) );
  NAND2_X1 U10417 ( .A1(n9627), .A2(n9626), .ZN(n9628) );
  NOR2_X1 U10418 ( .A1(n9629), .A2(n9628), .ZN(n9630) );
  AND2_X1 U10419 ( .A1(n9631), .A2(n9630), .ZN(n11878) );
  XNOR2_X1 U10420 ( .A(n9632), .B(n11303), .ZN(n11937) );
  XNOR2_X1 U10421 ( .A(n11883), .B(n10335), .ZN(n9633) );
  NAND4_X1 U10422 ( .A1(n11937), .A2(n9633), .A3(n11887), .A4(n11879), .ZN(
        n9656) );
  XNOR2_X1 U10423 ( .A(n9635), .B(n9634), .ZN(n9655) );
  NAND2_X1 U10424 ( .A1(n10493), .A2(n9636), .ZN(n11913) );
  AOI21_X1 U10425 ( .B1(n11259), .B2(n9470), .A(n9638), .ZN(n9640) );
  NAND2_X1 U10426 ( .A1(data_addr_o_4_), .A2(n9639), .ZN(n11906) );
  NAND4_X1 U10427 ( .A1(n11913), .A2(n9640), .A3(n11906), .A4(n11908), .ZN(
        n9641) );
  NOR2_X1 U10428 ( .A1(n11915), .A2(n9641), .ZN(n9651) );
  NAND2_X1 U10429 ( .A1(data_addr_o_6_), .A2(n9642), .ZN(n11900) );
  NAND2_X1 U10430 ( .A1(data_addr_o_5_), .A2(n9647), .ZN(n11899) );
  NAND2_X1 U10431 ( .A1(n11900), .A2(n11899), .ZN(n9648) );
  OAI22_X1 U10432 ( .A1(n10130), .A2(n9472), .B1(n11259), .B2(n9470), .ZN(
        n9644) );
  INV_X1 U10433 ( .A(n9644), .ZN(n9645) );
  OAI211_X1 U10434 ( .C1(n11255), .C2(n9647), .A(n9646), .B(n9645), .ZN(n11905) );
  NOR2_X1 U10435 ( .A1(n9648), .A2(n11905), .ZN(n9650) );
  NAND2_X1 U10436 ( .A1(data_addr_o_9_), .A2(n9649), .ZN(n11896) );
  NAND4_X1 U10437 ( .A1(n11928), .A2(n9651), .A3(n9650), .A4(n11896), .ZN(
        n9652) );
  NOR2_X1 U10438 ( .A1(n9652), .A2(n11922), .ZN(n9653) );
  NAND4_X1 U10439 ( .A1(n11888), .A2(n9653), .A3(n11893), .A4(n11933), .ZN(
        n9654) );
  NOR3_X1 U10440 ( .A1(n9656), .A2(n9655), .A3(n9654), .ZN(n9657) );
  NAND2_X1 U10441 ( .A1(n11878), .A2(n9657), .ZN(n9660) );
  MUX2_X1 U10442 ( .A(pmp_cfg_i[32]), .B(pmp_cfg_i[33]), .S(n11019), .Z(n9659)
         );
  NAND2_X1 U10443 ( .A1(n9658), .A2(n9659), .ZN(n11927) );
  AOI21_X1 U10444 ( .B1(n9661), .B2(n9660), .A(n11927), .ZN(n9999) );
  NOR2_X1 U10445 ( .A1(pmp_addr_i[428]), .A2(n6154), .ZN(n9662) );
  NOR2_X1 U10446 ( .A1(pmp_addr_i[429]), .A2(n10338), .ZN(n9705) );
  NOR2_X1 U10447 ( .A1(n9662), .A2(n9705), .ZN(n9664) );
  NOR2_X1 U10448 ( .A1(pmp_addr_i[430]), .A2(n10047), .ZN(n9663) );
  NOR2_X1 U10449 ( .A1(pmp_addr_i[431]), .A2(n7995), .ZN(n9708) );
  NOR2_X1 U10450 ( .A1(n9663), .A2(n9708), .ZN(n9711) );
  NAND2_X1 U10451 ( .A1(n9664), .A2(n9711), .ZN(n9713) );
  NOR2_X1 U10452 ( .A1(pmp_addr_i[424]), .A2(n6141), .ZN(n9665) );
  NOR2_X1 U10453 ( .A1(pmp_addr_i[425]), .A2(n9508), .ZN(n9696) );
  NOR2_X1 U10454 ( .A1(n9665), .A2(n9696), .ZN(n9667) );
  NOR2_X1 U10455 ( .A1(pmp_addr_i[426]), .A2(n10005), .ZN(n9666) );
  NOR2_X1 U10456 ( .A1(pmp_addr_i[427]), .A2(n10342), .ZN(n9699) );
  NOR2_X1 U10457 ( .A1(n9666), .A2(n9699), .ZN(n9702) );
  NAND2_X1 U10458 ( .A1(n9667), .A2(n9702), .ZN(n9668) );
  NOR2_X1 U10459 ( .A1(n9713), .A2(n9668), .ZN(n9717) );
  NOR2_X1 U10460 ( .A1(pmp_addr_i[418]), .A2(n6123), .ZN(n9669) );
  NOR2_X1 U10461 ( .A1(pmp_addr_i[419]), .A2(n10346), .ZN(n9675) );
  NOR2_X1 U10462 ( .A1(n9669), .A2(n9675), .ZN(n9678) );
  NOR2_X1 U10463 ( .A1(pmp_addr_i[417]), .A2(n9350), .ZN(n9672) );
  NAND2_X1 U10464 ( .A1(pmp_addr_i[416]), .A2(n10651), .ZN(n9671) );
  NAND2_X1 U10465 ( .A1(pmp_addr_i[417]), .A2(n9350), .ZN(n9670) );
  OAI21_X1 U10466 ( .B1(n9672), .B2(n9671), .A(n9670), .ZN(n9677) );
  NAND2_X1 U10467 ( .A1(pmp_addr_i[418]), .A2(n6123), .ZN(n9674) );
  NAND2_X1 U10468 ( .A1(pmp_addr_i[419]), .A2(n6127), .ZN(n9673) );
  OAI21_X1 U10469 ( .B1(n9675), .B2(n9674), .A(n9673), .ZN(n9676) );
  AOI21_X1 U10470 ( .B1(n9678), .B2(n9677), .A(n9676), .ZN(n9693) );
  NOR2_X1 U10471 ( .A1(pmp_addr_i[420]), .A2(n10362), .ZN(n9679) );
  NOR2_X1 U10472 ( .A1(pmp_addr_i[421]), .A2(n6400), .ZN(n9684) );
  NOR2_X1 U10473 ( .A1(n9679), .A2(n9684), .ZN(n9681) );
  NOR2_X1 U10474 ( .A1(pmp_addr_i[422]), .A2(n8735), .ZN(n9680) );
  NOR2_X1 U10475 ( .A1(pmp_addr_i[423]), .A2(n6140), .ZN(n9687) );
  NOR2_X1 U10476 ( .A1(n9680), .A2(n9687), .ZN(n9690) );
  NAND2_X1 U10477 ( .A1(n9681), .A2(n9690), .ZN(n9692) );
  NAND2_X1 U10478 ( .A1(pmp_addr_i[420]), .A2(n10362), .ZN(n9683) );
  NAND2_X1 U10479 ( .A1(pmp_addr_i[421]), .A2(n6400), .ZN(n9682) );
  OAI21_X1 U10480 ( .B1(n9684), .B2(n9683), .A(n9682), .ZN(n9689) );
  NAND2_X1 U10481 ( .A1(pmp_addr_i[422]), .A2(n8735), .ZN(n9686) );
  NAND2_X1 U10482 ( .A1(pmp_addr_i[423]), .A2(n6140), .ZN(n9685) );
  OAI21_X1 U10483 ( .B1(n9687), .B2(n9686), .A(n9685), .ZN(n9688) );
  AOI21_X1 U10484 ( .B1(n9690), .B2(n9689), .A(n9688), .ZN(n9691) );
  OAI21_X1 U10485 ( .B1(n9693), .B2(n9692), .A(n9691), .ZN(n9716) );
  NAND2_X1 U10486 ( .A1(pmp_addr_i[424]), .A2(n7964), .ZN(n9695) );
  NAND2_X1 U10487 ( .A1(pmp_addr_i[425]), .A2(n10711), .ZN(n9694) );
  OAI21_X1 U10488 ( .B1(n9696), .B2(n9695), .A(n9694), .ZN(n9701) );
  NAND2_X1 U10489 ( .A1(pmp_addr_i[426]), .A2(n10005), .ZN(n9698) );
  NAND2_X1 U10490 ( .A1(pmp_addr_i[427]), .A2(n10342), .ZN(n9697) );
  OAI21_X1 U10491 ( .B1(n9699), .B2(n9698), .A(n9697), .ZN(n9700) );
  AOI21_X1 U10492 ( .B1(n9702), .B2(n9701), .A(n9700), .ZN(n9714) );
  NAND2_X1 U10493 ( .A1(pmp_addr_i[428]), .A2(n11334), .ZN(n9704) );
  NAND2_X1 U10494 ( .A1(pmp_addr_i[429]), .A2(n10338), .ZN(n9703) );
  OAI21_X1 U10495 ( .B1(n9705), .B2(n9704), .A(n9703), .ZN(n9710) );
  NAND2_X1 U10496 ( .A1(pmp_addr_i[430]), .A2(n10047), .ZN(n9707) );
  NAND2_X1 U10497 ( .A1(pmp_addr_i[431]), .A2(n8444), .ZN(n9706) );
  OAI21_X1 U10498 ( .B1(n9708), .B2(n9707), .A(n9706), .ZN(n9709) );
  AOI21_X1 U10499 ( .B1(n9711), .B2(n9710), .A(n9709), .ZN(n9712) );
  OAI21_X1 U10500 ( .B1(n9714), .B2(n9713), .A(n9712), .ZN(n9715) );
  AOI21_X1 U10501 ( .B1(n9717), .B2(n9716), .A(n9715), .ZN(n9775) );
  NOR2_X1 U10502 ( .A1(pmp_addr_i[432]), .A2(n10403), .ZN(n9718) );
  NOR2_X1 U10503 ( .A1(pmp_addr_i[433]), .A2(n9414), .ZN(n9733) );
  NOR2_X1 U10504 ( .A1(n9718), .A2(n9733), .ZN(n9720) );
  NOR2_X1 U10505 ( .A1(pmp_addr_i[434]), .A2(n10754), .ZN(n9719) );
  NOR2_X1 U10506 ( .A1(pmp_addr_i[435]), .A2(n9418), .ZN(n9736) );
  NOR2_X1 U10507 ( .A1(n9719), .A2(n9736), .ZN(n9739) );
  NAND2_X1 U10508 ( .A1(n9720), .A2(n9739), .ZN(n9724) );
  NOR2_X1 U10509 ( .A1(pmp_addr_i[436]), .A2(n9156), .ZN(n9721) );
  NOR2_X1 U10510 ( .A1(pmp_addr_i[437]), .A2(n10064), .ZN(n9742) );
  NOR2_X1 U10511 ( .A1(n9721), .A2(n9742), .ZN(n9723) );
  NOR2_X1 U10512 ( .A1(pmp_addr_i[438]), .A2(n10428), .ZN(n9722) );
  NOR2_X1 U10513 ( .A1(pmp_addr_i[439]), .A2(n6462), .ZN(n9745) );
  NOR2_X1 U10514 ( .A1(n9722), .A2(n9745), .ZN(n9748) );
  NAND2_X1 U10515 ( .A1(n9723), .A2(n9748), .ZN(n9750) );
  NOR2_X1 U10516 ( .A1(n9724), .A2(n9750), .ZN(n9730) );
  NOR2_X1 U10517 ( .A1(pmp_addr_i[440]), .A2(n10439), .ZN(n9725) );
  INV_X1 U10518 ( .A(n10616), .ZN(n10096) );
  NOR2_X1 U10519 ( .A1(pmp_addr_i[441]), .A2(n10096), .ZN(n9754) );
  NOR2_X1 U10520 ( .A1(n9725), .A2(n9754), .ZN(n9727) );
  NOR2_X1 U10521 ( .A1(pmp_addr_i[443]), .A2(n6216), .ZN(n9757) );
  NOR2_X1 U10522 ( .A1(pmp_addr_i[442]), .A2(n8807), .ZN(n9726) );
  NOR2_X1 U10523 ( .A1(n9757), .A2(n9726), .ZN(n9760) );
  NAND2_X1 U10524 ( .A1(n9727), .A2(n9760), .ZN(n9729) );
  NOR2_X1 U10525 ( .A1(pmp_addr_i[445]), .A2(data_addr_o_31__BAR), .ZN(n9763)
         );
  NOR2_X1 U10526 ( .A1(pmp_addr_i[444]), .A2(n8814), .ZN(n9728) );
  OR2_X1 U10527 ( .A1(n9763), .A2(n9728), .ZN(n9768) );
  NOR2_X1 U10528 ( .A1(n9729), .A2(n9768), .ZN(n9771) );
  NAND2_X1 U10529 ( .A1(n9730), .A2(n9771), .ZN(n9774) );
  NAND2_X1 U10530 ( .A1(pmp_addr_i[432]), .A2(n12184), .ZN(n9732) );
  NAND2_X1 U10531 ( .A1(pmp_addr_i[433]), .A2(n10414), .ZN(n9731) );
  OAI21_X1 U10532 ( .B1(n9733), .B2(n9732), .A(n9731), .ZN(n9738) );
  NAND2_X1 U10533 ( .A1(pmp_addr_i[434]), .A2(n6188), .ZN(n9735) );
  NAND2_X1 U10534 ( .A1(pmp_addr_i[435]), .A2(n9418), .ZN(n9734) );
  OAI21_X1 U10535 ( .B1(n9736), .B2(n9735), .A(n9734), .ZN(n9737) );
  AOI21_X1 U10536 ( .B1(n9739), .B2(n9738), .A(n9737), .ZN(n9751) );
  NAND2_X1 U10537 ( .A1(pmp_addr_i[436]), .A2(n9156), .ZN(n9741) );
  NAND2_X1 U10538 ( .A1(pmp_addr_i[437]), .A2(n10064), .ZN(n9740) );
  OAI21_X1 U10539 ( .B1(n9742), .B2(n9741), .A(n9740), .ZN(n9747) );
  NAND2_X1 U10540 ( .A1(pmp_addr_i[438]), .A2(n10428), .ZN(n9744) );
  NAND2_X1 U10541 ( .A1(pmp_addr_i[439]), .A2(n6462), .ZN(n9743) );
  OAI21_X1 U10542 ( .B1(n9745), .B2(n9744), .A(n9743), .ZN(n9746) );
  AOI21_X1 U10543 ( .B1(n9748), .B2(n9747), .A(n9746), .ZN(n9749) );
  OAI21_X1 U10544 ( .B1(n9751), .B2(n9750), .A(n9749), .ZN(n9772) );
  NAND2_X1 U10545 ( .A1(pmp_addr_i[440]), .A2(n10439), .ZN(n9753) );
  NAND2_X1 U10546 ( .A1(pmp_addr_i[441]), .A2(n10096), .ZN(n9752) );
  OAI21_X1 U10547 ( .B1(n9754), .B2(n9753), .A(n9752), .ZN(n9759) );
  NAND2_X1 U10548 ( .A1(pmp_addr_i[442]), .A2(n10443), .ZN(n9756) );
  NAND2_X1 U10549 ( .A1(pmp_addr_i[443]), .A2(n10100), .ZN(n9755) );
  OAI21_X1 U10550 ( .B1(n9757), .B2(n9756), .A(n9755), .ZN(n9758) );
  AOI21_X1 U10551 ( .B1(n9760), .B2(n9759), .A(n9758), .ZN(n9769) );
  NAND2_X1 U10552 ( .A1(pmp_addr_i[444]), .A2(n8814), .ZN(n9762) );
  NAND2_X1 U10553 ( .A1(pmp_addr_i[445]), .A2(n10107), .ZN(n9761) );
  OAI21_X1 U10554 ( .B1(n9763), .B2(n9762), .A(n9761), .ZN(n9766) );
  INV_X1 U10555 ( .A(n9764), .ZN(n9765) );
  NOR2_X1 U10556 ( .A1(n9766), .A2(n9765), .ZN(n9767) );
  OAI21_X1 U10557 ( .B1(n9769), .B2(n9768), .A(n9767), .ZN(n9770) );
  AOI21_X1 U10558 ( .B1(n9772), .B2(n9771), .A(n9770), .ZN(n9773) );
  OAI21_X1 U10559 ( .B1(n9775), .B2(n9774), .A(n9773), .ZN(n9913) );
  NAND2_X1 U10560 ( .A1(n9842), .A2(n7995), .ZN(n9952) );
  INV_X1 U10561 ( .A(n9952), .ZN(n9776) );
  INV_X1 U10562 ( .A(n9939), .ZN(n9843) );
  NOR2_X1 U10563 ( .A1(n9843), .A2(n10857), .ZN(n9845) );
  NOR2_X1 U10564 ( .A1(n9776), .A2(n9845), .ZN(n9778) );
  INV_X1 U10565 ( .A(n9934), .ZN(n9847) );
  NOR2_X1 U10566 ( .A1(n9847), .A2(n9846), .ZN(n9777) );
  NOR2_X1 U10567 ( .A1(n4529), .A2(n10887), .ZN(n9850) );
  NOR2_X1 U10568 ( .A1(n9777), .A2(n9850), .ZN(n9853) );
  NAND2_X1 U10569 ( .A1(n9778), .A2(n9853), .ZN(n9782) );
  INV_X1 U10570 ( .A(n9914), .ZN(n9854) );
  NOR2_X1 U10571 ( .A1(n9854), .A2(n10891), .ZN(n9779) );
  INV_X1 U10572 ( .A(n9916), .ZN(n9855) );
  NOR2_X1 U10573 ( .A1(n9855), .A2(n9529), .ZN(n9858) );
  NOR2_X1 U10574 ( .A1(n9779), .A2(n9858), .ZN(n9781) );
  INV_X1 U10575 ( .A(n9917), .ZN(n9859) );
  NOR2_X1 U10576 ( .A1(n9859), .A2(data_addr_o_23_), .ZN(n9780) );
  NOR2_X1 U10577 ( .A1(n9860), .A2(n10899), .ZN(n9863) );
  NOR2_X1 U10578 ( .A1(n9780), .A2(n9863), .ZN(n9866) );
  NOR2_X1 U10579 ( .A1(n9782), .A2(n9868), .ZN(n9872) );
  NOR2_X1 U10580 ( .A1(n10129), .A2(n9973), .ZN(n9786) );
  NOR2_X1 U10581 ( .A1(n10818), .A2(n9967), .ZN(n9785) );
  NAND2_X1 U10582 ( .A1(n10818), .A2(n9967), .ZN(n11976) );
  OAI21_X1 U10583 ( .B1(n9786), .B2(n9785), .A(n11976), .ZN(n9789) );
  NAND2_X1 U10584 ( .A1(n12058), .A2(n9787), .ZN(n9970) );
  AND2_X1 U10585 ( .A1(n10135), .A2(n9974), .ZN(n9788) );
  AOI21_X1 U10586 ( .B1(n9789), .B2(n9970), .A(n9788), .ZN(n9797) );
  OR2_X1 U10587 ( .A1(data_addr_o_5_), .A2(n9971), .ZN(n9791) );
  OR2_X1 U10588 ( .A1(n10358), .A2(n3554), .ZN(n9794) );
  NAND2_X1 U10589 ( .A1(n9791), .A2(n9794), .ZN(n9796) );
  AND2_X1 U10590 ( .A1(n10486), .A2(n9971), .ZN(n9793) );
  AND2_X1 U10591 ( .A1(n10358), .A2(n3554), .ZN(n9792) );
  AOI21_X1 U10592 ( .B1(n9794), .B2(n9793), .A(n9792), .ZN(n9795) );
  OAI21_X1 U10593 ( .B1(n9797), .B2(n9796), .A(n9795), .ZN(n9817) );
  OR2_X1 U10594 ( .A1(n9805), .A2(n9979), .ZN(n9808) );
  OR2_X1 U10595 ( .A1(n7816), .A2(n4476), .ZN(n9800) );
  NAND2_X1 U10596 ( .A1(n9808), .A2(n9800), .ZN(n9804) );
  OR2_X1 U10597 ( .A1(data_addr_o_9_), .A2(n9978), .ZN(n9803) );
  OR2_X1 U10598 ( .A1(data_addr_o_10_), .A2(n9966), .ZN(n9811) );
  NAND2_X1 U10599 ( .A1(n9803), .A2(n9811), .ZN(n9813) );
  NOR2_X1 U10600 ( .A1(n9804), .A2(n9813), .ZN(n9816) );
  AND2_X1 U10601 ( .A1(n7816), .A2(n4476), .ZN(n9807) );
  AND2_X1 U10602 ( .A1(n9805), .A2(n9979), .ZN(n9806) );
  AOI21_X1 U10603 ( .B1(n9808), .B2(n9807), .A(n9806), .ZN(n9814) );
  AND2_X1 U10604 ( .A1(data_addr_o_9_), .A2(n9978), .ZN(n9810) );
  AND2_X1 U10605 ( .A1(data_addr_o_10_), .A2(n9966), .ZN(n9809) );
  AOI21_X1 U10606 ( .B1(n9811), .B2(n9810), .A(n9809), .ZN(n9812) );
  OAI21_X1 U10607 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(n9815) );
  AOI21_X1 U10608 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n9841) );
  NOR2_X1 U10609 ( .A1(n11014), .A2(n9986), .ZN(n9835) );
  NOR2_X1 U10610 ( .A1(n10657), .A2(n4497), .ZN(n9818) );
  NOR2_X1 U10611 ( .A1(n9835), .A2(n9818), .ZN(n9838) );
  OR2_X1 U10612 ( .A1(data_addr_o_11_), .A2(n9965), .ZN(n9820) );
  OR2_X1 U10613 ( .A1(n10499), .A2(n9983), .ZN(n9827) );
  NAND2_X1 U10614 ( .A1(n9820), .A2(n9827), .ZN(n9823) );
  OR2_X1 U10615 ( .A1(data_addr_o_13_), .A2(n9982), .ZN(n9822) );
  OR2_X1 U10616 ( .A1(data_addr_o_14_), .A2(n9988), .ZN(n9830) );
  NAND2_X1 U10617 ( .A1(n9822), .A2(n9830), .ZN(n9832) );
  NOR2_X1 U10618 ( .A1(n9823), .A2(n9832), .ZN(n9824) );
  NAND2_X1 U10619 ( .A1(n9838), .A2(n9824), .ZN(n9840) );
  AND2_X1 U10620 ( .A1(data_addr_o_11_), .A2(n9965), .ZN(n9826) );
  AND2_X1 U10621 ( .A1(n10499), .A2(n9983), .ZN(n9825) );
  AOI21_X1 U10622 ( .B1(n9827), .B2(n9826), .A(n9825), .ZN(n9833) );
  AND2_X1 U10623 ( .A1(data_addr_o_13_), .A2(n9982), .ZN(n9829) );
  AND2_X1 U10624 ( .A1(data_addr_o_14_), .A2(n9988), .ZN(n9828) );
  AOI21_X1 U10625 ( .B1(n9830), .B2(n9829), .A(n9828), .ZN(n9831) );
  OAI21_X1 U10626 ( .B1(n9833), .B2(n9832), .A(n9831), .ZN(n9837) );
  NAND2_X1 U10627 ( .A1(n10657), .A2(n4497), .ZN(n11991) );
  NAND2_X1 U10628 ( .A1(n11014), .A2(n9986), .ZN(n9834) );
  OAI21_X1 U10629 ( .B1(n9835), .B2(n11991), .A(n9834), .ZN(n9836) );
  AOI21_X1 U10630 ( .B1(n9838), .B2(n9837), .A(n9836), .ZN(n9839) );
  OAI21_X1 U10631 ( .B1(n9841), .B2(n9840), .A(n9839), .ZN(n9871) );
  OR2_X1 U10632 ( .A1(n9842), .A2(n7995), .ZN(n11946) );
  NAND2_X1 U10633 ( .A1(n9843), .A2(n10857), .ZN(n9844) );
  OAI21_X1 U10634 ( .B1(n9845), .B2(n11946), .A(n9844), .ZN(n9852) );
  NAND2_X1 U10635 ( .A1(n9847), .A2(n9846), .ZN(n9849) );
  NAND2_X1 U10636 ( .A1(n4529), .A2(n10887), .ZN(n9848) );
  OAI21_X1 U10637 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9851) );
  AOI21_X1 U10638 ( .B1(n9853), .B2(n9852), .A(n9851), .ZN(n9869) );
  NAND2_X1 U10639 ( .A1(n9854), .A2(n10891), .ZN(n9857) );
  NAND2_X1 U10640 ( .A1(n9855), .A2(n11313), .ZN(n9856) );
  OAI21_X1 U10641 ( .B1(n9858), .B2(n9857), .A(n9856), .ZN(n9865) );
  NAND2_X1 U10642 ( .A1(n9859), .A2(n10898), .ZN(n9862) );
  NAND2_X1 U10643 ( .A1(n9860), .A2(n10899), .ZN(n9861) );
  OAI21_X1 U10644 ( .B1(n9863), .B2(n9862), .A(n9861), .ZN(n9864) );
  AOI21_X1 U10645 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(n9867) );
  OAI21_X1 U10646 ( .B1(n9869), .B2(n9868), .A(n9867), .ZN(n9870) );
  AOI21_X1 U10647 ( .B1(n9872), .B2(n9871), .A(n9870), .ZN(n9910) );
  INV_X1 U10648 ( .A(n9924), .ZN(n9881) );
  NOR2_X1 U10649 ( .A1(n9881), .A2(n10903), .ZN(n9873) );
  INV_X1 U10650 ( .A(n9925), .ZN(n9882) );
  NOR2_X1 U10651 ( .A1(n9882), .A2(n10904), .ZN(n9885) );
  NOR2_X1 U10652 ( .A1(n9873), .A2(n9885), .ZN(n9875) );
  INV_X1 U10653 ( .A(n9926), .ZN(n9887) );
  NOR2_X1 U10654 ( .A1(n9887), .A2(n9886), .ZN(n9874) );
  INV_X1 U10655 ( .A(n9927), .ZN(n9888) );
  NOR2_X1 U10656 ( .A1(n9888), .A2(n10635), .ZN(n9891) );
  NOR2_X1 U10657 ( .A1(n9874), .A2(n9891), .ZN(n9894) );
  NAND2_X1 U10658 ( .A1(n9875), .A2(n9894), .ZN(n9879) );
  INV_X1 U10659 ( .A(n9956), .ZN(n9895) );
  NOR2_X1 U10660 ( .A1(n9895), .A2(n9955), .ZN(n9876) );
  INV_X1 U10661 ( .A(n9957), .ZN(n9896) );
  NOR2_X1 U10662 ( .A1(n9896), .A2(n10919), .ZN(n9899) );
  NOR2_X1 U10663 ( .A1(n9876), .A2(n9899), .ZN(n9878) );
  NOR2_X1 U10664 ( .A1(n4567), .A2(n24), .ZN(n9877) );
  NOR2_X1 U10665 ( .A1(n9877), .A2(pmp_addr_i[414]), .ZN(n9903) );
  NAND2_X1 U10666 ( .A1(n9878), .A2(n9903), .ZN(n9905) );
  NOR2_X1 U10667 ( .A1(n9879), .A2(n9905), .ZN(n9880) );
  NAND2_X1 U10668 ( .A1(n9880), .A2(n4459), .ZN(n9909) );
  NAND2_X1 U10669 ( .A1(n9881), .A2(n10903), .ZN(n9884) );
  NAND2_X1 U10670 ( .A1(n9882), .A2(n10904), .ZN(n9883) );
  OAI21_X1 U10671 ( .B1(n9885), .B2(n9884), .A(n9883), .ZN(n9893) );
  NAND2_X1 U10672 ( .A1(n9887), .A2(n9886), .ZN(n9890) );
  NAND2_X1 U10673 ( .A1(n9888), .A2(n10914), .ZN(n9889) );
  OAI21_X1 U10674 ( .B1(n9891), .B2(n9890), .A(n9889), .ZN(n9892) );
  AOI21_X1 U10675 ( .B1(n9894), .B2(n9893), .A(n9892), .ZN(n9906) );
  NAND2_X1 U10676 ( .A1(n9895), .A2(n9955), .ZN(n9898) );
  NAND2_X1 U10677 ( .A1(n9896), .A2(n10919), .ZN(n9897) );
  OAI21_X1 U10678 ( .B1(n9899), .B2(n9898), .A(n9897), .ZN(n9902) );
  NAND2_X1 U10679 ( .A1(n4567), .A2(n24), .ZN(n9900) );
  NOR2_X1 U10680 ( .A1(n9900), .A2(pmp_addr_i[414]), .ZN(n9901) );
  AOI21_X1 U10681 ( .B1(n9903), .B2(n9902), .A(n9901), .ZN(n9904) );
  OAI21_X1 U10682 ( .B1(n9906), .B2(n9905), .A(n9904), .ZN(n9907) );
  NAND2_X1 U10683 ( .A1(n9907), .A2(n4459), .ZN(n9908) );
  OAI21_X1 U10684 ( .B1(n9910), .B2(n9909), .A(n9908), .ZN(n9912) );
  XNOR2_X1 U10685 ( .A(n9914), .B(n10202), .ZN(n9922) );
  XNOR2_X1 U10686 ( .A(n9916), .B(n9915), .ZN(n9921) );
  XNOR2_X1 U10687 ( .A(n9917), .B(n10898), .ZN(n9920) );
  XNOR2_X1 U10688 ( .A(n9918), .B(n10738), .ZN(n9919) );
  NAND4_X1 U10689 ( .A1(n9922), .A2(n9921), .A3(n9920), .A4(n9919), .ZN(n9933)
         );
  XNOR2_X1 U10690 ( .A(n9924), .B(n9923), .ZN(n9931) );
  XNOR2_X1 U10691 ( .A(n9925), .B(n10904), .ZN(n9930) );
  XNOR2_X1 U10692 ( .A(n9926), .B(n10746), .ZN(n9929) );
  XNOR2_X1 U10693 ( .A(n9927), .B(n10914), .ZN(n9928) );
  NAND4_X1 U10694 ( .A1(n9931), .A2(n9930), .A3(n9929), .A4(n9928), .ZN(n9932)
         );
  OR2_X1 U10695 ( .A1(n9933), .A2(n9932), .ZN(n9963) );
  XNOR2_X1 U10696 ( .A(n9934), .B(n9846), .ZN(n9938) );
  XNOR2_X1 U10697 ( .A(n9936), .B(n9935), .ZN(n9937) );
  AND2_X1 U10698 ( .A1(n9938), .A2(n9937), .ZN(n9961) );
  XNOR2_X1 U10699 ( .A(n9939), .B(n10297), .ZN(n9954) );
  AOI22_X1 U10700 ( .A1(n9942), .A2(n9941), .B1(n11334), .B2(n9940), .ZN(n9951) );
  OAI22_X1 U10701 ( .A1(n9966), .A2(n11343), .B1(data_addr_o_11_), .B2(n9965), 
        .ZN(n9945) );
  OAI22_X1 U10702 ( .A1(data_addr_o_9_), .A2(n9978), .B1(n10281), .B2(n9979), 
        .ZN(n9944) );
  OAI22_X1 U10703 ( .A1(n4476), .A2(n7816), .B1(n10358), .B2(n3554), .ZN(n9943) );
  NOR3_X1 U10704 ( .A1(n9945), .A2(n9944), .A3(n9943), .ZN(n9950) );
  AOI22_X1 U10705 ( .A1(n9948), .A2(n9947), .B1(n11006), .B2(n9946), .ZN(n9949) );
  NAND4_X1 U10706 ( .A1(n9952), .A2(n9951), .A3(n9950), .A4(n9949), .ZN(n9953)
         );
  NOR2_X1 U10707 ( .A1(n9954), .A2(n9953), .ZN(n9960) );
  XNOR2_X1 U10708 ( .A(n9956), .B(n9955), .ZN(n9959) );
  XNOR2_X1 U10709 ( .A(n9957), .B(n10919), .ZN(n9958) );
  NAND4_X1 U10710 ( .A1(n9961), .A2(n9960), .A3(n9959), .A4(n9958), .ZN(n9962)
         );
  NOR2_X1 U10711 ( .A1(n9963), .A2(n9962), .ZN(n11945) );
  XNOR2_X1 U10712 ( .A(n9964), .B(n12123), .ZN(n9993) );
  NAND2_X1 U10713 ( .A1(n8246), .A2(n9965), .ZN(n11986) );
  NAND2_X1 U10714 ( .A1(data_addr_o_10_), .A2(n9966), .ZN(n11974) );
  NAND2_X1 U10715 ( .A1(n11986), .A2(n11974), .ZN(n9977) );
  OAI22_X1 U10716 ( .A1(n10958), .A2(n9967), .B1(n10129), .B2(n9973), .ZN(
        n9968) );
  INV_X1 U10717 ( .A(n9968), .ZN(n9969) );
  OAI211_X1 U10718 ( .C1(n11255), .C2(n9971), .A(n9970), .B(n9969), .ZN(n11983) );
  NAND2_X1 U10719 ( .A1(n10655), .A2(n3554), .ZN(n11970) );
  AOI21_X1 U10720 ( .B1(n11259), .B2(n9973), .A(n9972), .ZN(n9975) );
  NAND2_X1 U10721 ( .A1(data_addr_o_4_), .A2(n9974), .ZN(n11982) );
  NAND4_X1 U10722 ( .A1(n11970), .A2(n9975), .A3(n11982), .A4(n11976), .ZN(
        n9976) );
  NOR3_X1 U10723 ( .A1(n9977), .A2(n11983), .A3(n9976), .ZN(n9985) );
  NAND2_X1 U10724 ( .A1(data_addr_o_9_), .A2(n9978), .ZN(n11987) );
  NAND2_X1 U10725 ( .A1(n10494), .A2(n9979), .ZN(n11971) );
  NAND2_X1 U10726 ( .A1(n11987), .A2(n11971), .ZN(n9981) );
  NAND2_X1 U10727 ( .A1(n10493), .A2(n4476), .ZN(n11955) );
  OAI21_X1 U10728 ( .B1(n11291), .B2(n9980), .A(n11955), .ZN(n11956) );
  NOR2_X1 U10729 ( .A1(n9981), .A2(n11956), .ZN(n9984) );
  NAND2_X1 U10730 ( .A1(n9982), .A2(data_addr_o_13_), .ZN(n11951) );
  NAND2_X1 U10731 ( .A1(n9983), .A2(data_addr_o_12_), .ZN(n11993) );
  NAND4_X1 U10732 ( .A1(n9985), .A2(n9984), .A3(n11951), .A4(n11993), .ZN(
        n9991) );
  XNOR2_X1 U10733 ( .A(n9987), .B(n9986), .ZN(n9990) );
  NAND2_X1 U10734 ( .A1(n9988), .A2(n9066), .ZN(n11961) );
  NAND2_X1 U10735 ( .A1(n11961), .A2(n11991), .ZN(n9989) );
  NOR3_X1 U10736 ( .A1(n9991), .A2(n9990), .A3(n9989), .ZN(n9992) );
  NAND4_X1 U10737 ( .A1(n11945), .A2(n9993), .A3(n9992), .A4(n11946), .ZN(
        n9996) );
  MUX2_X1 U10738 ( .A(pmp_cfg_i[104]), .B(pmp_cfg_i[105]), .S(n11019), .Z(
        n9995) );
  NAND2_X1 U10739 ( .A1(n9994), .A2(n9995), .ZN(n11998) );
  AOI21_X1 U10740 ( .B1(n9997), .B2(n9996), .A(n11998), .ZN(n9998) );
  NOR2_X1 U10741 ( .A1(n9999), .A2(n9998), .ZN(n11028) );
  NOR2_X1 U10742 ( .A1(pmp_addr_i[364]), .A2(n10000), .ZN(n10001) );
  NOR2_X1 U10743 ( .A1(pmp_addr_i[365]), .A2(n10338), .ZN(n10046) );
  NOR2_X1 U10744 ( .A1(n10001), .A2(n10046), .ZN(n10003) );
  NOR2_X1 U10746 ( .A1(pmp_addr_i[366]), .A2(n10047), .ZN(n10002) );
  NOR2_X1 U10747 ( .A1(pmp_addr_i[367]), .A2(n8757), .ZN(n10050) );
  NOR2_X1 U10748 ( .A1(n10002), .A2(n10050), .ZN(n10053) );
  NAND2_X1 U10749 ( .A1(n10003), .A2(n10053), .ZN(n10055) );
  NOR2_X1 U10750 ( .A1(pmp_addr_i[360]), .A2(n6141), .ZN(n10004) );
  NOR2_X1 U10751 ( .A1(pmp_addr_i[361]), .A2(n9508), .ZN(n10037) );
  NOR2_X1 U10752 ( .A1(n10004), .A2(n10037), .ZN(n10007) );
  NOR2_X1 U10753 ( .A1(pmp_addr_i[362]), .A2(n10005), .ZN(n10006) );
  NOR2_X1 U10754 ( .A1(pmp_addr_i[363]), .A2(n11006), .ZN(n10040) );
  NOR2_X1 U10755 ( .A1(n10006), .A2(n10040), .ZN(n10043) );
  NAND2_X1 U10756 ( .A1(n10007), .A2(n10043), .ZN(n10008) );
  NOR2_X1 U10757 ( .A1(n10055), .A2(n10008), .ZN(n10059) );
  NOR2_X1 U10758 ( .A1(pmp_addr_i[354]), .A2(n10351), .ZN(n10009) );
  NOR2_X1 U10759 ( .A1(pmp_addr_i[355]), .A2(n10346), .ZN(n10016) );
  NOR2_X1 U10760 ( .A1(n10009), .A2(n10016), .ZN(n10019) );
  NOR2_X1 U10761 ( .A1(pmp_addr_i[353]), .A2(n10010), .ZN(n10013) );
  NAND2_X1 U10762 ( .A1(pmp_addr_i[352]), .A2(n10651), .ZN(n10012) );
  NAND2_X1 U10763 ( .A1(pmp_addr_i[353]), .A2(n10010), .ZN(n10011) );
  OAI21_X1 U10764 ( .B1(n10013), .B2(n10012), .A(n10011), .ZN(n10018) );
  NAND2_X1 U10765 ( .A1(pmp_addr_i[354]), .A2(n8406), .ZN(n10015) );
  NAND2_X1 U10766 ( .A1(pmp_addr_i[355]), .A2(n6127), .ZN(n10014) );
  OAI21_X1 U10767 ( .B1(n10016), .B2(n10015), .A(n10014), .ZN(n10017) );
  AOI21_X1 U10768 ( .B1(n10019), .B2(n10018), .A(n10017), .ZN(n10034) );
  NOR2_X1 U10769 ( .A1(pmp_addr_i[356]), .A2(n9363), .ZN(n10020) );
  NOR2_X1 U10770 ( .A1(pmp_addr_i[357]), .A2(n6400), .ZN(n10025) );
  NOR2_X1 U10771 ( .A1(n10020), .A2(n10025), .ZN(n10022) );
  NOR2_X1 U10772 ( .A1(pmp_addr_i[358]), .A2(n29), .ZN(n10021) );
  NOR2_X1 U10773 ( .A1(pmp_addr_i[359]), .A2(n6140), .ZN(n10028) );
  NOR2_X1 U10774 ( .A1(n10021), .A2(n10028), .ZN(n10031) );
  NAND2_X1 U10775 ( .A1(n10022), .A2(n10031), .ZN(n10033) );
  NAND2_X1 U10776 ( .A1(pmp_addr_i[356]), .A2(n9363), .ZN(n10024) );
  NAND2_X1 U10777 ( .A1(pmp_addr_i[357]), .A2(n7152), .ZN(n10023) );
  OAI21_X1 U10778 ( .B1(n10025), .B2(n10024), .A(n10023), .ZN(n10030) );
  NAND2_X1 U10779 ( .A1(pmp_addr_i[358]), .A2(n8735), .ZN(n10027) );
  NAND2_X1 U10780 ( .A1(pmp_addr_i[359]), .A2(n10501), .ZN(n10026) );
  OAI21_X1 U10781 ( .B1(n10028), .B2(n10027), .A(n10026), .ZN(n10029) );
  AOI21_X1 U10782 ( .B1(n10031), .B2(n10030), .A(n10029), .ZN(n10032) );
  OAI21_X1 U10783 ( .B1(n10034), .B2(n10033), .A(n10032), .ZN(n10058) );
  NAND2_X1 U10784 ( .A1(pmp_addr_i[360]), .A2(n10701), .ZN(n10036) );
  NAND2_X1 U10785 ( .A1(pmp_addr_i[361]), .A2(n9508), .ZN(n10035) );
  OAI21_X1 U10786 ( .B1(n10037), .B2(n10036), .A(n10035), .ZN(n10042) );
  NAND2_X1 U10787 ( .A1(pmp_addr_i[362]), .A2(n7976), .ZN(n10039) );
  NAND2_X1 U10788 ( .A1(pmp_addr_i[363]), .A2(n11006), .ZN(n10038) );
  OAI21_X1 U10789 ( .B1(n10040), .B2(n10039), .A(n10038), .ZN(n10041) );
  AOI21_X1 U10790 ( .B1(n10043), .B2(n10042), .A(n10041), .ZN(n10056) );
  NAND2_X1 U10791 ( .A1(pmp_addr_i[364]), .A2(n10000), .ZN(n10045) );
  NAND2_X1 U10792 ( .A1(pmp_addr_i[365]), .A2(n10338), .ZN(n10044) );
  OAI21_X1 U10793 ( .B1(n10046), .B2(n10045), .A(n10044), .ZN(n10052) );
  NAND2_X1 U10794 ( .A1(pmp_addr_i[366]), .A2(n10047), .ZN(n10049) );
  NAND2_X1 U10795 ( .A1(pmp_addr_i[367]), .A2(n8757), .ZN(n10048) );
  OAI21_X1 U10796 ( .B1(n10050), .B2(n10049), .A(n10048), .ZN(n10051) );
  AOI21_X1 U10797 ( .B1(n10053), .B2(n10052), .A(n10051), .ZN(n10054) );
  OAI21_X1 U10798 ( .B1(n10056), .B2(n10055), .A(n10054), .ZN(n10057) );
  AOI21_X1 U10799 ( .B1(n10059), .B2(n10058), .A(n10057), .ZN(n10121) );
  NOR2_X1 U10800 ( .A1(pmp_addr_i[368]), .A2(n10060), .ZN(n10061) );
  NOR2_X1 U10801 ( .A1(pmp_addr_i[369]), .A2(n10753), .ZN(n10077) );
  NOR2_X1 U10802 ( .A1(n10061), .A2(n10077), .ZN(n10063) );
  NOR2_X1 U10803 ( .A1(pmp_addr_i[370]), .A2(n6188), .ZN(n10062) );
  NOR2_X1 U10804 ( .A1(pmp_addr_i[371]), .A2(n6192), .ZN(n10080) );
  NOR2_X1 U10805 ( .A1(n10062), .A2(n10080), .ZN(n10083) );
  NAND2_X1 U10806 ( .A1(n10063), .A2(n10083), .ZN(n10068) );
  NOR2_X1 U10807 ( .A1(pmp_addr_i[372]), .A2(n9425), .ZN(n10065) );
  NOR2_X1 U10808 ( .A1(pmp_addr_i[373]), .A2(n10064), .ZN(n10086) );
  NOR2_X1 U10809 ( .A1(n10065), .A2(n10086), .ZN(n10067) );
  NOR2_X1 U10810 ( .A1(pmp_addr_i[374]), .A2(n9163), .ZN(n10066) );
  NOR2_X1 U10811 ( .A1(pmp_addr_i[375]), .A2(n10768), .ZN(n10089) );
  NOR2_X1 U10812 ( .A1(n10066), .A2(n10089), .ZN(n10092) );
  NAND2_X1 U10813 ( .A1(n10067), .A2(n10092), .ZN(n10094) );
  NOR2_X1 U10814 ( .A1(n10068), .A2(n10094), .ZN(n10074) );
  NOR2_X1 U10815 ( .A1(pmp_addr_i[376]), .A2(n6202), .ZN(n10069) );
  NOR2_X1 U10816 ( .A1(pmp_addr_i[377]), .A2(n10096), .ZN(n10099) );
  NOR2_X1 U10817 ( .A1(n10069), .A2(n10099), .ZN(n10071) );
  NOR2_X1 U10818 ( .A1(pmp_addr_i[379]), .A2(n10100), .ZN(n10103) );
  NOR2_X1 U10819 ( .A1(pmp_addr_i[378]), .A2(n8807), .ZN(n10070) );
  NOR2_X1 U10820 ( .A1(n10103), .A2(n10070), .ZN(n10106) );
  NAND2_X1 U10821 ( .A1(n10071), .A2(n10106), .ZN(n10073) );
  NOR2_X1 U10822 ( .A1(pmp_addr_i[381]), .A2(data_addr_o_31__BAR), .ZN(n10110)
         );
  NOR2_X1 U10823 ( .A1(pmp_addr_i[380]), .A2(n8814), .ZN(n10072) );
  OR2_X1 U10824 ( .A1(n10110), .A2(n10072), .ZN(n10114) );
  NOR2_X1 U10825 ( .A1(n10073), .A2(n10114), .ZN(n10117) );
  NAND2_X1 U10826 ( .A1(n10074), .A2(n10117), .ZN(n10120) );
  NAND2_X1 U10827 ( .A1(pmp_addr_i[368]), .A2(n12184), .ZN(n10076) );
  NAND2_X1 U10828 ( .A1(pmp_addr_i[369]), .A2(n9414), .ZN(n10075) );
  OAI21_X1 U10829 ( .B1(n10077), .B2(n10076), .A(n10075), .ZN(n10082) );
  NAND2_X1 U10830 ( .A1(pmp_addr_i[370]), .A2(n10754), .ZN(n10079) );
  NAND2_X1 U10831 ( .A1(pmp_addr_i[371]), .A2(n6192), .ZN(n10078) );
  OAI21_X1 U10832 ( .B1(n10080), .B2(n10079), .A(n10078), .ZN(n10081) );
  AOI21_X1 U10833 ( .B1(n10083), .B2(n10082), .A(n10081), .ZN(n10095) );
  NAND2_X1 U10834 ( .A1(pmp_addr_i[372]), .A2(n9425), .ZN(n10085) );
  NAND2_X1 U10835 ( .A1(pmp_addr_i[373]), .A2(n10064), .ZN(n10084) );
  OAI21_X1 U10836 ( .B1(n10086), .B2(n10085), .A(n10084), .ZN(n10091) );
  NAND2_X1 U10837 ( .A1(pmp_addr_i[374]), .A2(n9163), .ZN(n10088) );
  NAND2_X1 U10838 ( .A1(pmp_addr_i[375]), .A2(n6462), .ZN(n10087) );
  OAI21_X1 U10839 ( .B1(n10089), .B2(n10088), .A(n10087), .ZN(n10090) );
  AOI21_X1 U10840 ( .B1(n10092), .B2(n10091), .A(n10090), .ZN(n10093) );
  OAI21_X1 U10841 ( .B1(n10095), .B2(n10094), .A(n10093), .ZN(n10118) );
  NAND2_X1 U10842 ( .A1(pmp_addr_i[376]), .A2(n6202), .ZN(n10098) );
  NAND2_X1 U10843 ( .A1(pmp_addr_i[377]), .A2(n10096), .ZN(n10097) );
  OAI21_X1 U10844 ( .B1(n10099), .B2(n10098), .A(n10097), .ZN(n10105) );
  NAND2_X1 U10845 ( .A1(pmp_addr_i[378]), .A2(n10778), .ZN(n10102) );
  NAND2_X1 U10846 ( .A1(pmp_addr_i[379]), .A2(n10100), .ZN(n10101) );
  OAI21_X1 U10847 ( .B1(n10103), .B2(n10102), .A(n10101), .ZN(n10104) );
  AOI21_X1 U10848 ( .B1(n10106), .B2(n10105), .A(n10104), .ZN(n10115) );
  NAND2_X1 U10849 ( .A1(pmp_addr_i[380]), .A2(n8814), .ZN(n10109) );
  NAND2_X1 U10850 ( .A1(pmp_addr_i[381]), .A2(n10107), .ZN(n10108) );
  OAI21_X1 U10851 ( .B1(n10110), .B2(n10109), .A(n10108), .ZN(n10112) );
  NOR2_X1 U10852 ( .A1(n10112), .A2(n1548), .ZN(n10113) );
  OAI21_X1 U10853 ( .B1(n10115), .B2(n10114), .A(n10113), .ZN(n10116) );
  AOI21_X1 U10854 ( .B1(n10118), .B2(n10117), .A(n10116), .ZN(n10119) );
  OAI21_X1 U10855 ( .B1(n10121), .B2(n10120), .A(n10119), .ZN(n10332) );
  NOR2_X1 U10856 ( .A1(n34), .A2(n10202), .ZN(n10122) );
  INV_X1 U10857 ( .A(n10270), .ZN(n10203) );
  NOR2_X1 U10858 ( .A1(n10203), .A2(n9915), .ZN(n10206) );
  NOR2_X1 U10859 ( .A1(n10122), .A2(n10206), .ZN(n10124) );
  INV_X1 U10860 ( .A(n10259), .ZN(n10208) );
  NOR2_X1 U10861 ( .A1(n10208), .A2(n10899), .ZN(n10211) );
  INV_X1 U10862 ( .A(n10279), .ZN(n10207) );
  NOR2_X1 U10863 ( .A1(n10207), .A2(n10898), .ZN(n10123) );
  NAND2_X1 U10864 ( .A1(n10124), .A2(n10214), .ZN(n10216) );
  INV_X1 U10865 ( .A(n10261), .ZN(n10194) );
  NOR2_X1 U10866 ( .A1(n10194), .A2(n10886), .ZN(n10125) );
  INV_X1 U10867 ( .A(n10296), .ZN(n10195) );
  NOR2_X1 U10868 ( .A1(n10195), .A2(n10887), .ZN(n10198) );
  NOR2_X1 U10869 ( .A1(n10125), .A2(n10198), .ZN(n10201) );
  INV_X1 U10870 ( .A(n10298), .ZN(n10191) );
  NOR2_X1 U10871 ( .A1(n10191), .A2(n10857), .ZN(n10193) );
  NOR2_X1 U10872 ( .A1(n5973), .A2(n6813), .ZN(n10126) );
  NOR2_X1 U10873 ( .A1(n10193), .A2(n10126), .ZN(n10127) );
  NAND2_X1 U10874 ( .A1(n10201), .A2(n10127), .ZN(n10128) );
  NOR2_X1 U10875 ( .A1(n10216), .A2(n10128), .ZN(n10220) );
  NOR2_X1 U10876 ( .A1(n10129), .A2(n6012), .ZN(n10133) );
  NOR2_X1 U10877 ( .A1(n10130), .A2(n10319), .ZN(n10132) );
  NAND2_X1 U10878 ( .A1(n10130), .A2(n10319), .ZN(n10131) );
  OAI21_X1 U10879 ( .B1(n10133), .B2(n10132), .A(n10131), .ZN(n10138) );
  OR2_X1 U10880 ( .A1(n10135), .A2(n12059), .ZN(n10137) );
  AND2_X1 U10881 ( .A1(n10135), .A2(n12059), .ZN(n10136) );
  AOI21_X1 U10882 ( .B1(n10138), .B2(n10137), .A(n10136), .ZN(n10144) );
  NAND2_X1 U10883 ( .A1(n11291), .A2(n10307), .ZN(n12030) );
  OR2_X1 U10884 ( .A1(n10655), .A2(n10306), .ZN(n10141) );
  NAND2_X1 U10885 ( .A1(n12030), .A2(n10141), .ZN(n10143) );
  AND2_X1 U10886 ( .A1(n10824), .A2(n6014), .ZN(n12043) );
  AND2_X1 U10887 ( .A1(n10655), .A2(n10306), .ZN(n10140) );
  AOI21_X1 U10888 ( .B1(n10141), .B2(n12043), .A(n10140), .ZN(n10142) );
  OAI21_X1 U10889 ( .B1(n10144), .B2(n10143), .A(n10142), .ZN(n10164) );
  OR2_X1 U10890 ( .A1(n10836), .A2(n10322), .ZN(n10154) );
  OR2_X1 U10891 ( .A1(n10493), .A2(n10309), .ZN(n10147) );
  NAND2_X1 U10892 ( .A1(n10154), .A2(n10147), .ZN(n10151) );
  OR2_X1 U10893 ( .A1(data_addr_o_9_), .A2(n10305), .ZN(n10150) );
  OR2_X1 U10894 ( .A1(data_addr_o_10_), .A2(n10317), .ZN(n10158) );
  NAND2_X1 U10895 ( .A1(n10150), .A2(n10158), .ZN(n10160) );
  NOR2_X1 U10896 ( .A1(n10151), .A2(n10160), .ZN(n10163) );
  AND2_X1 U10897 ( .A1(n7816), .A2(n10309), .ZN(n10153) );
  AND2_X1 U10898 ( .A1(n9805), .A2(n10322), .ZN(n10152) );
  AOI21_X1 U10899 ( .B1(n10154), .B2(n10153), .A(n10152), .ZN(n10161) );
  AND2_X1 U10900 ( .A1(data_addr_o_9_), .A2(n10305), .ZN(n10157) );
  AND2_X1 U10901 ( .A1(data_addr_o_10_), .A2(n10317), .ZN(n10156) );
  AOI21_X1 U10902 ( .B1(n10158), .B2(n10157), .A(n10156), .ZN(n10159) );
  OAI21_X1 U10903 ( .B1(n10161), .B2(n10160), .A(n10159), .ZN(n10162) );
  AOI21_X1 U10904 ( .B1(n10164), .B2(n10163), .A(n10162), .ZN(n10190) );
  NOR2_X1 U10905 ( .A1(n10335), .A2(n6003), .ZN(n10184) );
  NOR2_X1 U10906 ( .A1(data_addr_o_15_), .A2(n3010), .ZN(n10165) );
  NOR2_X1 U10907 ( .A1(n10184), .A2(n10165), .ZN(n10187) );
  OR2_X1 U10908 ( .A1(n10508), .A2(n10318), .ZN(n10168) );
  OR2_X1 U10909 ( .A1(n31), .A2(n10316), .ZN(n10176) );
  NAND2_X1 U10910 ( .A1(n10168), .A2(n10176), .ZN(n10172) );
  OR2_X1 U10911 ( .A1(n10847), .A2(n10315), .ZN(n10171) );
  OR2_X1 U10912 ( .A1(n10848), .A2(n10314), .ZN(n10179) );
  NAND2_X1 U10913 ( .A1(n10171), .A2(n10179), .ZN(n10181) );
  NOR2_X1 U10914 ( .A1(n10172), .A2(n10181), .ZN(n10173) );
  NAND2_X1 U10915 ( .A1(n10187), .A2(n10173), .ZN(n10189) );
  AND2_X1 U10916 ( .A1(n10508), .A2(n10318), .ZN(n10175) );
  AND2_X1 U10917 ( .A1(n31), .A2(n10316), .ZN(n10174) );
  AOI21_X1 U10918 ( .B1(n10176), .B2(n10175), .A(n10174), .ZN(n10182) );
  AND2_X1 U10919 ( .A1(n10847), .A2(n10315), .ZN(n10178) );
  AND2_X1 U10920 ( .A1(n10848), .A2(n10314), .ZN(n10177) );
  AOI21_X1 U10921 ( .B1(n10179), .B2(n10178), .A(n10177), .ZN(n10180) );
  OAI21_X1 U10922 ( .B1(n10182), .B2(n10181), .A(n10180), .ZN(n10186) );
  NAND2_X1 U10923 ( .A1(data_addr_o_15_), .A2(n3010), .ZN(n12023) );
  NAND2_X1 U10924 ( .A1(n9987), .A2(n6003), .ZN(n10183) );
  OAI21_X1 U10925 ( .B1(n10184), .B2(n12023), .A(n10183), .ZN(n10185) );
  AOI21_X1 U10926 ( .B1(n10187), .B2(n10186), .A(n10185), .ZN(n10188) );
  OAI21_X1 U10927 ( .B1(n10190), .B2(n10189), .A(n10188), .ZN(n10219) );
  OR2_X1 U10928 ( .A1(n10290), .A2(n8444), .ZN(n12055) );
  NAND2_X1 U10929 ( .A1(n10191), .A2(n10857), .ZN(n10192) );
  OAI21_X1 U10930 ( .B1(n10193), .B2(n12055), .A(n10192), .ZN(n10200) );
  NAND2_X1 U10931 ( .A1(n10194), .A2(n9846), .ZN(n10197) );
  NAND2_X1 U10932 ( .A1(n10195), .A2(n10887), .ZN(n10196) );
  OAI21_X1 U10933 ( .B1(n10198), .B2(n10197), .A(n10196), .ZN(n10199) );
  AOI21_X1 U10934 ( .B1(n10201), .B2(n10200), .A(n10199), .ZN(n10217) );
  NAND2_X1 U10935 ( .A1(n34), .A2(n10202), .ZN(n10205) );
  NAND2_X1 U10936 ( .A1(n10203), .A2(n9915), .ZN(n10204) );
  OAI21_X1 U10937 ( .B1(n10206), .B2(n10205), .A(n10204), .ZN(n10213) );
  NAND2_X1 U10938 ( .A1(n10207), .A2(n10898), .ZN(n10210) );
  NAND2_X1 U10939 ( .A1(n10208), .A2(n10899), .ZN(n10209) );
  OAI21_X1 U10940 ( .B1(n10211), .B2(n10210), .A(n10209), .ZN(n10212) );
  AOI21_X1 U10941 ( .B1(n10214), .B2(n10213), .A(n10212), .ZN(n10215) );
  OAI21_X1 U10942 ( .B1(n10217), .B2(n10216), .A(n10215), .ZN(n10218) );
  AOI21_X1 U10943 ( .B1(n10220), .B2(n10219), .A(n10218), .ZN(n10255) );
  INV_X1 U10944 ( .A(n10269), .ZN(n10229) );
  NOR2_X1 U10945 ( .A1(n10229), .A2(n10903), .ZN(n10221) );
  INV_X1 U10946 ( .A(n10268), .ZN(n10230) );
  NOR2_X1 U10947 ( .A1(n10230), .A2(n10267), .ZN(n10233) );
  NOR2_X1 U10948 ( .A1(n10221), .A2(n10233), .ZN(n10223) );
  INV_X1 U10949 ( .A(n10278), .ZN(n10234) );
  NOR2_X1 U10950 ( .A1(n10234), .A2(n10746), .ZN(n10222) );
  NOR2_X1 U10951 ( .A1(n3077), .A2(n10914), .ZN(n10237) );
  NOR2_X1 U10952 ( .A1(n10222), .A2(n10237), .ZN(n10240) );
  NAND2_X1 U10953 ( .A1(n10223), .A2(n10240), .ZN(n10227) );
  INV_X1 U10954 ( .A(n10277), .ZN(n10241) );
  NOR2_X1 U10955 ( .A1(n10241), .A2(n10918), .ZN(n10224) );
  INV_X1 U10956 ( .A(n10258), .ZN(n10242) );
  NOR2_X1 U10957 ( .A1(n10242), .A2(data_addr_o_30_), .ZN(n10245) );
  NOR2_X1 U10958 ( .A1(n10224), .A2(n10245), .ZN(n10226) );
  NOR2_X1 U10959 ( .A1(n3087), .A2(n24), .ZN(n10225) );
  NOR2_X1 U10960 ( .A1(n10225), .A2(pmp_addr_i[350]), .ZN(n10249) );
  NAND2_X1 U10961 ( .A1(n10228), .A2(n3052), .ZN(n10254) );
  NAND2_X1 U10962 ( .A1(n10229), .A2(n10903), .ZN(n10232) );
  NAND2_X1 U10963 ( .A1(n10230), .A2(n10267), .ZN(n10231) );
  OAI21_X1 U10964 ( .B1(n10233), .B2(n10232), .A(n10231), .ZN(n10239) );
  NAND2_X1 U10965 ( .A1(n10234), .A2(n10746), .ZN(n10236) );
  NAND2_X1 U10966 ( .A1(n3077), .A2(n10747), .ZN(n10235) );
  OAI21_X1 U10967 ( .B1(n10237), .B2(n10236), .A(n10235), .ZN(n10238) );
  AOI21_X1 U10968 ( .B1(n10240), .B2(n10239), .A(n10238), .ZN(n10251) );
  NAND2_X1 U10969 ( .A1(n10241), .A2(n10918), .ZN(n10244) );
  NAND2_X1 U10970 ( .A1(n10242), .A2(data_addr_o_30_), .ZN(n10243) );
  OAI21_X1 U10971 ( .B1(n10245), .B2(n10244), .A(n10243), .ZN(n10248) );
  NAND2_X1 U10972 ( .A1(n3087), .A2(n24), .ZN(n10246) );
  NOR2_X1 U10973 ( .A1(n10246), .A2(pmp_addr_i[350]), .ZN(n10247) );
  AOI21_X1 U10974 ( .B1(n10249), .B2(n10248), .A(n10247), .ZN(n10250) );
  NAND2_X1 U10975 ( .A1(n10252), .A2(n3052), .ZN(n10253) );
  OAI21_X1 U10976 ( .B1(n10255), .B2(n10254), .A(n10253), .ZN(n10257) );
  XNOR2_X1 U10977 ( .A(n10258), .B(data_addr_o_30_), .ZN(n10265) );
  XNOR2_X1 U10978 ( .A(n10259), .B(n10899), .ZN(n10264) );
  XNOR2_X1 U10979 ( .A(n10260), .B(n10891), .ZN(n10263) );
  XNOR2_X1 U10980 ( .A(n10261), .B(n10886), .ZN(n10262) );
  NAND4_X1 U10981 ( .A1(n10265), .A2(n10264), .A3(n10263), .A4(n10262), .ZN(
        n10276) );
  XNOR2_X1 U10982 ( .A(n10266), .B(n10747), .ZN(n10274) );
  XNOR2_X1 U10983 ( .A(n10268), .B(n10267), .ZN(n10273) );
  XNOR2_X1 U10984 ( .A(n10269), .B(n9923), .ZN(n10272) );
  XNOR2_X1 U10985 ( .A(n10270), .B(n9915), .ZN(n10271) );
  NAND4_X1 U10986 ( .A1(n10274), .A2(n10273), .A3(n10272), .A4(n10271), .ZN(
        n10275) );
  OR2_X1 U10987 ( .A1(n10276), .A2(n10275), .ZN(n10303) );
  XNOR2_X1 U10988 ( .A(n10277), .B(n10918), .ZN(n10294) );
  XNOR2_X1 U10989 ( .A(n10278), .B(n9886), .ZN(n10293) );
  XNOR2_X1 U10990 ( .A(n10279), .B(data_addr_o_23_), .ZN(n10292) );
  OAI22_X1 U10991 ( .A1(n10314), .A2(data_addr_o_14_), .B1(n11309), .B2(n3010), 
        .ZN(n10284) );
  OAI22_X1 U10992 ( .A1(n11343), .A2(n10317), .B1(n10281), .B2(n10322), .ZN(
        n10283) );
  OAI22_X1 U10993 ( .A1(n10309), .A2(n7816), .B1(n11331), .B2(n10306), .ZN(
        n10282) );
  NOR3_X1 U10994 ( .A1(n10284), .A2(n10283), .A3(n10282), .ZN(n10288) );
  OAI22_X1 U10995 ( .A1(n10318), .A2(data_addr_o_11_), .B1(data_addr_o_9_), 
        .B2(n10305), .ZN(n10286) );
  OAI22_X1 U10996 ( .A1(n10316), .A2(data_addr_o_12_), .B1(data_addr_i[13]), 
        .B2(n10315), .ZN(n10285) );
  NOR2_X1 U10997 ( .A1(n10286), .A2(n10285), .ZN(n10287) );
  NAND2_X1 U10998 ( .A1(n10288), .A2(n10287), .ZN(n10289) );
  AOI21_X1 U10999 ( .B1(n10290), .B2(n8444), .A(n10289), .ZN(n10291) );
  NAND4_X1 U11000 ( .A1(n10294), .A2(n10293), .A3(n10292), .A4(n10291), .ZN(
        n10301) );
  XNOR2_X1 U11001 ( .A(n10296), .B(n10295), .ZN(n10300) );
  XNOR2_X1 U11002 ( .A(n10298), .B(n10297), .ZN(n10299) );
  OR3_X1 U11003 ( .A1(n10301), .A2(n10300), .A3(n10299), .ZN(n10302) );
  NOR2_X1 U11004 ( .A1(n10303), .A2(n10302), .ZN(n12007) );
  XNOR2_X1 U11005 ( .A(n10304), .B(n10107), .ZN(n10330) );
  XNOR2_X1 U11006 ( .A(n12051), .B(n11004), .ZN(n10328) );
  NAND2_X1 U11007 ( .A1(data_addr_o_9_), .A2(n10305), .ZN(n12022) );
  NAND2_X1 U11008 ( .A1(n10358), .A2(n10306), .ZN(n12037) );
  NAND2_X1 U11009 ( .A1(n12022), .A2(n12037), .ZN(n12044) );
  XNOR2_X1 U11010 ( .A(n10824), .B(n10307), .ZN(n10312) );
  XNOR2_X1 U11011 ( .A(n11259), .B(n10308), .ZN(n10310) );
  NAND2_X1 U11012 ( .A1(n7816), .A2(n10309), .ZN(n12038) );
  NAND4_X1 U11013 ( .A1(n10312), .A2(n10311), .A3(n10310), .A4(n12038), .ZN(
        n10313) );
  NOR2_X1 U11014 ( .A1(n12044), .A2(n10313), .ZN(n10327) );
  NAND2_X1 U11015 ( .A1(n9066), .A2(n10314), .ZN(n12036) );
  NAND2_X1 U11016 ( .A1(n6649), .A2(n10315), .ZN(n12012) );
  NAND2_X1 U11017 ( .A1(data_addr_o_12_), .A2(n10316), .ZN(n12017) );
  NAND4_X1 U11018 ( .A1(n12036), .A2(n12023), .A3(n12012), .A4(n12017), .ZN(
        n10325) );
  NAND2_X1 U11019 ( .A1(data_addr_o_10_), .A2(n10317), .ZN(n12011) );
  NAND2_X1 U11020 ( .A1(data_addr_o_11_), .A2(n10318), .ZN(n12016) );
  XNOR2_X1 U11021 ( .A(n11288), .B(n12059), .ZN(n10321) );
  XNOR2_X1 U11022 ( .A(n10958), .B(n10319), .ZN(n10320) );
  NOR2_X1 U11023 ( .A1(n10321), .A2(n10320), .ZN(n10323) );
  NAND2_X1 U11024 ( .A1(n10281), .A2(n10322), .ZN(n12033) );
  NAND4_X1 U11025 ( .A1(n12011), .A2(n12016), .A3(n10323), .A4(n12033), .ZN(
        n10324) );
  NOR2_X1 U11026 ( .A1(n10325), .A2(n10324), .ZN(n10326) );
  NAND4_X1 U11027 ( .A1(n12055), .A2(n10328), .A3(n10327), .A4(n10326), .ZN(
        n10329) );
  NOR2_X1 U11028 ( .A1(n10330), .A2(n10329), .ZN(n10331) );
  OR2_X1 U11029 ( .A1(n11019), .A2(pmp_cfg_i[88]), .ZN(n10334) );
  OAI211_X1 U11030 ( .C1(pmp_cfg_i[89]), .C2(n11021), .A(n10333), .B(n10334), 
        .ZN(n12054) );
  NOR2_X1 U11031 ( .A1(n7990), .A2(pmp_addr_i[206]), .ZN(n10337) );
  NOR2_X1 U11032 ( .A1(pmp_addr_i[207]), .A2(n8757), .ZN(n10389) );
  NOR2_X1 U11033 ( .A1(n10337), .A2(n10389), .ZN(n10392) );
  NOR2_X1 U11034 ( .A1(pmp_addr_i[204]), .A2(n10000), .ZN(n10339) );
  NOR2_X1 U11035 ( .A1(pmp_addr_i[205]), .A2(n10338), .ZN(n10386) );
  NOR2_X1 U11036 ( .A1(n10339), .A2(n10386), .ZN(n10340) );
  NAND2_X1 U11037 ( .A1(n10392), .A2(n10340), .ZN(n10394) );
  NOR2_X1 U11038 ( .A1(pmp_addr_i[200]), .A2(n10701), .ZN(n10341) );
  NOR2_X1 U11039 ( .A1(pmp_addr_i[201]), .A2(n9508), .ZN(n10377) );
  NOR2_X1 U11040 ( .A1(n10341), .A2(n10377), .ZN(n10344) );
  NOR2_X1 U11041 ( .A1(pmp_addr_i[202]), .A2(n10005), .ZN(n10343) );
  NOR2_X1 U11042 ( .A1(pmp_addr_i[203]), .A2(n10342), .ZN(n10380) );
  NOR2_X1 U11043 ( .A1(n10343), .A2(n10380), .ZN(n10383) );
  NAND2_X1 U11044 ( .A1(n10344), .A2(n10383), .ZN(n10345) );
  NOR2_X1 U11045 ( .A1(n10394), .A2(n10345), .ZN(n10398) );
  NOR2_X1 U11046 ( .A1(pmp_addr_i[194]), .A2(n6123), .ZN(n10347) );
  NOR2_X1 U11047 ( .A1(pmp_addr_i[195]), .A2(n10346), .ZN(n10354) );
  NOR2_X1 U11048 ( .A1(n10347), .A2(n10354), .ZN(n10357) );
  NOR2_X1 U11049 ( .A1(pmp_addr_i[193]), .A2(n9350), .ZN(n10350) );
  NAND2_X1 U11050 ( .A1(pmp_addr_i[192]), .A2(n10651), .ZN(n10349) );
  NAND2_X1 U11051 ( .A1(pmp_addr_i[193]), .A2(n9350), .ZN(n10348) );
  OAI21_X1 U11052 ( .B1(n10350), .B2(n10349), .A(n10348), .ZN(n10356) );
  NAND2_X1 U11053 ( .A1(pmp_addr_i[194]), .A2(n10351), .ZN(n10353) );
  NAND2_X1 U11054 ( .A1(pmp_addr_i[195]), .A2(n6127), .ZN(n10352) );
  OAI21_X1 U11055 ( .B1(n10354), .B2(n10353), .A(n10352), .ZN(n10355) );
  AOI21_X1 U11056 ( .B1(n10357), .B2(n10356), .A(n10355), .ZN(n10374) );
  INV_X1 U11057 ( .A(n10358), .ZN(n10362) );
  NOR2_X1 U11058 ( .A1(pmp_addr_i[196]), .A2(n10362), .ZN(n10359) );
  NOR2_X1 U11059 ( .A1(pmp_addr_i[197]), .A2(n6400), .ZN(n10365) );
  NOR2_X1 U11060 ( .A1(n10359), .A2(n10365), .ZN(n10361) );
  NOR2_X1 U11061 ( .A1(pmp_addr_i[198]), .A2(n8735), .ZN(n10360) );
  NOR2_X1 U11062 ( .A1(pmp_addr_i[199]), .A2(n10501), .ZN(n10368) );
  NOR2_X1 U11063 ( .A1(n10360), .A2(n10368), .ZN(n10371) );
  NAND2_X1 U11064 ( .A1(n10361), .A2(n10371), .ZN(n10373) );
  NAND2_X1 U11065 ( .A1(pmp_addr_i[196]), .A2(n10362), .ZN(n10364) );
  NAND2_X1 U11066 ( .A1(pmp_addr_i[197]), .A2(n7152), .ZN(n10363) );
  OAI21_X1 U11067 ( .B1(n10365), .B2(n10364), .A(n10363), .ZN(n10370) );
  NAND2_X1 U11068 ( .A1(pmp_addr_i[198]), .A2(n8735), .ZN(n10367) );
  NAND2_X1 U11069 ( .A1(pmp_addr_i[199]), .A2(n9367), .ZN(n10366) );
  OAI21_X1 U11070 ( .B1(n10368), .B2(n10367), .A(n10366), .ZN(n10369) );
  AOI21_X1 U11071 ( .B1(n10371), .B2(n10370), .A(n10369), .ZN(n10372) );
  OAI21_X1 U11072 ( .B1(n10374), .B2(n10373), .A(n10372), .ZN(n10397) );
  NAND2_X1 U11073 ( .A1(pmp_addr_i[200]), .A2(n10701), .ZN(n10376) );
  NAND2_X1 U11074 ( .A1(pmp_addr_i[201]), .A2(n9508), .ZN(n10375) );
  OAI21_X1 U11075 ( .B1(n10377), .B2(n10376), .A(n10375), .ZN(n10382) );
  NAND2_X1 U11076 ( .A1(pmp_addr_i[202]), .A2(n10005), .ZN(n10379) );
  NAND2_X1 U11077 ( .A1(pmp_addr_i[203]), .A2(n10342), .ZN(n10378) );
  OAI21_X1 U11078 ( .B1(n10380), .B2(n10379), .A(n10378), .ZN(n10381) );
  AOI21_X1 U11079 ( .B1(n10383), .B2(n10382), .A(n10381), .ZN(n10395) );
  NAND2_X1 U11080 ( .A1(pmp_addr_i[204]), .A2(n10000), .ZN(n10385) );
  NAND2_X1 U11081 ( .A1(pmp_addr_i[205]), .A2(n10721), .ZN(n10384) );
  OAI21_X1 U11082 ( .B1(n10386), .B2(n10385), .A(n10384), .ZN(n10391) );
  NAND2_X1 U11083 ( .A1(n10047), .A2(pmp_addr_i[206]), .ZN(n10388) );
  NAND2_X1 U11084 ( .A1(pmp_addr_i[207]), .A2(n7995), .ZN(n10387) );
  OAI21_X1 U11085 ( .B1(n10389), .B2(n10388), .A(n10387), .ZN(n10390) );
  AOI21_X1 U11086 ( .B1(n10392), .B2(n10391), .A(n10390), .ZN(n10393) );
  OAI21_X1 U11087 ( .B1(n10395), .B2(n10394), .A(n10393), .ZN(n10396) );
  AOI21_X1 U11088 ( .B1(n10398), .B2(n10397), .A(n10396), .ZN(n10463) );
  NOR2_X1 U11089 ( .A1(pmp_addr_i[212]), .A2(n9425), .ZN(n10399) );
  INV_X1 U11090 ( .A(n10737), .ZN(n10424) );
  NOR2_X1 U11091 ( .A1(pmp_addr_i[213]), .A2(n10424), .ZN(n10427) );
  NOR2_X1 U11092 ( .A1(n10399), .A2(n10427), .ZN(n10401) );
  INV_X1 U11093 ( .A(data_addr_i[24]), .ZN(n10428) );
  NOR2_X1 U11094 ( .A1(pmp_addr_i[214]), .A2(n10428), .ZN(n10400) );
  INV_X1 U11095 ( .A(n10614), .ZN(n10429) );
  NOR2_X1 U11096 ( .A1(pmp_addr_i[215]), .A2(n10429), .ZN(n10432) );
  NOR2_X1 U11097 ( .A1(n10400), .A2(n10432), .ZN(n10435) );
  NAND2_X1 U11098 ( .A1(n10401), .A2(n10435), .ZN(n10437) );
  NOR2_X1 U11099 ( .A1(pmp_addr_i[211]), .A2(n6192), .ZN(n10420) );
  NOR2_X1 U11100 ( .A1(pmp_addr_i[210]), .A2(n6188), .ZN(n10402) );
  NOR2_X1 U11101 ( .A1(n10420), .A2(n10402), .ZN(n10423) );
  INV_X1 U11102 ( .A(data_addr_i[19]), .ZN(n10414) );
  NOR2_X1 U11103 ( .A1(pmp_addr_i[209]), .A2(n10414), .ZN(n10417) );
  NOR2_X1 U11104 ( .A1(pmp_addr_i[208]), .A2(n10403), .ZN(n10404) );
  NOR2_X1 U11105 ( .A1(n10417), .A2(n10404), .ZN(n10405) );
  NAND2_X1 U11106 ( .A1(n10423), .A2(n10405), .ZN(n10406) );
  NOR2_X1 U11107 ( .A1(n10437), .A2(n10406), .ZN(n10412) );
  INV_X1 U11108 ( .A(data_addr_i[26]), .ZN(n10439) );
  NOR2_X1 U11109 ( .A1(pmp_addr_i[216]), .A2(n10439), .ZN(n10407) );
  NOR2_X1 U11110 ( .A1(pmp_addr_i[217]), .A2(n6212), .ZN(n10442) );
  NOR2_X1 U11111 ( .A1(n10407), .A2(n10442), .ZN(n10409) );
  INV_X1 U11112 ( .A(data_addr_i[28]), .ZN(n10443) );
  NOR2_X1 U11113 ( .A1(pmp_addr_i[218]), .A2(n10443), .ZN(n10408) );
  NOR2_X1 U11114 ( .A1(pmp_addr_i[219]), .A2(n10782), .ZN(n10446) );
  NOR2_X1 U11115 ( .A1(n10408), .A2(n10446), .ZN(n10449) );
  NAND2_X1 U11116 ( .A1(n10409), .A2(n10449), .ZN(n10411) );
  NOR2_X1 U11117 ( .A1(pmp_addr_i[220]), .A2(n8814), .ZN(n10410) );
  NOR2_X1 U11118 ( .A1(pmp_addr_i[221]), .A2(data_addr_o_31__BAR), .ZN(n10452)
         );
  OR2_X1 U11119 ( .A1(n10410), .A2(n10452), .ZN(n10456) );
  NOR2_X1 U11120 ( .A1(n10411), .A2(n10456), .ZN(n10459) );
  NAND2_X1 U11121 ( .A1(n10412), .A2(n10459), .ZN(n10462) );
  NAND2_X1 U11122 ( .A1(pmp_addr_i[208]), .A2(n12184), .ZN(n10416) );
  NAND2_X1 U11123 ( .A1(pmp_addr_i[209]), .A2(n10414), .ZN(n10415) );
  OAI21_X1 U11124 ( .B1(n10417), .B2(n10416), .A(n10415), .ZN(n10422) );
  NAND2_X1 U11125 ( .A1(pmp_addr_i[210]), .A2(n10754), .ZN(n10419) );
  NAND2_X1 U11126 ( .A1(pmp_addr_i[211]), .A2(n9418), .ZN(n10418) );
  OAI21_X1 U11127 ( .B1(n10420), .B2(n10419), .A(n10418), .ZN(n10421) );
  AOI21_X1 U11128 ( .B1(n10423), .B2(n10422), .A(n10421), .ZN(n10438) );
  NAND2_X1 U11129 ( .A1(pmp_addr_i[212]), .A2(n9156), .ZN(n10426) );
  NAND2_X1 U11130 ( .A1(pmp_addr_i[213]), .A2(n10424), .ZN(n10425) );
  OAI21_X1 U11131 ( .B1(n10427), .B2(n10426), .A(n10425), .ZN(n10434) );
  NAND2_X1 U11132 ( .A1(pmp_addr_i[214]), .A2(n10428), .ZN(n10431) );
  NAND2_X1 U11133 ( .A1(pmp_addr_i[215]), .A2(n10429), .ZN(n10430) );
  OAI21_X1 U11134 ( .B1(n10432), .B2(n10431), .A(n10430), .ZN(n10433) );
  AOI21_X1 U11135 ( .B1(n10435), .B2(n10434), .A(n10433), .ZN(n10436) );
  OAI21_X1 U11136 ( .B1(n10438), .B2(n10437), .A(n10436), .ZN(n10460) );
  NAND2_X1 U11137 ( .A1(pmp_addr_i[216]), .A2(n10439), .ZN(n10441) );
  NAND2_X1 U11138 ( .A1(pmp_addr_i[217]), .A2(n9438), .ZN(n10440) );
  OAI21_X1 U11139 ( .B1(n10442), .B2(n10441), .A(n10440), .ZN(n10448) );
  NAND2_X1 U11140 ( .A1(pmp_addr_i[218]), .A2(n10443), .ZN(n10445) );
  NAND2_X1 U11141 ( .A1(pmp_addr_i[219]), .A2(n6216), .ZN(n10444) );
  OAI21_X1 U11142 ( .B1(n10446), .B2(n10445), .A(n10444), .ZN(n10447) );
  AOI21_X1 U11143 ( .B1(n10449), .B2(n10448), .A(n10447), .ZN(n10457) );
  NAND2_X1 U11144 ( .A1(pmp_addr_i[220]), .A2(n8814), .ZN(n10451) );
  NAND2_X1 U11145 ( .A1(pmp_addr_i[221]), .A2(data_addr_o_31__BAR), .ZN(n10450) );
  OAI21_X1 U11146 ( .B1(n10452), .B2(n10451), .A(n10450), .ZN(n10454) );
  NOR2_X1 U11147 ( .A1(n10454), .A2(n397), .ZN(n10455) );
  OAI21_X1 U11148 ( .B1(n10457), .B2(n10456), .A(n10455), .ZN(n10458) );
  AOI21_X1 U11149 ( .B1(n10460), .B2(n10459), .A(n10458), .ZN(n10461) );
  OAI21_X1 U11150 ( .B1(n10463), .B2(n10462), .A(n10461), .ZN(n10593) );
  NOR2_X1 U11151 ( .A1(n11004), .A2(n637), .ZN(n10523) );
  NOR2_X1 U11152 ( .A1(data_addr_o_15_), .A2(n10658), .ZN(n10465) );
  NOR2_X1 U11153 ( .A1(n10523), .A2(n10465), .ZN(n10526) );
  AOI22_X1 U11154 ( .A1(n10519), .A2(n11334), .B1(n10517), .B2(n10466), .ZN(
        n10617) );
  NAND2_X1 U11155 ( .A1(n10526), .A2(n10617), .ZN(n10471) );
  NOR2_X1 U11156 ( .A1(n10530), .A2(n718), .ZN(n10533) );
  NOR2_X1 U11157 ( .A1(n10886), .A2(n742), .ZN(n10467) );
  NOR2_X1 U11158 ( .A1(n10533), .A2(n10467), .ZN(n10536) );
  NOR2_X1 U11159 ( .A1(n10857), .A2(n628), .ZN(n10529) );
  NAND2_X1 U11160 ( .A1(n8757), .A2(n10527), .ZN(n10607) );
  INV_X1 U11161 ( .A(n10607), .ZN(n10469) );
  NOR2_X1 U11162 ( .A1(n10529), .A2(n10469), .ZN(n10470) );
  NAND2_X1 U11163 ( .A1(n10536), .A2(n10470), .ZN(n10538) );
  NOR2_X1 U11164 ( .A1(n10471), .A2(n10538), .ZN(n10542) );
  INV_X1 U11165 ( .A(n10652), .ZN(n10472) );
  NOR2_X1 U11166 ( .A1(n10129), .A2(n10472), .ZN(n10477) );
  NAND2_X1 U11167 ( .A1(n10473), .A2(n10474), .ZN(n10598) );
  INV_X1 U11168 ( .A(n10598), .ZN(n10476) );
  INV_X1 U11169 ( .A(n10474), .ZN(n10475) );
  NAND2_X1 U11170 ( .A1(n22), .A2(n10475), .ZN(n11537) );
  OAI21_X1 U11171 ( .B1(n10477), .B2(n10476), .A(n11537), .ZN(n10482) );
  OR2_X1 U11172 ( .A1(n10479), .A2(n10650), .ZN(n10481) );
  AND2_X1 U11173 ( .A1(n10479), .A2(n10650), .ZN(n10480) );
  AOI21_X1 U11174 ( .B1(n10482), .B2(n10481), .A(n10480), .ZN(n10490) );
  OAI22_X1 U11175 ( .A1(n10654), .A2(n10953), .B1(n11255), .B2(n10483), .ZN(
        n10595) );
  OR2_X1 U11176 ( .A1(n11331), .A2(n10654), .ZN(n10488) );
  AND2_X1 U11177 ( .A1(n10486), .A2(n10483), .ZN(n11544) );
  AND2_X1 U11178 ( .A1(n11331), .A2(n10654), .ZN(n10487) );
  AOI21_X1 U11179 ( .B1(n10488), .B2(n11544), .A(n10487), .ZN(n10489) );
  OAI21_X1 U11180 ( .B1(n10490), .B2(n10595), .A(n10489), .ZN(n10497) );
  NOR2_X1 U11181 ( .A1(n10494), .A2(n672), .ZN(n10594) );
  NOR2_X1 U11182 ( .A1(n10493), .A2(n4843), .ZN(n10600) );
  NOR2_X1 U11183 ( .A1(n10594), .A2(n10600), .ZN(n10496) );
  NAND2_X1 U11184 ( .A1(n10493), .A2(n4843), .ZN(n11547) );
  NAND2_X1 U11185 ( .A1(n10494), .A2(n672), .ZN(n11541) );
  OAI21_X1 U11186 ( .B1(n10594), .B2(n11547), .A(n11541), .ZN(n10495) );
  AOI21_X1 U11187 ( .B1(n10497), .B2(n10496), .A(n10495), .ZN(n10515) );
  OAI22_X1 U11188 ( .A1(n10500), .A2(n10499), .B1(n10498), .B2(data_addr_o_11_), .ZN(n10603) );
  INV_X1 U11189 ( .A(n10603), .ZN(n10512) );
  AOI22_X1 U11190 ( .A1(n10502), .A2(n10701), .B1(n10501), .B2(n10503), .ZN(
        n10608) );
  NAND2_X1 U11191 ( .A1(n10512), .A2(n10608), .ZN(n10514) );
  NOR2_X1 U11192 ( .A1(n10838), .A2(n643), .ZN(n10505) );
  NAND2_X1 U11193 ( .A1(n10504), .A2(n4848), .ZN(n11529) );
  NAND2_X1 U11194 ( .A1(n10838), .A2(n643), .ZN(n11527) );
  OAI21_X1 U11195 ( .B1(n10505), .B2(n11529), .A(n11527), .ZN(n10511) );
  NOR2_X1 U11196 ( .A1(n31), .A2(n10500), .ZN(n10509) );
  NAND2_X1 U11197 ( .A1(n10508), .A2(n10498), .ZN(n11552) );
  NAND2_X1 U11198 ( .A1(n31), .A2(n10500), .ZN(n11520) );
  OAI21_X1 U11199 ( .B1(n10509), .B2(n11552), .A(n11520), .ZN(n10510) );
  AOI21_X1 U11200 ( .B1(n10512), .B2(n10511), .A(n10510), .ZN(n10513) );
  OAI21_X1 U11201 ( .B1(n10515), .B2(n10514), .A(n10513), .ZN(n10541) );
  INV_X1 U11202 ( .A(n10519), .ZN(n10516) );
  NOR2_X1 U11203 ( .A1(n10516), .A2(n10848), .ZN(n10520) );
  OR2_X1 U11204 ( .A1(n10517), .A2(n11006), .ZN(n11566) );
  OR2_X1 U11205 ( .A1(n10519), .A2(n10518), .ZN(n11560) );
  OAI21_X1 U11206 ( .B1(n10520), .B2(n11566), .A(n11560), .ZN(n10525) );
  NAND2_X1 U11207 ( .A1(data_addr_o_15_), .A2(n10658), .ZN(n10522) );
  NAND2_X1 U11208 ( .A1(n11004), .A2(n637), .ZN(n10521) );
  OAI21_X1 U11209 ( .B1(n10523), .B2(n10522), .A(n10521), .ZN(n10524) );
  AOI21_X1 U11210 ( .B1(n10526), .B2(n10525), .A(n10524), .ZN(n10539) );
  NAND2_X1 U11211 ( .A1(data_addr_o_17_), .A2(n4857), .ZN(n11559) );
  NAND2_X1 U11212 ( .A1(n10857), .A2(n628), .ZN(n10528) );
  OAI21_X1 U11213 ( .B1(n10529), .B2(n11559), .A(n10528), .ZN(n10535) );
  NAND2_X1 U11214 ( .A1(n10886), .A2(n742), .ZN(n10532) );
  NAND2_X1 U11215 ( .A1(n10530), .A2(n718), .ZN(n10531) );
  OAI21_X1 U11216 ( .B1(n10533), .B2(n10532), .A(n10531), .ZN(n10534) );
  AOI21_X1 U11217 ( .B1(n10536), .B2(n10535), .A(n10534), .ZN(n10537) );
  OAI21_X1 U11218 ( .B1(n10539), .B2(n10538), .A(n10537), .ZN(n10540) );
  AOI21_X1 U11219 ( .B1(n10542), .B2(n10541), .A(n10540), .ZN(n10591) );
  NOR2_X1 U11220 ( .A1(n9529), .A2(n713), .ZN(n10557) );
  NOR2_X1 U11221 ( .A1(n10891), .A2(n746), .ZN(n10543) );
  NOR2_X1 U11222 ( .A1(n10557), .A2(n10543), .ZN(n10545) );
  INV_X1 U11223 ( .A(n10628), .ZN(n10558) );
  NOR2_X1 U11224 ( .A1(n10899), .A2(n10558), .ZN(n10561) );
  NOR2_X1 U11225 ( .A1(n10898), .A2(n768), .ZN(n10544) );
  NOR2_X1 U11226 ( .A1(n10561), .A2(n10544), .ZN(n10564) );
  NAND2_X1 U11227 ( .A1(n10545), .A2(n10564), .ZN(n10549) );
  NOR2_X1 U11228 ( .A1(n10914), .A2(n731), .ZN(n10570) );
  NOR2_X1 U11229 ( .A1(n11322), .A2(n753), .ZN(n10546) );
  NOR2_X1 U11230 ( .A1(n10570), .A2(n10546), .ZN(n10573) );
  NOR2_X1 U11231 ( .A1(data_addr_o_26_), .A2(n698), .ZN(n10567) );
  NOR2_X1 U11232 ( .A1(n10903), .A2(n771), .ZN(n10547) );
  NOR2_X1 U11233 ( .A1(n10567), .A2(n10547), .ZN(n10548) );
  NAND2_X1 U11234 ( .A1(n10573), .A2(n10548), .ZN(n10575) );
  NOR2_X1 U11235 ( .A1(n10549), .A2(n10575), .ZN(n10554) );
  INV_X1 U11236 ( .A(n10661), .ZN(n10580) );
  NOR2_X1 U11237 ( .A1(n10580), .A2(n24), .ZN(n10550) );
  NOR2_X1 U11238 ( .A1(n10550), .A2(pmp_addr_i[190]), .ZN(n10584) );
  NOR2_X1 U11239 ( .A1(data_addr_o_30_), .A2(n724), .ZN(n10579) );
  NOR2_X1 U11240 ( .A1(n10918), .A2(n756), .ZN(n10551) );
  NOR2_X1 U11241 ( .A1(n10579), .A2(n10551), .ZN(n10552) );
  NAND2_X1 U11242 ( .A1(n10584), .A2(n10552), .ZN(n10553) );
  NOR2_X1 U11243 ( .A1(n10553), .A2(pmp_addr_i[191]), .ZN(n10587) );
  NAND2_X1 U11244 ( .A1(n10554), .A2(n10587), .ZN(n10590) );
  NAND2_X1 U11245 ( .A1(n10891), .A2(n746), .ZN(n10556) );
  NAND2_X1 U11246 ( .A1(n11313), .A2(n713), .ZN(n10555) );
  OAI21_X1 U11247 ( .B1(n10557), .B2(n10556), .A(n10555), .ZN(n10563) );
  NAND2_X1 U11248 ( .A1(n10898), .A2(n768), .ZN(n10560) );
  NAND2_X1 U11249 ( .A1(n10899), .A2(n10558), .ZN(n10559) );
  OAI21_X1 U11250 ( .B1(n10561), .B2(n10560), .A(n10559), .ZN(n10562) );
  AOI21_X1 U11251 ( .B1(n10564), .B2(n10563), .A(n10562), .ZN(n10576) );
  NAND2_X1 U11252 ( .A1(n10903), .A2(n771), .ZN(n10566) );
  NAND2_X1 U11253 ( .A1(data_addr_o_26_), .A2(n698), .ZN(n10565) );
  OAI21_X1 U11254 ( .B1(n10567), .B2(n10566), .A(n10565), .ZN(n10572) );
  NAND2_X1 U11255 ( .A1(n9886), .A2(n753), .ZN(n10569) );
  NAND2_X1 U11256 ( .A1(n10914), .A2(n731), .ZN(n10568) );
  OAI21_X1 U11257 ( .B1(n10570), .B2(n10569), .A(n10568), .ZN(n10571) );
  AOI21_X1 U11258 ( .B1(n10573), .B2(n10572), .A(n10571), .ZN(n10574) );
  OAI21_X1 U11259 ( .B1(n10576), .B2(n10575), .A(n10574), .ZN(n10588) );
  NAND2_X1 U11260 ( .A1(n10918), .A2(n756), .ZN(n10578) );
  NAND2_X1 U11261 ( .A1(n10919), .A2(n724), .ZN(n10577) );
  OAI21_X1 U11262 ( .B1(n10579), .B2(n10578), .A(n10577), .ZN(n10583) );
  NAND2_X1 U11263 ( .A1(n10580), .A2(n24), .ZN(n10581) );
  NOR2_X1 U11264 ( .A1(n10581), .A2(pmp_addr_i[190]), .ZN(n10582) );
  AOI21_X1 U11265 ( .B1(n10584), .B2(n10583), .A(n10582), .ZN(n10585) );
  NOR2_X1 U11266 ( .A1(n10585), .A2(pmp_addr_i[191]), .ZN(n10586) );
  AOI21_X1 U11267 ( .B1(n10588), .B2(n10587), .A(n10586), .ZN(n10589) );
  OAI21_X1 U11268 ( .B1(n10591), .B2(n10590), .A(n10589), .ZN(n10592) );
  NAND3_X1 U11269 ( .A1(n10593), .A2(n878), .A3(n10592), .ZN(n10673) );
  NOR2_X1 U11270 ( .A1(n10595), .A2(n10594), .ZN(n10602) );
  AOI21_X1 U11271 ( .B1(n10651), .B2(n10652), .A(n10596), .ZN(n10597) );
  OAI211_X1 U11272 ( .C1(n10650), .C2(n11288), .A(n10598), .B(n10597), .ZN(
        n10599) );
  NOR2_X1 U11273 ( .A1(n10600), .A2(n10599), .ZN(n10601) );
  OAI211_X1 U11274 ( .C1(n10658), .C2(n10657), .A(n10602), .B(n10601), .ZN(
        n10604) );
  NOR2_X1 U11275 ( .A1(n10604), .A2(n10603), .ZN(n10610) );
  XNOR2_X1 U11276 ( .A(n10606), .B(n10605), .ZN(n10609) );
  NAND4_X1 U11277 ( .A1(n10610), .A2(n10609), .A3(n10608), .A4(n10607), .ZN(
        n10622) );
  XNOR2_X1 U11278 ( .A(n10612), .B(n10611), .ZN(n10620) );
  XNOR2_X1 U11279 ( .A(n10614), .B(n10613), .ZN(n10619) );
  XNOR2_X1 U11280 ( .A(n10616), .B(n10615), .ZN(n10618) );
  NAND4_X1 U11281 ( .A1(n10620), .A2(n10619), .A3(n10618), .A4(n10617), .ZN(
        n10621) );
  NOR2_X1 U11282 ( .A1(n10622), .A2(n10621), .ZN(n10647) );
  XNOR2_X1 U11283 ( .A(n10919), .B(n10623), .ZN(n10633) );
  XNOR2_X1 U11284 ( .A(n10967), .B(n10625), .ZN(n10632) );
  XNOR2_X1 U11285 ( .A(n10627), .B(n10626), .ZN(n10631) );
  XNOR2_X1 U11286 ( .A(n10629), .B(n10628), .ZN(n10630) );
  NAND4_X1 U11287 ( .A1(n10633), .A2(n10632), .A3(n10631), .A4(n10630), .ZN(
        n10645) );
  XNOR2_X1 U11288 ( .A(n10635), .B(n10634), .ZN(n10643) );
  XNOR2_X1 U11289 ( .A(n10530), .B(n10636), .ZN(n10642) );
  XNOR2_X1 U11290 ( .A(n10638), .B(n10637), .ZN(n10641) );
  XNOR2_X1 U11291 ( .A(data_addr_o_23_), .B(n10639), .ZN(n10640) );
  NAND4_X1 U11292 ( .A1(n10643), .A2(n10642), .A3(n10641), .A4(n10640), .ZN(
        n10644) );
  NOR2_X1 U11293 ( .A1(n10645), .A2(n10644), .ZN(n10646) );
  XNOR2_X1 U11295 ( .A(n11303), .B(n10648), .ZN(n11574) );
  NAND2_X1 U11296 ( .A1(data_addr_o_4_), .A2(n10650), .ZN(n11536) );
  OAI211_X1 U11297 ( .C1(n10652), .C2(n10651), .A(n11536), .B(n11537), .ZN(
        n10653) );
  NOR2_X1 U11298 ( .A1(n11544), .A2(n10653), .ZN(n10656) );
  NAND2_X1 U11299 ( .A1(n10655), .A2(n10654), .ZN(n11534) );
  NAND4_X1 U11300 ( .A1(n10656), .A2(n11541), .A3(n11547), .A4(n11534), .ZN(
        n10659) );
  AND2_X1 U11301 ( .A1(n10658), .A2(n10657), .ZN(n11523) );
  NOR2_X1 U11302 ( .A1(n10659), .A2(n11523), .ZN(n10660) );
  NAND4_X1 U11303 ( .A1(n10660), .A2(n11560), .A3(n11520), .A4(n11552), .ZN(
        n10664) );
  XOR2_X1 U11304 ( .A(n10662), .B(n10661), .Z(n10663) );
  NOR2_X1 U11305 ( .A1(n10664), .A2(n10663), .ZN(n10669) );
  NAND2_X1 U11306 ( .A1(n11559), .A2(n11566), .ZN(n10667) );
  XNOR2_X1 U11307 ( .A(n11004), .B(n11568), .ZN(n10665) );
  NAND3_X1 U11308 ( .A1(n10665), .A2(n11527), .A3(n11529), .ZN(n10666) );
  NOR2_X1 U11309 ( .A1(n10667), .A2(n10666), .ZN(n10668) );
  NAND4_X1 U11310 ( .A1(n11519), .A2(n11574), .A3(n10669), .A4(n10668), .ZN(
        n10672) );
  MUX2_X1 U11311 ( .A(pmp_cfg_i[48]), .B(pmp_cfg_i[49]), .S(n11019), .Z(n10671) );
  NAND2_X1 U11312 ( .A1(n10670), .A2(n10671), .ZN(n11549) );
  AOI21_X1 U11313 ( .B1(n10673), .B2(n10672), .A(n11549), .ZN(n11025) );
  NOR2_X1 U11314 ( .A1(n10047), .A2(pmp_addr_i[174]), .ZN(n10724) );
  INV_X1 U11315 ( .A(n11227), .ZN(n10721) );
  NOR2_X1 U11316 ( .A1(n10721), .A2(pmp_addr_i[173]), .ZN(n10674) );
  NOR2_X1 U11317 ( .A1(n10724), .A2(n10674), .ZN(n10676) );
  NOR2_X1 U11318 ( .A1(n10060), .A2(pmp_addr_i[176]), .ZN(n10727) );
  NOR2_X1 U11319 ( .A1(n7995), .A2(pmp_addr_i[175]), .ZN(n10675) );
  NOR2_X1 U11320 ( .A1(n10727), .A2(n10675), .ZN(n10729) );
  NAND2_X1 U11321 ( .A1(n10676), .A2(n10729), .ZN(n10733) );
  INV_X1 U11322 ( .A(data_addr_o_11_), .ZN(n10711) );
  NOR2_X1 U11323 ( .A1(n10711), .A2(pmp_addr_i[169]), .ZN(n10677) );
  NOR2_X1 U11324 ( .A1(n9947), .A2(pmp_addr_i[170]), .ZN(n10714) );
  NOR2_X1 U11325 ( .A1(n10677), .A2(n10714), .ZN(n10679) );
  NOR2_X1 U11326 ( .A1(n11006), .A2(pmp_addr_i[171]), .ZN(n10678) );
  NOR2_X1 U11327 ( .A1(n6154), .A2(pmp_addr_i[172]), .ZN(n10717) );
  NOR2_X1 U11328 ( .A1(n10678), .A2(n10717), .ZN(n10720) );
  NAND2_X1 U11329 ( .A1(n10679), .A2(n10720), .ZN(n10680) );
  NOR2_X1 U11330 ( .A1(n10733), .A2(n10680), .ZN(n10736) );
  NOR2_X1 U11331 ( .A1(n6127), .A2(pmp_addr_i[163]), .ZN(n10681) );
  NOR2_X1 U11332 ( .A1(n10362), .A2(pmp_addr_i[164]), .ZN(n10690) );
  NOR2_X1 U11333 ( .A1(n10681), .A2(n10690), .ZN(n10693) );
  OR2_X1 U11334 ( .A1(n9350), .A2(pmp_addr_i[161]), .ZN(n10684) );
  AND2_X1 U11335 ( .A1(n10651), .A2(pmp_addr_i[160]), .ZN(n10683) );
  AND2_X1 U11336 ( .A1(n9350), .A2(pmp_addr_i[161]), .ZN(n10682) );
  AOI21_X1 U11337 ( .B1(n10684), .B2(n10683), .A(n10682), .ZN(n10687) );
  NOR2_X1 U11338 ( .A1(n8406), .A2(pmp_addr_i[162]), .ZN(n10686) );
  NAND2_X1 U11339 ( .A1(n6123), .A2(pmp_addr_i[162]), .ZN(n10685) );
  OAI21_X1 U11340 ( .B1(n10687), .B2(n10686), .A(n10685), .ZN(n10692) );
  NAND2_X1 U11341 ( .A1(n6127), .A2(pmp_addr_i[163]), .ZN(n10689) );
  NAND2_X1 U11342 ( .A1(n9363), .A2(pmp_addr_i[164]), .ZN(n10688) );
  OAI21_X1 U11343 ( .B1(n10690), .B2(n10689), .A(n10688), .ZN(n10691) );
  AOI21_X1 U11344 ( .B1(n10693), .B2(n10692), .A(n10691), .ZN(n10710) );
  NOR2_X1 U11345 ( .A1(n8735), .A2(pmp_addr_i[166]), .ZN(n10700) );
  INV_X1 U11346 ( .A(n7816), .ZN(n10697) );
  NOR2_X1 U11347 ( .A1(n10697), .A2(pmp_addr_i[165]), .ZN(n10694) );
  NOR2_X1 U11348 ( .A1(n10700), .A2(n10694), .ZN(n10696) );
  NOR2_X1 U11349 ( .A1(n6140), .A2(pmp_addr_i[167]), .ZN(n10695) );
  NOR2_X1 U11351 ( .A1(n10701), .A2(pmp_addr_i[168]), .ZN(n10704) );
  NOR2_X1 U11352 ( .A1(n10695), .A2(n10704), .ZN(n10707) );
  NAND2_X1 U11353 ( .A1(n10696), .A2(n10707), .ZN(n10709) );
  NAND2_X1 U11354 ( .A1(n10697), .A2(pmp_addr_i[165]), .ZN(n10699) );
  NAND2_X1 U11355 ( .A1(n8735), .A2(pmp_addr_i[166]), .ZN(n10698) );
  OAI21_X1 U11356 ( .B1(n10700), .B2(n10699), .A(n10698), .ZN(n10706) );
  NAND2_X1 U11357 ( .A1(n10501), .A2(pmp_addr_i[167]), .ZN(n10703) );
  NAND2_X1 U11358 ( .A1(n10701), .A2(pmp_addr_i[168]), .ZN(n10702) );
  OAI21_X1 U11359 ( .B1(n10704), .B2(n10703), .A(n10702), .ZN(n10705) );
  AOI21_X1 U11360 ( .B1(n10707), .B2(n10706), .A(n10705), .ZN(n10708) );
  OAI21_X1 U11361 ( .B1(n10710), .B2(n10709), .A(n10708), .ZN(n10735) );
  NAND2_X1 U11362 ( .A1(n10711), .A2(pmp_addr_i[169]), .ZN(n10713) );
  NAND2_X1 U11363 ( .A1(n7976), .A2(pmp_addr_i[170]), .ZN(n10712) );
  OAI21_X1 U11364 ( .B1(n10714), .B2(n10713), .A(n10712), .ZN(n10719) );
  NAND2_X1 U11365 ( .A1(n10342), .A2(pmp_addr_i[171]), .ZN(n10716) );
  NAND2_X1 U11366 ( .A1(n6154), .A2(pmp_addr_i[172]), .ZN(n10715) );
  OAI21_X1 U11367 ( .B1(n10717), .B2(n10716), .A(n10715), .ZN(n10718) );
  AOI21_X1 U11368 ( .B1(n10720), .B2(n10719), .A(n10718), .ZN(n10732) );
  NAND2_X1 U11369 ( .A1(n10721), .A2(pmp_addr_i[173]), .ZN(n10723) );
  NAND2_X1 U11370 ( .A1(n7057), .A2(pmp_addr_i[174]), .ZN(n10722) );
  OAI21_X1 U11371 ( .B1(n10724), .B2(n10723), .A(n10722), .ZN(n10730) );
  NAND2_X1 U11372 ( .A1(n8757), .A2(pmp_addr_i[175]), .ZN(n10726) );
  NAND2_X1 U11373 ( .A1(n10060), .A2(pmp_addr_i[176]), .ZN(n10725) );
  OAI21_X1 U11374 ( .B1(n10727), .B2(n10726), .A(n10725), .ZN(n10728) );
  AOI21_X1 U11375 ( .B1(n10730), .B2(n10729), .A(n10728), .ZN(n10731) );
  OAI21_X1 U11376 ( .B1(n10733), .B2(n10732), .A(n10731), .ZN(n10734) );
  AOI21_X1 U11377 ( .B1(n10736), .B2(n10735), .A(n10734), .ZN(n10800) );
  INV_X1 U11378 ( .A(n10737), .ZN(n10764) );
  NOR2_X1 U11379 ( .A1(n10764), .A2(pmp_addr_i[181]), .ZN(n10739) );
  NOR2_X1 U11380 ( .A1(n10428), .A2(pmp_addr_i[182]), .ZN(n10767) );
  NOR2_X1 U11381 ( .A1(n10739), .A2(n10767), .ZN(n10741) );
  INV_X1 U11382 ( .A(n10903), .ZN(n10768) );
  NOR2_X1 U11383 ( .A1(n10768), .A2(pmp_addr_i[183]), .ZN(n10740) );
  NOR2_X1 U11384 ( .A1(n10439), .A2(pmp_addr_i[184]), .ZN(n10771) );
  NOR2_X1 U11385 ( .A1(n10740), .A2(n10771), .ZN(n10774) );
  NAND2_X1 U11386 ( .A1(n10741), .A2(n10774), .ZN(n10776) );
  NOR2_X1 U11387 ( .A1(n9418), .A2(pmp_addr_i[179]), .ZN(n10742) );
  NOR2_X1 U11388 ( .A1(n9425), .A2(pmp_addr_i[180]), .ZN(n10760) );
  NOR2_X1 U11389 ( .A1(n10742), .A2(n10760), .ZN(n10763) );
  INV_X1 U11390 ( .A(n10886), .ZN(n10753) );
  NOR2_X1 U11391 ( .A1(n10753), .A2(pmp_addr_i[177]), .ZN(n10743) );
  INV_X1 U11392 ( .A(data_addr_i[20]), .ZN(n10754) );
  NOR2_X1 U11393 ( .A1(n10754), .A2(pmp_addr_i[178]), .ZN(n10757) );
  NOR2_X1 U11394 ( .A1(n10743), .A2(n10757), .ZN(n10744) );
  NAND2_X1 U11395 ( .A1(n10763), .A2(n10744), .ZN(n10745) );
  NOR2_X1 U11396 ( .A1(n10776), .A2(n10745), .ZN(n10752) );
  NOR2_X1 U11397 ( .A1(n6212), .A2(pmp_addr_i[185]), .ZN(n10748) );
  INV_X1 U11398 ( .A(n10747), .ZN(n10778) );
  NOR2_X1 U11399 ( .A1(n10778), .A2(pmp_addr_i[186]), .ZN(n10781) );
  NOR2_X1 U11400 ( .A1(n10748), .A2(n10781), .ZN(n10750) );
  INV_X1 U11401 ( .A(data_addr_o_29_), .ZN(n10782) );
  NOR2_X1 U11402 ( .A1(n10782), .A2(pmp_addr_i[187]), .ZN(n10749) );
  NOR2_X1 U11403 ( .A1(n8814), .A2(pmp_addr_i[188]), .ZN(n10785) );
  NOR2_X1 U11404 ( .A1(n10749), .A2(n10785), .ZN(n10788) );
  NAND2_X1 U11405 ( .A1(n10750), .A2(n10788), .ZN(n10751) );
  NOR2_X1 U11406 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[189]), .ZN(n10793)
         );
  NOR2_X1 U11407 ( .A1(n10751), .A2(n10793), .ZN(n10796) );
  NAND2_X1 U11408 ( .A1(n10752), .A2(n10796), .ZN(n10799) );
  NAND2_X1 U11409 ( .A1(n10753), .A2(pmp_addr_i[177]), .ZN(n10756) );
  NAND2_X1 U11410 ( .A1(n10754), .A2(pmp_addr_i[178]), .ZN(n10755) );
  OAI21_X1 U11411 ( .B1(n10757), .B2(n10756), .A(n10755), .ZN(n10762) );
  NAND2_X1 U11412 ( .A1(n6192), .A2(pmp_addr_i[179]), .ZN(n10759) );
  NAND2_X1 U11413 ( .A1(n9156), .A2(pmp_addr_i[180]), .ZN(n10758) );
  OAI21_X1 U11414 ( .B1(n10760), .B2(n10759), .A(n10758), .ZN(n10761) );
  AOI21_X1 U11415 ( .B1(n10763), .B2(n10762), .A(n10761), .ZN(n10777) );
  NAND2_X1 U11416 ( .A1(n10764), .A2(pmp_addr_i[181]), .ZN(n10766) );
  NAND2_X1 U11417 ( .A1(n9163), .A2(pmp_addr_i[182]), .ZN(n10765) );
  OAI21_X1 U11418 ( .B1(n10767), .B2(n10766), .A(n10765), .ZN(n10773) );
  NAND2_X1 U11419 ( .A1(n10768), .A2(pmp_addr_i[183]), .ZN(n10770) );
  NAND2_X1 U11420 ( .A1(n6202), .A2(pmp_addr_i[184]), .ZN(n10769) );
  OAI21_X1 U11421 ( .B1(n10771), .B2(n10770), .A(n10769), .ZN(n10772) );
  AOI21_X1 U11422 ( .B1(n10774), .B2(n10773), .A(n10772), .ZN(n10775) );
  OAI21_X1 U11423 ( .B1(n10777), .B2(n10776), .A(n10775), .ZN(n10797) );
  NAND2_X1 U11424 ( .A1(n6212), .A2(pmp_addr_i[185]), .ZN(n10780) );
  NAND2_X1 U11425 ( .A1(n10778), .A2(pmp_addr_i[186]), .ZN(n10779) );
  OAI21_X1 U11426 ( .B1(n10781), .B2(n10780), .A(n10779), .ZN(n10787) );
  NAND2_X1 U11427 ( .A1(n10782), .A2(pmp_addr_i[187]), .ZN(n10784) );
  NAND2_X1 U11428 ( .A1(n8494), .A2(pmp_addr_i[188]), .ZN(n10783) );
  OAI21_X1 U11429 ( .B1(n10785), .B2(n10784), .A(n10783), .ZN(n10786) );
  AOI21_X1 U11430 ( .B1(n10788), .B2(n10787), .A(n10786), .ZN(n10794) );
  NAND2_X1 U11431 ( .A1(data_addr_o_31__BAR), .A2(pmp_addr_i[189]), .ZN(n10790) );
  INV_X1 U11432 ( .A(pmp_addr_i[190]), .ZN(n10789) );
  NAND2_X1 U11433 ( .A1(n10790), .A2(n10789), .ZN(n10791) );
  NOR2_X1 U11434 ( .A1(n10791), .A2(pmp_addr_i[191]), .ZN(n10792) );
  OAI21_X1 U11435 ( .B1(n10794), .B2(n10793), .A(n10792), .ZN(n10795) );
  AOI21_X1 U11436 ( .B1(n10797), .B2(n10796), .A(n10795), .ZN(n10798) );
  OAI21_X1 U11437 ( .B1(n10800), .B2(n10799), .A(n10798), .ZN(n10938) );
  NOR2_X1 U11438 ( .A1(n10857), .A2(n5220), .ZN(n10860) );
  INV_X1 U11439 ( .A(n10965), .ZN(n10856) );
  NOR2_X1 U11440 ( .A1(n6813), .A2(n10856), .ZN(n10801) );
  NOR2_X1 U11441 ( .A1(n10860), .A2(n10801), .ZN(n10863) );
  NOR2_X1 U11442 ( .A1(n11004), .A2(n11015), .ZN(n10855) );
  NOR2_X1 U11443 ( .A1(n11309), .A2(n10948), .ZN(n10804) );
  NOR2_X1 U11444 ( .A1(n10855), .A2(n10804), .ZN(n10805) );
  NAND2_X1 U11445 ( .A1(n10863), .A2(n10805), .ZN(n10866) );
  NOR2_X1 U11446 ( .A1(n10508), .A2(n10946), .ZN(n10808) );
  NOR2_X1 U11447 ( .A1(n31), .A2(n10939), .ZN(n10846) );
  NOR2_X1 U11448 ( .A1(n10808), .A2(n10846), .ZN(n10811) );
  NOR2_X1 U11449 ( .A1(n10847), .A2(n10947), .ZN(n10810) );
  NOR2_X1 U11450 ( .A1(n10848), .A2(n10945), .ZN(n10850) );
  NOR2_X1 U11451 ( .A1(n10810), .A2(n10850), .ZN(n10853) );
  NAND2_X1 U11452 ( .A1(n10811), .A2(n10853), .ZN(n10812) );
  NOR2_X1 U11453 ( .A1(n10866), .A2(n10812), .ZN(n10869) );
  NOR2_X1 U11454 ( .A1(n10824), .A2(n10963), .ZN(n10815) );
  NOR2_X1 U11455 ( .A1(data_addr_o_6_), .A2(n10952), .ZN(n10825) );
  NOR2_X1 U11456 ( .A1(n10815), .A2(n10825), .ZN(n10828) );
  INV_X1 U11457 ( .A(n10957), .ZN(n10816) );
  OR2_X1 U11458 ( .A1(data_addr_o_2_), .A2(n10816), .ZN(n10821) );
  INV_X1 U11459 ( .A(n10956), .ZN(n10817) );
  OR2_X1 U11460 ( .A1(n10818), .A2(n10817), .ZN(n10820) );
  AND2_X1 U11461 ( .A1(n10818), .A2(n10817), .ZN(n10819) );
  AOI21_X1 U11462 ( .B1(n10821), .B2(n10820), .A(n10819), .ZN(n10823) );
  NOR2_X1 U11463 ( .A1(n10135), .A2(n5898), .ZN(n10822) );
  NAND2_X1 U11464 ( .A1(n10479), .A2(n5898), .ZN(n11379) );
  OAI21_X1 U11465 ( .B1(n10823), .B2(n10822), .A(n11379), .ZN(n10827) );
  NAND2_X1 U11466 ( .A1(n10824), .A2(n10963), .ZN(n11373) );
  NAND2_X1 U11467 ( .A1(data_addr_o_6_), .A2(n10952), .ZN(n11374) );
  OAI21_X1 U11468 ( .B1(n10825), .B2(n11373), .A(n11374), .ZN(n10826) );
  AOI21_X1 U11469 ( .B1(n10828), .B2(n10827), .A(n10826), .ZN(n10845) );
  NOR2_X1 U11470 ( .A1(n10836), .A2(n10941), .ZN(n10837) );
  NOR2_X1 U11471 ( .A1(n7816), .A2(n10954), .ZN(n10831) );
  NOR2_X1 U11472 ( .A1(n10837), .A2(n10831), .ZN(n10835) );
  NOR2_X1 U11473 ( .A1(data_addr_o_9_), .A2(n10940), .ZN(n10834) );
  NOR2_X1 U11474 ( .A1(n10838), .A2(n10942), .ZN(n10839) );
  NOR2_X1 U11475 ( .A1(n10834), .A2(n10839), .ZN(n10842) );
  NAND2_X1 U11476 ( .A1(n10835), .A2(n10842), .ZN(n10844) );
  NAND2_X1 U11477 ( .A1(n7816), .A2(n10954), .ZN(n11387) );
  NAND2_X1 U11478 ( .A1(n10836), .A2(n10941), .ZN(n11363) );
  OAI21_X1 U11479 ( .B1(n10837), .B2(n11387), .A(n11363), .ZN(n10841) );
  NAND2_X1 U11480 ( .A1(n8237), .A2(n10940), .ZN(n11360) );
  NAND2_X1 U11481 ( .A1(n10838), .A2(n10942), .ZN(n11356) );
  OAI21_X1 U11482 ( .B1(n10839), .B2(n11360), .A(n11356), .ZN(n10840) );
  AOI21_X1 U11483 ( .B1(n10842), .B2(n10841), .A(n10840), .ZN(n10843) );
  OAI21_X1 U11484 ( .B1(n10845), .B2(n10844), .A(n10843), .ZN(n10868) );
  NAND2_X1 U11485 ( .A1(n8246), .A2(n10946), .ZN(n11396) );
  NAND2_X1 U11486 ( .A1(n31), .A2(n10939), .ZN(n11394) );
  OAI21_X1 U11487 ( .B1(n10846), .B2(n11396), .A(n11394), .ZN(n10852) );
  NAND2_X1 U11488 ( .A1(n10847), .A2(n10947), .ZN(n10849) );
  NAND2_X1 U11489 ( .A1(n10848), .A2(n10945), .ZN(n11359) );
  OAI21_X1 U11490 ( .B1(n10850), .B2(n10849), .A(n11359), .ZN(n10851) );
  AOI21_X1 U11491 ( .B1(n10853), .B2(n10852), .A(n10851), .ZN(n10865) );
  NAND2_X1 U11492 ( .A1(n11309), .A2(n10948), .ZN(n11365) );
  NAND2_X1 U11493 ( .A1(n11004), .A2(n11015), .ZN(n10854) );
  OAI21_X1 U11494 ( .B1(n10855), .B2(n11365), .A(n10854), .ZN(n10862) );
  NAND2_X1 U11495 ( .A1(data_addr_o_17_), .A2(n10856), .ZN(n10859) );
  NAND2_X1 U11496 ( .A1(n10857), .A2(n5220), .ZN(n10858) );
  OAI21_X1 U11497 ( .B1(n10860), .B2(n10859), .A(n10858), .ZN(n10861) );
  AOI21_X1 U11498 ( .B1(n10863), .B2(n10862), .A(n10861), .ZN(n10864) );
  OAI21_X1 U11499 ( .B1(n10866), .B2(n10865), .A(n10864), .ZN(n10867) );
  AOI21_X1 U11500 ( .B1(n10869), .B2(n10868), .A(n10867), .ZN(n10936) );
  NOR2_X1 U11501 ( .A1(n10898), .A2(n5207), .ZN(n10870) );
  NOR2_X1 U11502 ( .A1(n10899), .A2(n5205), .ZN(n10902) );
  NOR2_X1 U11503 ( .A1(n10870), .A2(n10902), .ZN(n10872) );
  NOR2_X1 U11504 ( .A1(n10903), .A2(n5211), .ZN(n10871) );
  NOR2_X1 U11505 ( .A1(n10904), .A2(n5199), .ZN(n10907) );
  NOR2_X1 U11506 ( .A1(n10871), .A2(n10907), .ZN(n10910) );
  NAND2_X1 U11507 ( .A1(n10872), .A2(n10910), .ZN(n10912) );
  NOR2_X1 U11508 ( .A1(n10891), .A2(n5190), .ZN(n10873) );
  NOR2_X1 U11509 ( .A1(n9529), .A2(n5180), .ZN(n10894) );
  NOR2_X1 U11510 ( .A1(n10873), .A2(n10894), .ZN(n10897) );
  INV_X1 U11511 ( .A(n10968), .ZN(n10885) );
  NOR2_X1 U11512 ( .A1(n10886), .A2(n10885), .ZN(n10874) );
  NOR2_X1 U11513 ( .A1(n10887), .A2(n5186), .ZN(n10890) );
  NOR2_X1 U11514 ( .A1(n10874), .A2(n10890), .ZN(n10875) );
  NAND2_X1 U11515 ( .A1(n10897), .A2(n10875), .ZN(n10876) );
  NOR2_X1 U11516 ( .A1(n10912), .A2(n10876), .ZN(n10884) );
  NOR2_X1 U11517 ( .A1(n9886), .A2(n5161), .ZN(n10877) );
  NOR2_X1 U11518 ( .A1(n10914), .A2(n5159), .ZN(n10917) );
  NOR2_X1 U11519 ( .A1(n10877), .A2(n10917), .ZN(n10879) );
  NOR2_X1 U11520 ( .A1(n10918), .A2(n5155), .ZN(n10878) );
  NOR2_X1 U11521 ( .A1(n10919), .A2(n5151), .ZN(n10922) );
  NOR2_X1 U11522 ( .A1(n10878), .A2(n10922), .ZN(n10925) );
  NAND2_X1 U11523 ( .A1(n10879), .A2(n10925), .ZN(n10883) );
  NOR2_X1 U11524 ( .A1(n24), .A2(n5166), .ZN(n10880) );
  NOR2_X1 U11525 ( .A1(n10880), .A2(pmp_addr_i[158]), .ZN(n10882) );
  INV_X1 U11526 ( .A(pmp_addr_i[159]), .ZN(n10881) );
  NAND2_X1 U11527 ( .A1(n10882), .A2(n10881), .ZN(n10929) );
  NOR2_X1 U11528 ( .A1(n10883), .A2(n10929), .ZN(n10932) );
  NAND2_X1 U11529 ( .A1(n10884), .A2(n10932), .ZN(n10935) );
  NAND2_X1 U11530 ( .A1(n10886), .A2(n10885), .ZN(n10889) );
  NAND2_X1 U11531 ( .A1(n10887), .A2(n5186), .ZN(n10888) );
  OAI21_X1 U11532 ( .B1(n10890), .B2(n10889), .A(n10888), .ZN(n10896) );
  NAND2_X1 U11533 ( .A1(n10891), .A2(n5190), .ZN(n10893) );
  NAND2_X1 U11534 ( .A1(n11313), .A2(n5180), .ZN(n10892) );
  OAI21_X1 U11535 ( .B1(n10894), .B2(n10893), .A(n10892), .ZN(n10895) );
  AOI21_X1 U11536 ( .B1(n10897), .B2(n10896), .A(n10895), .ZN(n10913) );
  NAND2_X1 U11537 ( .A1(n10898), .A2(n5207), .ZN(n10901) );
  NAND2_X1 U11538 ( .A1(n10899), .A2(n5205), .ZN(n10900) );
  OAI21_X1 U11539 ( .B1(n10902), .B2(n10901), .A(n10900), .ZN(n10909) );
  NAND2_X1 U11540 ( .A1(n10903), .A2(n5211), .ZN(n10906) );
  NAND2_X1 U11541 ( .A1(n10904), .A2(n5199), .ZN(n10905) );
  OAI21_X1 U11542 ( .B1(n10907), .B2(n10906), .A(n10905), .ZN(n10908) );
  AOI21_X1 U11543 ( .B1(n10910), .B2(n10909), .A(n10908), .ZN(n10911) );
  OAI21_X1 U11544 ( .B1(n10913), .B2(n10912), .A(n10911), .ZN(n10933) );
  NAND2_X1 U11545 ( .A1(n11322), .A2(n5161), .ZN(n10916) );
  NAND2_X1 U11546 ( .A1(n10914), .A2(n5159), .ZN(n10915) );
  OAI21_X1 U11547 ( .B1(n10917), .B2(n10916), .A(n10915), .ZN(n10924) );
  NAND2_X1 U11548 ( .A1(n10918), .A2(n5155), .ZN(n10921) );
  NAND2_X1 U11549 ( .A1(n10919), .A2(n5151), .ZN(n10920) );
  OAI21_X1 U11550 ( .B1(n10922), .B2(n10921), .A(n10920), .ZN(n10923) );
  AOI21_X1 U11551 ( .B1(n10925), .B2(n10924), .A(n10923), .ZN(n10930) );
  NAND2_X1 U11552 ( .A1(n24), .A2(n5166), .ZN(n10926) );
  NOR2_X1 U11553 ( .A1(n10926), .A2(pmp_addr_i[158]), .ZN(n10927) );
  NAND2_X1 U11554 ( .A1(n10927), .A2(n10881), .ZN(n10928) );
  OAI21_X1 U11555 ( .B1(n10930), .B2(n10929), .A(n10928), .ZN(n10931) );
  AOI21_X1 U11556 ( .B1(n10933), .B2(n10932), .A(n10931), .ZN(n10934) );
  OAI21_X1 U11557 ( .B1(n10936), .B2(n10935), .A(n10934), .ZN(n10937) );
  NAND3_X1 U11558 ( .A1(n10938), .A2(n161), .A3(n10937), .ZN(n11023) );
  OAI22_X1 U11559 ( .A1(n10940), .A2(data_addr_o_9_), .B1(data_addr_o_12_), 
        .B2(n10939), .ZN(n10944) );
  OAI22_X1 U11560 ( .A1(n11343), .A2(n10942), .B1(n10836), .B2(n10941), .ZN(
        n10943) );
  OR2_X1 U11561 ( .A1(n10944), .A2(n10943), .ZN(n10951) );
  OAI22_X1 U11562 ( .A1(n10946), .A2(data_addr_o_11_), .B1(data_addr_o_14_), 
        .B2(n10945), .ZN(n10950) );
  OAI22_X1 U11563 ( .A1(n10948), .A2(n11309), .B1(n6649), .B2(n10947), .ZN(
        n10949) );
  NOR3_X1 U11564 ( .A1(n10951), .A2(n10950), .A3(n10949), .ZN(n10972) );
  OAI22_X1 U11565 ( .A1(n10954), .A2(n7816), .B1(n10953), .B2(n10952), .ZN(
        n10955) );
  INV_X1 U11566 ( .A(n10955), .ZN(n10962) );
  OAI22_X1 U11567 ( .A1(n10958), .A2(n10817), .B1(n10129), .B2(n10816), .ZN(
        n10959) );
  AOI21_X1 U11568 ( .B1(n10960), .B2(n12058), .A(n10959), .ZN(n10961) );
  OAI211_X1 U11569 ( .C1(n10963), .C2(n11255), .A(n10962), .B(n10961), .ZN(
        n10964) );
  AOI21_X1 U11570 ( .B1(n8444), .B2(n10965), .A(n10964), .ZN(n10971) );
  XNOR2_X1 U11571 ( .A(n11298), .B(n10966), .ZN(n10970) );
  XNOR2_X1 U11572 ( .A(n11283), .B(n10968), .ZN(n10969) );
  NAND4_X1 U11573 ( .A1(n10972), .A2(n10971), .A3(n10970), .A4(n10969), .ZN(
        n10978) );
  XNOR2_X1 U11574 ( .A(n10635), .B(n10973), .ZN(n10976) );
  XNOR2_X1 U11575 ( .A(data_addr_o_30_), .B(n10974), .ZN(n10975) );
  NAND2_X1 U11576 ( .A1(n10976), .A2(n10975), .ZN(n10977) );
  NOR2_X1 U11577 ( .A1(n10978), .A2(n10977), .ZN(n10998) );
  XNOR2_X1 U11578 ( .A(n11285), .B(n10979), .ZN(n10986) );
  XNOR2_X1 U11579 ( .A(n11312), .B(n10980), .ZN(n10985) );
  XNOR2_X1 U11580 ( .A(n11313), .B(n10981), .ZN(n10984) );
  XNOR2_X1 U11581 ( .A(data_addr_o_23_), .B(n10982), .ZN(n10983) );
  NAND4_X1 U11582 ( .A1(n10986), .A2(n10985), .A3(n10984), .A4(n10983), .ZN(
        n10996) );
  XNOR2_X1 U11583 ( .A(n10899), .B(n10987), .ZN(n10994) );
  XNOR2_X1 U11584 ( .A(n11320), .B(n10988), .ZN(n10993) );
  XNOR2_X1 U11585 ( .A(data_addr_o_26_), .B(n10989), .ZN(n10992) );
  XNOR2_X1 U11586 ( .A(n11322), .B(n10990), .ZN(n10991) );
  NAND4_X1 U11587 ( .A1(n10994), .A2(n10993), .A3(n10992), .A4(n10991), .ZN(
        n10995) );
  NOR2_X1 U11588 ( .A1(n10996), .A2(n10995), .ZN(n10997) );
  AND2_X1 U11589 ( .A1(n10998), .A2(n10997), .ZN(n11405) );
  AND2_X1 U11590 ( .A1(data_addr_o_17_), .A2(n10856), .ZN(n11369) );
  NAND4_X1 U11591 ( .A1(n11360), .A2(n11356), .A3(n11396), .A4(n11363), .ZN(
        n10999) );
  NOR2_X1 U11592 ( .A1(n11369), .A2(n10999), .ZN(n11011) );
  NAND2_X1 U11593 ( .A1(n11365), .A2(n11394), .ZN(n11003) );
  AOI21_X1 U11594 ( .B1(n11259), .B2(n10816), .A(pmp_cfg_i[43]), .ZN(n11000)
         );
  NAND2_X1 U11595 ( .A1(n22), .A2(n10817), .ZN(n11376) );
  AND3_X1 U11596 ( .A1(n11379), .A2(n11000), .A3(n11376), .ZN(n11001) );
  NAND4_X1 U11597 ( .A1(n11387), .A2(n11373), .A3(n11374), .A4(n11001), .ZN(
        n11002) );
  NOR2_X1 U11598 ( .A1(n11003), .A2(n11002), .ZN(n11010) );
  AND2_X1 U11599 ( .A1(n11004), .A2(n11015), .ZN(n11355) );
  OAI21_X1 U11600 ( .B1(n11006), .B2(n11005), .A(n11359), .ZN(n11371) );
  NOR2_X1 U11601 ( .A1(n11355), .A2(n11371), .ZN(n11009) );
  XNOR2_X1 U11602 ( .A(n12123), .B(n11007), .ZN(n11008) );
  NAND4_X1 U11603 ( .A1(n11011), .A2(n11010), .A3(n11009), .A4(n11008), .ZN(
        n11016) );
  XNOR2_X1 U11604 ( .A(n11303), .B(n11012), .ZN(n11013) );
  OAI21_X1 U11605 ( .B1(n11015), .B2(n11014), .A(n11013), .ZN(n11401) );
  NOR2_X1 U11606 ( .A1(n11016), .A2(n11401), .ZN(n11017) );
  NAND2_X1 U11607 ( .A1(n11405), .A2(n11017), .ZN(n11022) );
  OR2_X1 U11608 ( .A1(n11019), .A2(pmp_cfg_i[40]), .ZN(n11020) );
  OAI211_X1 U11609 ( .C1(pmp_cfg_i[41]), .C2(n11021), .A(n11018), .B(n11020), 
        .ZN(n11377) );
  AOI21_X1 U11610 ( .B1(n11023), .B2(n11022), .A(n11377), .ZN(n11024) );
  NOR2_X1 U11611 ( .A1(n11025), .A2(n11024), .ZN(n11026) );
  INV_X1 U11612 ( .A(n11030), .ZN(n11051) );
  NAND2_X1 U11613 ( .A1(n11032), .A2(n11031), .ZN(n11048) );
  INV_X1 U11614 ( .A(n11033), .ZN(n11041) );
  NAND2_X1 U11615 ( .A1(n7139), .A2(n11035), .ZN(n11036) );
  OAI211_X1 U11616 ( .C1(n11038), .C2(n11037), .A(n11036), .B(pmp_cfg_i[59]), 
        .ZN(n11039) );
  AOI21_X1 U11617 ( .B1(n11041), .B2(n11040), .A(n11039), .ZN(n11046) );
  INV_X1 U11618 ( .A(n11042), .ZN(n11044) );
  NAND2_X1 U11619 ( .A1(n11044), .A2(n11043), .ZN(n11045) );
  NAND4_X1 U11620 ( .A1(n11048), .A2(n11047), .A3(n11046), .A4(n11045), .ZN(
        n11049) );
  AOI21_X1 U11621 ( .B1(n11051), .B2(n11050), .A(n11049), .ZN(n11080) );
  NOR2_X1 U11622 ( .A1(n11054), .A2(n11052), .ZN(n11053) );
  MUX2_X1 U11623 ( .A(n11054), .B(n11053), .S(n9987), .Z(n11061) );
  INV_X1 U11624 ( .A(n11055), .ZN(n11058) );
  OAI22_X1 U11625 ( .A1(n11059), .A2(n11058), .B1(n11057), .B2(n11056), .ZN(
        n11060) );
  NOR2_X1 U11626 ( .A1(n11061), .A2(n11060), .ZN(n11079) );
  INV_X1 U11627 ( .A(n11062), .ZN(n11063) );
  OAI22_X1 U11628 ( .A1(n11066), .A2(n11065), .B1(n11064), .B2(n11063), .ZN(
        n11071) );
  OAI22_X1 U11629 ( .A1(n11069), .A2(n11068), .B1(n11067), .B2(pmp_addr_i[229]), .ZN(n11070) );
  NOR2_X1 U11630 ( .A1(n11071), .A2(n11070), .ZN(n11078) );
  AOI21_X1 U11631 ( .B1(n11074), .B2(n11073), .A(n11072), .ZN(n11075) );
  NAND2_X1 U11632 ( .A1(n11076), .A2(n11075), .ZN(n11077) );
  NAND4_X1 U11633 ( .A1(n11080), .A2(n11079), .A3(n11078), .A4(n11077), .ZN(
        n11081) );
  NOR2_X1 U11634 ( .A1(n11082), .A2(n11081), .ZN(n12091) );
  NAND2_X1 U11635 ( .A1(n12091), .A2(n12089), .ZN(n11354) );
  INV_X1 U11636 ( .A(n11083), .ZN(n11144) );
  INV_X1 U11637 ( .A(n11084), .ZN(n11088) );
  INV_X1 U11638 ( .A(n11085), .ZN(n11086) );
  AOI21_X1 U11639 ( .B1(n11088), .B2(n11087), .A(n11086), .ZN(n11089) );
  OAI21_X1 U11640 ( .B1(n11091), .B2(n11090), .A(n11089), .ZN(n11092) );
  AOI21_X1 U11641 ( .B1(n11094), .B2(n11093), .A(n11092), .ZN(n11132) );
  INV_X1 U11642 ( .A(n11095), .ZN(n11110) );
  NOR2_X1 U11643 ( .A1(n11097), .A2(pmp_addr_i[448]), .ZN(n11096) );
  MUX2_X1 U11644 ( .A(n11097), .B(n11096), .S(n10818), .Z(n11099) );
  NOR2_X1 U11645 ( .A1(n11099), .A2(n11098), .ZN(n11105) );
  OR2_X1 U11646 ( .A1(n11101), .A2(n11100), .ZN(n11102) );
  MUX2_X1 U11647 ( .A(n11103), .B(n11102), .S(n10479), .Z(n11104) );
  OAI211_X1 U11648 ( .C1(n11107), .C2(n11106), .A(n11105), .B(n11104), .ZN(
        n11108) );
  AOI21_X1 U11649 ( .B1(n11110), .B2(n11109), .A(n11108), .ZN(n11131) );
  OAI22_X1 U11650 ( .A1(n11114), .A2(n11113), .B1(n11112), .B2(n11111), .ZN(
        n11119) );
  INV_X1 U11651 ( .A(n11115), .ZN(n11116) );
  NOR2_X1 U11652 ( .A1(n11117), .A2(n11116), .ZN(n11118) );
  NOR2_X1 U11653 ( .A1(n11119), .A2(n11118), .ZN(n11130) );
  NAND2_X1 U11654 ( .A1(n11120), .A2(n11122), .ZN(n11121) );
  MUX2_X1 U11655 ( .A(n11122), .B(n11121), .S(n11255), .Z(n11123) );
  OAI21_X1 U11656 ( .B1(n11124), .B2(pmp_addr_i[454]), .A(n11123), .ZN(n11128)
         );
  NOR2_X1 U11657 ( .A1(n11126), .A2(n11125), .ZN(n11127) );
  NOR2_X1 U11658 ( .A1(n11128), .A2(n11127), .ZN(n11129) );
  NAND4_X1 U11659 ( .A1(n11132), .A2(n11131), .A3(n11130), .A4(n11129), .ZN(
        n11142) );
  NOR2_X1 U11660 ( .A1(n11134), .A2(n11133), .ZN(n11137) );
  OAI21_X1 U11661 ( .B1(n11137), .B2(n7841), .A(n11136), .ZN(n11141) );
  MUX2_X1 U11662 ( .A(n11139), .B(n11138), .S(n9987), .Z(n11140) );
  NOR3_X1 U11663 ( .A1(n11142), .A2(n11141), .A3(n11140), .ZN(n11143) );
  NAND2_X1 U11664 ( .A1(n11144), .A2(n11143), .ZN(n12079) );
  INV_X1 U11665 ( .A(n12079), .ZN(n11146) );
  NAND2_X1 U11666 ( .A1(n11146), .A2(n11145), .ZN(n11353) );
  INV_X1 U11668 ( .A(n11148), .ZN(n11172) );
  INV_X1 U11669 ( .A(n11149), .ZN(n11163) );
  INV_X1 U11670 ( .A(n11151), .ZN(n11160) );
  INV_X1 U11671 ( .A(pmp_addr_i[64]), .ZN(n11153) );
  NAND2_X1 U11672 ( .A1(n6254), .A2(n11153), .ZN(n11159) );
  INV_X1 U11673 ( .A(n11154), .ZN(n11157) );
  INV_X1 U11674 ( .A(n11155), .ZN(n11156) );
  NOR2_X1 U11675 ( .A1(n11157), .A2(n11156), .ZN(n11158) );
  OAI211_X1 U11676 ( .C1(n6259), .C2(n11160), .A(n11159), .B(n11158), .ZN(
        n11161) );
  AOI21_X1 U11677 ( .B1(n11163), .B2(n11162), .A(n11161), .ZN(n11170) );
  OAI21_X1 U11678 ( .B1(n11166), .B2(n11165), .A(n11164), .ZN(n11168) );
  NAND2_X1 U11679 ( .A1(n11168), .A2(n11167), .ZN(n11169) );
  OAI211_X1 U11680 ( .C1(n11172), .C2(n11171), .A(n11170), .B(n11169), .ZN(
        n11182) );
  OAI22_X1 U11681 ( .A1(n11176), .A2(n11175), .B1(n11174), .B2(n11173), .ZN(
        n11181) );
  OAI22_X1 U11682 ( .A1(n11179), .A2(pmp_addr_i[73]), .B1(n11178), .B2(n11177), 
        .ZN(n11180) );
  NOR3_X1 U11683 ( .A1(n11182), .A2(n11181), .A3(n11180), .ZN(n11202) );
  MUX2_X1 U11684 ( .A(n11184), .B(n11183), .S(n9066), .Z(n11189) );
  OAI21_X1 U11685 ( .B1(n11185), .B2(n2056), .A(n11187), .ZN(n11186) );
  MUX2_X1 U11686 ( .A(n11187), .B(n11186), .S(n11309), .Z(n11188) );
  NAND2_X1 U11687 ( .A1(n11189), .A2(n11188), .ZN(n11190) );
  AOI21_X1 U11688 ( .B1(n11192), .B2(n11191), .A(n11190), .ZN(n11201) );
  AND2_X1 U11689 ( .A1(n11194), .A2(n11193), .ZN(n11195) );
  MUX2_X1 U11690 ( .A(n11196), .B(n11195), .S(n9987), .Z(n11197) );
  AOI21_X1 U11691 ( .B1(n11199), .B2(n11198), .A(n11197), .ZN(n11200) );
  NAND4_X1 U11692 ( .A1(n12230), .A2(n11202), .A3(n11201), .A4(n11200), .ZN(
        n12072) );
  INV_X1 U11693 ( .A(n12072), .ZN(n11205) );
  NAND2_X1 U11694 ( .A1(n11205), .A2(n11204), .ZN(n11352) );
  AND2_X1 U11695 ( .A1(data_addr_o_9_), .A2(n158), .ZN(n11243) );
  AND2_X1 U11696 ( .A1(data_addr_o_11_), .A2(n11335), .ZN(n11268) );
  AOI22_X1 U11697 ( .A1(n11243), .A2(n11207), .B1(n11268), .B2(n11206), .ZN(
        n11224) );
  AND2_X1 U11698 ( .A1(data_addr_o_14_), .A2(n11208), .ZN(n11269) );
  INV_X1 U11699 ( .A(n11209), .ZN(n11212) );
  AND2_X1 U11700 ( .A1(n10499), .A2(n11336), .ZN(n11244) );
  INV_X1 U11701 ( .A(n11210), .ZN(n11211) );
  AOI22_X1 U11702 ( .A1(n11269), .A2(n11212), .B1(n11244), .B2(n11211), .ZN(
        n11223) );
  INV_X1 U11703 ( .A(n11213), .ZN(n11342) );
  AND2_X1 U11704 ( .A1(data_addr_o_10_), .A2(n11342), .ZN(n11242) );
  INV_X1 U11705 ( .A(n11214), .ZN(n11216) );
  AND2_X1 U11706 ( .A1(data_addr_i[13]), .A2(n330), .ZN(n11267) );
  AOI22_X1 U11707 ( .A1(n11242), .A2(n11216), .B1(n11267), .B2(n11215), .ZN(
        n11222) );
  AND2_X1 U11708 ( .A1(n9805), .A2(n159), .ZN(n11245) );
  AND2_X1 U11709 ( .A1(data_addr_o_7_), .A2(n11345), .ZN(n11256) );
  INV_X1 U11710 ( .A(n11218), .ZN(n11219) );
  AOI22_X1 U11711 ( .A1(n11245), .A2(n11220), .B1(n11256), .B2(n11219), .ZN(
        n11221) );
  NAND4_X1 U11712 ( .A1(n11224), .A2(n11223), .A3(n11222), .A4(n11221), .ZN(
        n11281) );
  INV_X1 U11713 ( .A(n11225), .ZN(n11275) );
  AND2_X1 U11714 ( .A1(data_addr_o_16_), .A2(n328), .ZN(n11274) );
  NAND2_X1 U11715 ( .A1(n11274), .A2(n11226), .ZN(n11240) );
  NAND2_X1 U11716 ( .A1(n11227), .A2(n329), .ZN(n11271) );
  INV_X1 U11717 ( .A(n11228), .ZN(n11286) );
  NAND2_X1 U11718 ( .A1(data_addr_o_3_), .A2(n11286), .ZN(n11252) );
  NAND2_X1 U11719 ( .A1(data_addr_o_4_), .A2(n11229), .ZN(n11231) );
  OAI211_X1 U11720 ( .C1(n11252), .C2(pmp_addr_i[0]), .A(n11231), .B(n11230), 
        .ZN(n11232) );
  AOI21_X1 U11721 ( .B1(n11233), .B2(data_addr_o_5_), .A(n11232), .ZN(n11236)
         );
  AND2_X1 U11722 ( .A1(data_addr_o_6_), .A2(n324), .ZN(n11257) );
  NAND2_X1 U11723 ( .A1(n11257), .A2(n11234), .ZN(n11235) );
  OAI211_X1 U11724 ( .C1(n11271), .C2(n11237), .A(n11236), .B(n11235), .ZN(
        n11238) );
  INV_X1 U11725 ( .A(n11238), .ZN(n11239) );
  OAI211_X1 U11726 ( .C1(n11241), .C2(n11275), .A(n11240), .B(n11239), .ZN(
        n11280) );
  INV_X1 U11727 ( .A(n11242), .ZN(n11249) );
  INV_X1 U11728 ( .A(n11243), .ZN(n11248) );
  INV_X1 U11729 ( .A(n11244), .ZN(n11247) );
  INV_X1 U11730 ( .A(n11245), .ZN(n11246) );
  NAND4_X1 U11731 ( .A1(n11249), .A2(n11248), .A3(n11247), .A4(n11246), .ZN(
        n11266) );
  INV_X1 U11732 ( .A(n11250), .ZN(n11251) );
  NAND2_X1 U11733 ( .A1(n11252), .A2(n11251), .ZN(n11253) );
  AOI21_X1 U11734 ( .B1(n11255), .B2(n11254), .A(n11253), .ZN(n11264) );
  INV_X1 U11735 ( .A(n11256), .ZN(n11263) );
  INV_X1 U11736 ( .A(n11257), .ZN(n11262) );
  XNOR2_X1 U11737 ( .A(n11259), .B(n11258), .ZN(n11260) );
  AOI21_X1 U11738 ( .B1(n10135), .B2(n11287), .A(n11260), .ZN(n11261) );
  NAND4_X1 U11739 ( .A1(n11264), .A2(n11263), .A3(n11262), .A4(n11261), .ZN(
        n11265) );
  NOR2_X1 U11740 ( .A1(n11266), .A2(n11265), .ZN(n11278) );
  INV_X1 U11741 ( .A(n11267), .ZN(n11273) );
  INV_X1 U11742 ( .A(n11268), .ZN(n11272) );
  INV_X1 U11743 ( .A(n11269), .ZN(n11270) );
  AND4_X1 U11744 ( .A1(n11273), .A2(n11272), .A3(n11271), .A4(n11270), .ZN(
        n11277) );
  INV_X1 U11745 ( .A(n11274), .ZN(n11276) );
  NAND4_X1 U11746 ( .A1(n11278), .A2(n11277), .A3(n11276), .A4(n11275), .ZN(
        n11279) );
  OAI21_X1 U11747 ( .B1(n11281), .B2(n11280), .A(n11279), .ZN(n11302) );
  XNOR2_X1 U11748 ( .A(n11283), .B(n11282), .ZN(n11294) );
  XNOR2_X1 U11749 ( .A(n11285), .B(n11284), .ZN(n11293) );
  OAI22_X1 U11750 ( .A1(n11288), .A2(n11287), .B1(n10130), .B2(n11286), .ZN(
        n11289) );
  AOI21_X1 U11751 ( .B1(n11291), .B2(n11290), .A(n11289), .ZN(n11292) );
  AND3_X1 U11752 ( .A1(n11294), .A2(n11293), .A3(n11292), .ZN(n11301) );
  XNOR2_X1 U11753 ( .A(data_addr_o_23_), .B(n11295), .ZN(n11300) );
  XNOR2_X1 U11754 ( .A(n11298), .B(n11297), .ZN(n11299) );
  NAND4_X1 U11755 ( .A1(n11302), .A2(n11301), .A3(n11300), .A4(n11299), .ZN(
        n12083) );
  INV_X1 U11756 ( .A(n12083), .ZN(n11350) );
  XNOR2_X1 U11757 ( .A(n11303), .B(pmp_addr_i[27]), .ZN(n11307) );
  XNOR2_X1 U11758 ( .A(data_addr_o_30_), .B(n11304), .ZN(n11306) );
  AND2_X1 U11759 ( .A1(n11307), .A2(n11306), .ZN(n11317) );
  INV_X1 U11760 ( .A(n11308), .ZN(n11311) );
  OAI22_X1 U11761 ( .A1(n9987), .A2(n328), .B1(n11309), .B2(n329), .ZN(n11310)
         );
  NOR2_X1 U11762 ( .A1(n11311), .A2(n11310), .ZN(n11316) );
  XNOR2_X1 U11763 ( .A(n11312), .B(pmp_addr_i[19]), .ZN(n11315) );
  XNOR2_X1 U11764 ( .A(n11313), .B(pmp_addr_i[20]), .ZN(n11314) );
  NAND4_X1 U11765 ( .A1(n11317), .A2(n11316), .A3(n11315), .A4(n11314), .ZN(
        n11328) );
  XNOR2_X1 U11766 ( .A(n10635), .B(n11318), .ZN(n11326) );
  XNOR2_X1 U11767 ( .A(n11320), .B(pmp_addr_i[23]), .ZN(n11325) );
  XNOR2_X1 U11768 ( .A(n11322), .B(n11321), .ZN(n11324) );
  XNOR2_X1 U11769 ( .A(n10738), .B(pmp_addr_i[22]), .ZN(n11323) );
  NAND4_X1 U11770 ( .A1(n11326), .A2(n11325), .A3(n11324), .A4(n11323), .ZN(
        n11327) );
  NOR2_X1 U11771 ( .A1(n11328), .A2(n11327), .ZN(n12082) );
  XNOR2_X1 U11772 ( .A(data_addr_o_26_), .B(pmp_addr_i[24]), .ZN(n11341) );
  OAI21_X1 U11773 ( .B1(n11331), .B2(n324), .A(n11330), .ZN(n11332) );
  AOI21_X1 U11774 ( .B1(n11334), .B2(n11333), .A(n11332), .ZN(n11340) );
  OAI22_X1 U11775 ( .A1(data_addr_o_11_), .A2(n11335), .B1(n8237), .B2(n158), 
        .ZN(n11338) );
  OAI22_X1 U11776 ( .A1(data_addr_o_12_), .A2(n11336), .B1(data_addr_o_13_), 
        .B2(n330), .ZN(n11337) );
  NOR2_X1 U11777 ( .A1(n11338), .A2(n11337), .ZN(n11339) );
  AND3_X1 U11778 ( .A1(n11341), .A2(n11340), .A3(n11339), .ZN(n12081) );
  OAI22_X1 U11779 ( .A1(n11343), .A2(n11342), .B1(n9805), .B2(n159), .ZN(
        n11347) );
  OAI21_X1 U11780 ( .B1(n7816), .B2(n11345), .A(n3758), .ZN(n11346) );
  NOR2_X1 U11781 ( .A1(n11347), .A2(n11346), .ZN(n12080) );
  INV_X1 U11782 ( .A(n12080), .ZN(n11348) );
  NOR2_X1 U11783 ( .A1(n11348), .A2(pmp_addr_i[29]), .ZN(n11349) );
  NAND4_X1 U11784 ( .A1(n11350), .A2(n12082), .A3(n12081), .A4(n11349), .ZN(
        n11351) );
  AND4_X1 U11785 ( .A1(n11352), .A2(n11353), .A3(n11354), .A4(n11351), .ZN(
        n11581) );
  OAI22_X1 U11786 ( .A1(n10854), .A2(n11358), .B1(n11357), .B2(n11356), .ZN(
        n11368) );
  OAI22_X1 U11787 ( .A1(n11361), .A2(n11360), .B1(n11359), .B2(pmp_addr_i[171]), .ZN(n11367) );
  OAI22_X1 U11788 ( .A1(n11365), .A2(n11364), .B1(n11363), .B2(n11362), .ZN(
        n11366) );
  NOR3_X1 U11789 ( .A1(n11368), .A2(n11367), .A3(n11366), .ZN(n11404) );
  NAND2_X1 U11790 ( .A1(n11371), .A2(n11370), .ZN(n11391) );
  OAI22_X1 U11791 ( .A1(n11375), .A2(n11374), .B1(n11373), .B2(n11372), .ZN(
        n11389) );
  INV_X1 U11792 ( .A(pmp_addr_i[160]), .ZN(n11378) );
  AOI21_X1 U11793 ( .B1(n10819), .B2(n11378), .A(n11377), .ZN(n11385) );
  INV_X1 U11794 ( .A(n11379), .ZN(n11383) );
  OAI22_X1 U11795 ( .A1(n11383), .A2(n11382), .B1(n11381), .B2(n11380), .ZN(
        n11384) );
  OAI211_X1 U11796 ( .C1(n11387), .C2(n11386), .A(n11385), .B(n11384), .ZN(
        n11388) );
  NOR2_X1 U11797 ( .A1(n11389), .A2(n11388), .ZN(n11390) );
  OAI211_X1 U11798 ( .C1(n10859), .C2(n11392), .A(n11391), .B(n11390), .ZN(
        n11393) );
  INV_X1 U11799 ( .A(n11393), .ZN(n11403) );
  NOR2_X1 U11800 ( .A1(n11395), .A2(n11394), .ZN(n11400) );
  INV_X1 U11801 ( .A(n11396), .ZN(n11398) );
  AND2_X1 U11802 ( .A1(n11398), .A2(n11397), .ZN(n11399) );
  NOR3_X1 U11803 ( .A1(n11401), .A2(n11400), .A3(n11399), .ZN(n11402) );
  NAND4_X1 U11804 ( .A1(n11405), .A2(n11404), .A3(n11403), .A4(n11402), .ZN(
        n12074) );
  INV_X1 U11805 ( .A(n12074), .ZN(n11462) );
  INV_X1 U11806 ( .A(n11406), .ZN(n11407) );
  OAI22_X1 U11807 ( .A1(n9987), .A2(n11409), .B1(n11408), .B2(n11407), .ZN(
        n11416) );
  INV_X1 U11808 ( .A(n11410), .ZN(n11414) );
  OAI22_X1 U11809 ( .A1(n11414), .A2(n11413), .B1(n11412), .B2(n11411), .ZN(
        n11415) );
  OR2_X1 U11810 ( .A1(n11416), .A2(n11415), .ZN(n11441) );
  INV_X1 U11811 ( .A(n11418), .ZN(n11424) );
  INV_X1 U11812 ( .A(n11419), .ZN(n11422) );
  INV_X1 U11813 ( .A(n11420), .ZN(n11421) );
  AOI22_X1 U11814 ( .A1(n11424), .A2(n11423), .B1(n11422), .B2(n11421), .ZN(
        n11433) );
  NOR2_X1 U11815 ( .A1(n11426), .A2(n11425), .ZN(n11431) );
  INV_X1 U11816 ( .A(n11427), .ZN(n11428) );
  OAI211_X1 U11817 ( .C1(n11429), .C2(pmp_addr_i[384]), .A(pmp_cfg_i[99]), .B(
        n11428), .ZN(n11430) );
  NOR2_X1 U11818 ( .A1(n11431), .A2(n11430), .ZN(n11432) );
  OAI211_X1 U11819 ( .C1(n11434), .C2(n8535), .A(n11433), .B(n11432), .ZN(
        n11440) );
  OAI22_X1 U11820 ( .A1(n11438), .A2(n11437), .B1(n11436), .B2(n11435), .ZN(
        n11439) );
  NOR3_X1 U11821 ( .A1(n11441), .A2(n11440), .A3(n11439), .ZN(n11457) );
  INV_X1 U11822 ( .A(n11442), .ZN(n11445) );
  OAI21_X1 U11823 ( .B1(n11445), .B2(n11444), .A(n11443), .ZN(n11447) );
  AOI22_X1 U11824 ( .A1(n11449), .A2(n11448), .B1(n11447), .B2(n11446), .ZN(
        n11456) );
  NAND2_X1 U11825 ( .A1(n11451), .A2(n11450), .ZN(n11452) );
  NAND3_X1 U11826 ( .A1(n11454), .A2(n11453), .A3(n11452), .ZN(n11455) );
  NAND4_X1 U11827 ( .A1(n11458), .A2(n11457), .A3(n11456), .A4(n11455), .ZN(
        n12086) );
  INV_X1 U11828 ( .A(n12086), .ZN(n11460) );
  AOI22_X1 U11829 ( .A1(n11462), .A2(n11461), .B1(n11460), .B2(n11459), .ZN(
        n11580) );
  INV_X1 U11830 ( .A(n11464), .ZN(n11467) );
  INV_X1 U11831 ( .A(n11465), .ZN(n11466) );
  NAND2_X1 U11832 ( .A1(n11467), .A2(n11466), .ZN(n11472) );
  INV_X1 U11833 ( .A(n11468), .ZN(n11470) );
  NAND2_X1 U11834 ( .A1(n11470), .A2(n11469), .ZN(n11471) );
  OAI211_X1 U11835 ( .C1(n8252), .C2(n11473), .A(n11472), .B(n11471), .ZN(
        n11499) );
  INV_X1 U11836 ( .A(n11474), .ZN(n11480) );
  INV_X1 U11837 ( .A(n11475), .ZN(n11478) );
  INV_X1 U11838 ( .A(n11476), .ZN(n11477) );
  AOI22_X1 U11839 ( .A1(n11480), .A2(n11479), .B1(n11478), .B2(n11477), .ZN(
        n11490) );
  NAND2_X1 U11840 ( .A1(n8217), .A2(n11482), .ZN(n11483) );
  OAI211_X1 U11841 ( .C1(n11485), .C2(n11484), .A(n11483), .B(pmp_cfg_i[11]), 
        .ZN(n11486) );
  AOI21_X1 U11842 ( .B1(n11488), .B2(n11487), .A(n11486), .ZN(n11489) );
  OAI211_X1 U11843 ( .C1(n11492), .C2(n11491), .A(n11490), .B(n11489), .ZN(
        n11498) );
  INV_X1 U11844 ( .A(n11493), .ZN(n11496) );
  OAI22_X1 U11845 ( .A1(n11496), .A2(n11495), .B1(n11494), .B2(pmp_addr_i[38]), 
        .ZN(n11497) );
  NOR3_X1 U11846 ( .A1(n11499), .A2(n11498), .A3(n11497), .ZN(n11516) );
  INV_X1 U11847 ( .A(n11500), .ZN(n11511) );
  INV_X1 U11848 ( .A(n11501), .ZN(n11503) );
  NAND2_X1 U11849 ( .A1(n11503), .A2(n11502), .ZN(n11506) );
  INV_X1 U11850 ( .A(n11504), .ZN(n11505) );
  OAI211_X1 U11851 ( .C1(n11508), .C2(n11507), .A(n11506), .B(n11505), .ZN(
        n11509) );
  AOI21_X1 U11852 ( .B1(n11511), .B2(n11510), .A(n11509), .ZN(n11515) );
  NAND2_X1 U11853 ( .A1(n11513), .A2(n11512), .ZN(n11514) );
  NAND4_X1 U11854 ( .A1(n11517), .A2(n11516), .A3(n11515), .A4(n11514), .ZN(
        n12076) );
  INV_X1 U11855 ( .A(n12076), .ZN(n11518) );
  NAND2_X1 U11856 ( .A1(n11518), .A2(n12075), .ZN(n11579) );
  INV_X1 U11858 ( .A(n11520), .ZN(n11525) );
  INV_X1 U11859 ( .A(n11521), .ZN(n11524) );
  AOI22_X1 U11860 ( .A1(n11525), .A2(n11524), .B1(n11523), .B2(n11522), .ZN(
        n11558) );
  INV_X1 U11861 ( .A(n11526), .ZN(n11528) );
  OAI21_X1 U11862 ( .B1(n11529), .B2(n11528), .A(n11527), .ZN(n11532) );
  INV_X1 U11863 ( .A(n11530), .ZN(n11531) );
  NAND2_X1 U11864 ( .A1(n11532), .A2(n11531), .ZN(n11557) );
  INV_X1 U11865 ( .A(n11533), .ZN(n11542) );
  NAND2_X1 U11866 ( .A1(n10487), .A2(n11535), .ZN(n11540) );
  OAI21_X1 U11867 ( .B1(n11537), .B2(pmp_addr_i[192]), .A(pmp_cfg_i[51]), .ZN(
        n11538) );
  AOI21_X1 U11868 ( .B1(n10480), .B2(n651), .A(n11538), .ZN(n11539) );
  OAI211_X1 U11869 ( .C1(n11542), .C2(n11541), .A(n11540), .B(n11539), .ZN(
        n11551) );
  INV_X1 U11870 ( .A(n11543), .ZN(n11548) );
  INV_X1 U11871 ( .A(n11544), .ZN(n11546) );
  OAI22_X1 U11872 ( .A1(n11548), .A2(n11547), .B1(n11546), .B2(n11545), .ZN(
        n11550) );
  NOR3_X1 U11873 ( .A1(n11551), .A2(n11550), .A3(n11549), .ZN(n11556) );
  INV_X1 U11874 ( .A(n11552), .ZN(n11554) );
  NAND2_X1 U11875 ( .A1(n11554), .A2(n11553), .ZN(n11555) );
  AND4_X1 U11876 ( .A1(n11558), .A2(n11557), .A3(n11556), .A4(n11555), .ZN(
        n11575) );
  INV_X1 U11877 ( .A(n11559), .ZN(n11565) );
  INV_X1 U11878 ( .A(n11560), .ZN(n11563) );
  INV_X1 U11879 ( .A(n11561), .ZN(n11562) );
  AOI22_X1 U11880 ( .A1(n11565), .A2(n11564), .B1(n11563), .B2(n11562), .ZN(
        n11573) );
  INV_X1 U11881 ( .A(n11566), .ZN(n11571) );
  MUX2_X1 U11882 ( .A(n11568), .B(n11567), .S(n11004), .Z(n11569) );
  AOI21_X1 U11883 ( .B1(n11571), .B2(n11570), .A(n11569), .ZN(n11572) );
  NAND4_X1 U11884 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11576) );
  NOR2_X1 U11885 ( .A1(n11577), .A2(n11576), .ZN(n12094) );
  OAI22_X1 U11889 ( .A1(n11585), .A2(n11584), .B1(n8877), .B2(n11583), .ZN(
        n11593) );
  INV_X1 U11890 ( .A(n11586), .ZN(n11591) );
  INV_X1 U11891 ( .A(n11587), .ZN(n11588) );
  OAI22_X1 U11892 ( .A1(n11591), .A2(n11590), .B1(n11589), .B2(n11588), .ZN(
        n11592) );
  NOR2_X1 U11893 ( .A1(n11593), .A2(n11592), .ZN(n11612) );
  INV_X1 U11894 ( .A(n11594), .ZN(n11604) );
  INV_X1 U11895 ( .A(n11595), .ZN(n11597) );
  OAI211_X1 U11896 ( .C1(n11598), .C2(pmp_addr_i[256]), .A(n11597), .B(n11596), 
        .ZN(n11599) );
  INV_X1 U11897 ( .A(n11599), .ZN(n11600) );
  OAI21_X1 U11898 ( .B1(n11601), .B2(pmp_addr_i[259]), .A(n11600), .ZN(n11602)
         );
  AOI21_X1 U11899 ( .B1(n11604), .B2(n11603), .A(n11602), .ZN(n11611) );
  INV_X1 U11900 ( .A(n11605), .ZN(n11606) );
  OR2_X1 U11901 ( .A1(n11607), .A2(n11606), .ZN(n11608) );
  MUX2_X1 U11902 ( .A(n11609), .B(n11608), .S(n11014), .Z(n11610) );
  NAND3_X1 U11903 ( .A1(n11612), .A2(n11611), .A3(n11610), .ZN(n11630) );
  INV_X1 U11904 ( .A(n11613), .ZN(n11625) );
  INV_X1 U11905 ( .A(n11614), .ZN(n11619) );
  INV_X1 U11906 ( .A(n11615), .ZN(n11617) );
  AOI22_X1 U11907 ( .A1(n11619), .A2(n11618), .B1(n11617), .B2(n11616), .ZN(
        n11623) );
  NAND2_X1 U11908 ( .A1(n11621), .A2(n11620), .ZN(n11622) );
  OAI211_X1 U11909 ( .C1(n11625), .C2(n11624), .A(n11623), .B(n11622), .ZN(
        n11629) );
  NOR2_X1 U11910 ( .A1(n11627), .A2(n11626), .ZN(n11628) );
  NOR3_X1 U11911 ( .A1(n11630), .A2(n11629), .A3(n11628), .ZN(n11638) );
  INV_X1 U11912 ( .A(n11631), .ZN(n11632) );
  NAND2_X1 U11913 ( .A1(n11633), .A2(n11632), .ZN(n11637) );
  OR2_X1 U11914 ( .A1(n11635), .A2(n11634), .ZN(n11636) );
  NAND4_X1 U11915 ( .A1(n11639), .A2(n11638), .A3(n11637), .A4(n11636), .ZN(
        n12112) );
  INV_X1 U11916 ( .A(n11640), .ZN(n11645) );
  INV_X1 U11917 ( .A(n11641), .ZN(n11643) );
  AOI22_X1 U11918 ( .A1(n11645), .A2(n11644), .B1(n11643), .B2(n11642), .ZN(
        n11673) );
  INV_X1 U11919 ( .A(n11646), .ZN(n11651) );
  INV_X1 U11920 ( .A(n11647), .ZN(n11649) );
  AOI22_X1 U11921 ( .A1(n11651), .A2(n11650), .B1(n11649), .B2(n11648), .ZN(
        n11672) );
  INV_X1 U11922 ( .A(n11652), .ZN(n11656) );
  AOI22_X1 U11923 ( .A1(n11656), .A2(n11655), .B1(n11654), .B2(n11653), .ZN(
        n11671) );
  INV_X1 U11924 ( .A(n11657), .ZN(n11669) );
  INV_X1 U11925 ( .A(pmp_addr_i[320]), .ZN(n11660) );
  AOI21_X1 U11926 ( .B1(n9214), .B2(n11660), .A(n11659), .ZN(n11665) );
  INV_X1 U11927 ( .A(n11661), .ZN(n11663) );
  NAND2_X1 U11928 ( .A1(n11663), .A2(n11662), .ZN(n11664) );
  OAI211_X1 U11929 ( .C1(n11666), .C2(pmp_addr_i[323]), .A(n11665), .B(n11664), 
        .ZN(n11667) );
  AOI21_X1 U11930 ( .B1(n11669), .B2(n11668), .A(n11667), .ZN(n11670) );
  AND4_X1 U11931 ( .A1(n11673), .A2(n11672), .A3(n11671), .A4(n11670), .ZN(
        n11694) );
  INV_X1 U11932 ( .A(n11674), .ZN(n11675) );
  NAND2_X1 U11933 ( .A1(n11675), .A2(n11676), .ZN(n11679) );
  INV_X1 U11934 ( .A(n11676), .ZN(n11677) );
  AOI22_X1 U11935 ( .A1(n11679), .A2(n11678), .B1(pmp_addr_i[329]), .B2(n11677), .ZN(n11683) );
  MUX2_X1 U11936 ( .A(n11681), .B(n11680), .S(data_addr_o_16_), .Z(n11682) );
  NOR2_X1 U11937 ( .A1(n11683), .A2(n11682), .ZN(n11693) );
  INV_X1 U11938 ( .A(n11684), .ZN(n11685) );
  AOI21_X1 U11939 ( .B1(n11687), .B2(n11686), .A(n11685), .ZN(n11692) );
  INV_X1 U11940 ( .A(n11688), .ZN(n11690) );
  NAND2_X1 U11941 ( .A1(n11690), .A2(n11689), .ZN(n11691) );
  NAND4_X1 U11942 ( .A1(n11694), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(
        n11695) );
  NOR2_X1 U11943 ( .A1(n11696), .A2(n11695), .ZN(n12101) );
  INV_X1 U11944 ( .A(n11697), .ZN(n11757) );
  INV_X1 U11945 ( .A(n11699), .ZN(n11705) );
  INV_X1 U11946 ( .A(n11700), .ZN(n11703) );
  INV_X1 U11947 ( .A(n11701), .ZN(n11702) );
  AOI22_X1 U11948 ( .A1(n11705), .A2(n11704), .B1(n11703), .B2(n11702), .ZN(
        n11706) );
  OAI21_X1 U11949 ( .B1(n11707), .B2(n7370), .A(n11706), .ZN(n11721) );
  INV_X1 U11950 ( .A(n11708), .ZN(n11718) );
  INV_X1 U11951 ( .A(n11709), .ZN(n11711) );
  NAND2_X1 U11952 ( .A1(n11711), .A2(n11710), .ZN(n11717) );
  INV_X1 U11953 ( .A(n11712), .ZN(n11715) );
  INV_X1 U11954 ( .A(n11713), .ZN(n11714) );
  NAND2_X1 U11955 ( .A1(n11715), .A2(n11714), .ZN(n11716) );
  OAI211_X1 U11956 ( .C1(n11719), .C2(n11718), .A(n11717), .B(n11716), .ZN(
        n11720) );
  NOR2_X1 U11957 ( .A1(n11721), .A2(n11720), .ZN(n11755) );
  OR2_X1 U11958 ( .A1(n11723), .A2(n11722), .ZN(n11741) );
  INV_X1 U11959 ( .A(n11724), .ZN(n11731) );
  OAI21_X1 U11960 ( .B1(n11727), .B2(n11726), .A(n11725), .ZN(n11729) );
  AOI22_X1 U11961 ( .A1(n11731), .A2(n11730), .B1(n11729), .B2(n11728), .ZN(
        n11740) );
  INV_X1 U11962 ( .A(n11732), .ZN(n11737) );
  OAI21_X1 U11963 ( .B1(n11734), .B2(pmp_addr_i[96]), .A(n11733), .ZN(n11735)
         );
  AOI21_X1 U11964 ( .B1(n11737), .B2(n11736), .A(n11735), .ZN(n11738) );
  NAND4_X1 U11965 ( .A1(n11741), .A2(n11740), .A3(n11739), .A4(n11738), .ZN(
        n11744) );
  INV_X1 U11966 ( .A(n11742), .ZN(n11743) );
  NOR2_X1 U11967 ( .A1(n11744), .A2(n11743), .ZN(n11754) );
  OR2_X1 U11968 ( .A1(n11746), .A2(n11745), .ZN(n11753) );
  OAI21_X1 U11969 ( .B1(n11749), .B2(n11748), .A(n11747), .ZN(n11750) );
  NAND2_X1 U11970 ( .A1(n11751), .A2(n11750), .ZN(n11752) );
  NAND4_X1 U11971 ( .A1(n11755), .A2(n11754), .A3(n11753), .A4(n11752), .ZN(
        n11756) );
  NOR2_X1 U11972 ( .A1(n11757), .A2(n11756), .ZN(n12102) );
  AOI22_X1 U11975 ( .A1(n11763), .A2(n11762), .B1(n6536), .B2(n11761), .ZN(
        n11774) );
  INV_X1 U11976 ( .A(n11764), .ZN(n11768) );
  INV_X1 U11977 ( .A(n11765), .ZN(n11767) );
  AOI22_X1 U11978 ( .A1(n11768), .A2(n11767), .B1(n6507), .B2(n3877), .ZN(
        n11772) );
  NAND2_X1 U11979 ( .A1(n11770), .A2(n11769), .ZN(n11771) );
  NAND4_X1 U11980 ( .A1(n11774), .A2(n11773), .A3(n11772), .A4(n11771), .ZN(
        n11775) );
  NOR2_X1 U11981 ( .A1(n11776), .A2(n11775), .ZN(n12108) );
  INV_X1 U11982 ( .A(n11778), .ZN(n11780) );
  AOI22_X1 U11983 ( .A1(n6540), .A2(n11781), .B1(n11780), .B2(n11779), .ZN(
        n11787) );
  AOI22_X1 U11984 ( .A1(n6512), .A2(n11785), .B1(n6513), .B2(n11784), .ZN(
        n11786) );
  OAI211_X1 U11985 ( .C1(n11789), .C2(n11788), .A(n11787), .B(n11786), .ZN(
        n11795) );
  INV_X1 U11986 ( .A(n11790), .ZN(n11791) );
  NAND2_X1 U11987 ( .A1(data_addr_o_17_), .A2(n11791), .ZN(n11792) );
  NOR2_X1 U11988 ( .A1(n11793), .A2(n11792), .ZN(n11794) );
  NOR2_X1 U11989 ( .A1(n11795), .A2(n11794), .ZN(n12107) );
  INV_X1 U11990 ( .A(n11796), .ZN(n11797) );
  OAI21_X1 U11991 ( .B1(n11798), .B2(pmp_addr_i[480]), .A(n11797), .ZN(n11799)
         );
  NOR2_X1 U11992 ( .A1(n11800), .A2(n11799), .ZN(n11804) );
  NAND2_X1 U11993 ( .A1(n6539), .A2(n11802), .ZN(n11803) );
  OAI211_X1 U11994 ( .C1(n11806), .C2(n11805), .A(n11804), .B(n11803), .ZN(
        n11811) );
  INV_X1 U11995 ( .A(n11807), .ZN(n11808) );
  NOR2_X1 U11996 ( .A1(n11809), .A2(n11808), .ZN(n11810) );
  NOR2_X1 U11997 ( .A1(n11811), .A2(n11810), .ZN(n12106) );
  INV_X1 U11998 ( .A(n11812), .ZN(n12104) );
  INV_X1 U11999 ( .A(n12103), .ZN(n11813) );
  NOR2_X1 U12000 ( .A1(n12104), .A2(n11813), .ZN(n11814) );
  NAND4_X1 U12001 ( .A1(n12108), .A2(n12107), .A3(n12106), .A4(n11814), .ZN(
        n11815) );
  NOR2_X1 U12003 ( .A1(n11819), .A2(n11818), .ZN(n12070) );
  NAND2_X1 U12004 ( .A1(n11820), .A2(data_addr_o_16_), .ZN(n11822) );
  MUX2_X1 U12005 ( .A(n11822), .B(data_addr_o_16_), .S(n11821), .Z(n11875) );
  INV_X1 U12006 ( .A(n11823), .ZN(n11825) );
  NAND2_X1 U12007 ( .A1(n11825), .A2(n11824), .ZN(n11866) );
  INV_X1 U12008 ( .A(n11826), .ZN(n11829) );
  AOI21_X1 U12009 ( .B1(n11829), .B2(n11828), .A(n11827), .ZN(n11865) );
  INV_X1 U12010 ( .A(n11831), .ZN(n11832) );
  OAI21_X1 U12011 ( .B1(n11833), .B2(pmp_addr_i[288]), .A(n11832), .ZN(n11834)
         );
  AOI21_X1 U12012 ( .B1(n6831), .B2(n11835), .A(n11834), .ZN(n11836) );
  OAI211_X1 U12013 ( .C1(n11839), .C2(n11838), .A(n11837), .B(n11836), .ZN(
        n11840) );
  INV_X1 U12014 ( .A(n11840), .ZN(n11856) );
  INV_X1 U12015 ( .A(n11842), .ZN(n11845) );
  INV_X1 U12016 ( .A(n11843), .ZN(n11844) );
  OAI211_X1 U12017 ( .C1(n11846), .C2(n6848), .A(n11845), .B(n11844), .ZN(
        n11855) );
  AOI22_X1 U12018 ( .A1(n6851), .A2(n11850), .B1(n6847), .B2(n11849), .ZN(
        n11854) );
  NAND2_X1 U12019 ( .A1(n6861), .A2(n11852), .ZN(n11853) );
  NAND4_X1 U12020 ( .A1(n11856), .A2(n11855), .A3(n11854), .A4(n11853), .ZN(
        n11860) );
  AND2_X1 U12021 ( .A1(n11858), .A2(n11857), .ZN(n11859) );
  NOR2_X1 U12022 ( .A1(n11860), .A2(n11859), .ZN(n11864) );
  NAND2_X1 U12023 ( .A1(n6860), .A2(n11862), .ZN(n11863) );
  AND4_X1 U12024 ( .A1(n11866), .A2(n11865), .A3(n11864), .A4(n11863), .ZN(
        n11874) );
  NAND2_X1 U12025 ( .A1(n11868), .A2(n11867), .ZN(n11873) );
  INV_X1 U12026 ( .A(n11869), .ZN(n11871) );
  NAND2_X1 U12027 ( .A1(n11871), .A2(n11870), .ZN(n11872) );
  NAND4_X1 U12028 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n11877) );
  NOR2_X1 U12029 ( .A1(n11877), .A2(n11876), .ZN(n12116) );
  INV_X1 U12030 ( .A(n11878), .ZN(n11942) );
  INV_X1 U12031 ( .A(n11879), .ZN(n11881) );
  NAND2_X1 U12032 ( .A1(n11881), .A2(n11880), .ZN(n11886) );
  NAND2_X1 U12033 ( .A1(n11882), .A2(data_addr_o_16_), .ZN(n11884) );
  MUX2_X1 U12034 ( .A(n11884), .B(data_addr_o_16_), .S(n11883), .Z(n11885) );
  AND2_X1 U12035 ( .A1(n11886), .A2(n11885), .ZN(n11940) );
  INV_X1 U12036 ( .A(n11887), .ZN(n11892) );
  INV_X1 U12037 ( .A(n11888), .ZN(n11890) );
  AOI22_X1 U12038 ( .A1(n11892), .A2(n11891), .B1(n11890), .B2(n11889), .ZN(
        n11939) );
  INV_X1 U12039 ( .A(n11893), .ZN(n11895) );
  NAND2_X1 U12040 ( .A1(n11895), .A2(n11894), .ZN(n11926) );
  INV_X1 U12041 ( .A(n11897), .ZN(n11898) );
  OAI22_X1 U12042 ( .A1(n11901), .A2(n11900), .B1(n11899), .B2(n11898), .ZN(
        n11902) );
  AOI21_X1 U12043 ( .B1(n9496), .B2(n11903), .A(n11902), .ZN(n11925) );
  INV_X1 U12044 ( .A(n11904), .ZN(n11914) );
  INV_X1 U12045 ( .A(n11905), .ZN(n11912) );
  OAI21_X1 U12046 ( .B1(n11908), .B2(pmp_addr_i[128]), .A(n11907), .ZN(n11909)
         );
  AOI21_X1 U12047 ( .B1(n9476), .B2(n11910), .A(n11909), .ZN(n11911) );
  OAI211_X1 U12048 ( .C1(n11914), .C2(n11913), .A(n11912), .B(n11911), .ZN(
        n11920) );
  INV_X1 U12049 ( .A(n11915), .ZN(n11918) );
  INV_X1 U12050 ( .A(n11916), .ZN(n11917) );
  NOR2_X1 U12051 ( .A1(n11918), .A2(n11917), .ZN(n11919) );
  NOR2_X1 U12052 ( .A1(n11920), .A2(n11919), .ZN(n11924) );
  NAND2_X1 U12053 ( .A1(n11922), .A2(n11921), .ZN(n11923) );
  NAND4_X1 U12054 ( .A1(n11926), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11936) );
  INV_X1 U12055 ( .A(n11927), .ZN(n11932) );
  INV_X1 U12056 ( .A(n11928), .ZN(n11930) );
  NAND2_X1 U12057 ( .A1(n11930), .A2(n11929), .ZN(n11931) );
  OAI211_X1 U12058 ( .C1(n11934), .C2(n11933), .A(n11932), .B(n11931), .ZN(
        n11935) );
  NOR2_X1 U12059 ( .A1(n11936), .A2(n11935), .ZN(n11938) );
  NAND4_X1 U12060 ( .A1(n11940), .A2(n11939), .A3(n11938), .A4(n11937), .ZN(
        n11941) );
  NOR2_X1 U12061 ( .A1(n11942), .A2(n11941), .ZN(n12117) );
  AOI22_X1 U12062 ( .A1(n12116), .A2(n11944), .B1(n12117), .B2(n11943), .ZN(
        n12069) );
  INV_X1 U12063 ( .A(n11945), .ZN(n12005) );
  INV_X1 U12064 ( .A(n11946), .ZN(n11949) );
  INV_X1 U12065 ( .A(n11947), .ZN(n11948) );
  NAND2_X1 U12066 ( .A1(n11949), .A2(n11948), .ZN(n12003) );
  INV_X1 U12067 ( .A(n11950), .ZN(n11962) );
  INV_X1 U12068 ( .A(n11951), .ZN(n11953) );
  NAND2_X1 U12069 ( .A1(n11953), .A2(n11952), .ZN(n11960) );
  NOR2_X1 U12070 ( .A1(n11955), .A2(n11954), .ZN(n11957) );
  OAI21_X1 U12071 ( .B1(n11958), .B2(n11957), .A(n11956), .ZN(n11959) );
  OAI211_X1 U12072 ( .C1(n11962), .C2(n11961), .A(n11960), .B(n11959), .ZN(
        n11968) );
  INV_X1 U12073 ( .A(n11963), .ZN(n11964) );
  NOR2_X1 U12074 ( .A1(n11966), .A2(n11964), .ZN(n11965) );
  MUX2_X1 U12075 ( .A(n11966), .B(n11965), .S(data_addr_o_16_), .Z(n11967) );
  NOR2_X1 U12076 ( .A1(n11968), .A2(n11967), .ZN(n12002) );
  INV_X1 U12077 ( .A(n11969), .ZN(n11973) );
  AOI22_X1 U12078 ( .A1(n11973), .A2(n9792), .B1(n9806), .B2(n11972), .ZN(
        n12001) );
  INV_X1 U12079 ( .A(n11975), .ZN(n11981) );
  INV_X1 U12080 ( .A(n11976), .ZN(n11978) );
  NAND2_X1 U12081 ( .A1(n11978), .A2(n11977), .ZN(n11980) );
  OAI211_X1 U12082 ( .C1(n11982), .C2(n11981), .A(n11980), .B(n11979), .ZN(
        n11984) );
  AOI211_X1 U12083 ( .C1(n9809), .C2(n11985), .A(n11984), .B(n11983), .ZN(
        n11997) );
  AOI22_X1 U12084 ( .A1(n9826), .A2(n11989), .B1(n9810), .B2(n11988), .ZN(
        n11996) );
  OR2_X1 U12085 ( .A1(n11991), .A2(n11990), .ZN(n11995) );
  OR2_X1 U12086 ( .A1(n11993), .A2(n11992), .ZN(n11994) );
  NAND4_X1 U12087 ( .A1(n11997), .A2(n11996), .A3(n11995), .A4(n11994), .ZN(
        n11999) );
  NOR2_X1 U12088 ( .A1(n11999), .A2(n11998), .ZN(n12000) );
  NAND4_X1 U12089 ( .A1(n12003), .A2(n12002), .A3(n12001), .A4(n12000), .ZN(
        n12004) );
  NOR2_X1 U12090 ( .A1(n12005), .A2(n12004), .ZN(n12115) );
  NAND2_X1 U12091 ( .A1(n12115), .A2(n12006), .ZN(n12068) );
  INV_X1 U12092 ( .A(n12007), .ZN(n12065) );
  INV_X1 U12093 ( .A(n12008), .ZN(n12013) );
  INV_X1 U12094 ( .A(n12009), .ZN(n12010) );
  OAI22_X1 U12095 ( .A1(n12013), .A2(n12012), .B1(n12011), .B2(n12010), .ZN(
        n12020) );
  INV_X1 U12096 ( .A(n12014), .ZN(n12015) );
  OAI22_X1 U12097 ( .A1(n12018), .A2(n12017), .B1(n12016), .B2(n12015), .ZN(
        n12019) );
  NOR2_X1 U12098 ( .A1(n12020), .A2(n12019), .ZN(n12048) );
  OAI22_X1 U12099 ( .A1(n12024), .A2(n12023), .B1(n12022), .B2(n12021), .ZN(
        n12035) );
  INV_X1 U12100 ( .A(n12025), .ZN(n12032) );
  NOR2_X1 U12101 ( .A1(n12027), .A2(pmp_addr_i[352]), .ZN(n12026) );
  MUX2_X1 U12102 ( .A(n12027), .B(n12026), .S(n10130), .Z(n12029) );
  NOR2_X1 U12103 ( .A1(n12029), .A2(n12028), .ZN(n12031) );
  OAI211_X1 U12104 ( .C1(n12033), .C2(n12032), .A(n12031), .B(n12030), .ZN(
        n12034) );
  NOR2_X1 U12105 ( .A1(n12035), .A2(n12034), .ZN(n12047) );
  OAI22_X1 U12106 ( .A1(n12039), .A2(n12038), .B1(n12037), .B2(pmp_addr_i[355]), .ZN(n12040) );
  AOI21_X1 U12107 ( .B1(n10177), .B2(n12041), .A(n12040), .ZN(n12046) );
  OAI21_X1 U12108 ( .B1(n12044), .B2(n12043), .A(n12042), .ZN(n12045) );
  NAND4_X1 U12109 ( .A1(n12048), .A2(n12047), .A3(n12046), .A4(n12045), .ZN(
        n12053) );
  INV_X1 U12110 ( .A(n115), .ZN(n12049) );
  NOR2_X1 U12111 ( .A1(n12051), .A2(n12049), .ZN(n12050) );
  MUX2_X1 U12112 ( .A(n12051), .B(n12050), .S(n9987), .Z(n12052) );
  NOR3_X1 U12113 ( .A1(n12054), .A2(n12053), .A3(n12052), .ZN(n12063) );
  INV_X1 U12114 ( .A(n12055), .ZN(n12056) );
  NAND2_X1 U12115 ( .A1(n12056), .A2(n111), .ZN(n12062) );
  NAND2_X1 U12116 ( .A1(n12057), .A2(n12059), .ZN(n12060) );
  MUX2_X1 U12117 ( .A(n12060), .B(n12059), .S(n12058), .Z(n12061) );
  NAND3_X1 U12118 ( .A1(n12063), .A2(n12062), .A3(n12061), .ZN(n12064) );
  NOR2_X1 U12119 ( .A1(n12065), .A2(n12064), .ZN(n12118) );
  NAND2_X1 U12120 ( .A1(n12118), .A2(n12066), .ZN(n12067) );
  NAND4_X1 U12121 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n12067), .ZN(
        n12125) );
  OAI22_X1 U12122 ( .A1(n12074), .A2(n12073), .B1(n12072), .B2(n12071), .ZN(
        n12078) );
  NOR2_X1 U12123 ( .A1(n12076), .A2(n12075), .ZN(n12077) );
  NOR2_X1 U12124 ( .A1(n12078), .A2(n12077), .ZN(n12098) );
  NOR2_X1 U12125 ( .A1(n12079), .A2(n2590), .ZN(n12088) );
  NAND4_X1 U12126 ( .A1(n12082), .A2(pmp_addr_i[29]), .A3(n12081), .A4(n12080), 
        .ZN(n12084) );
  OAI22_X1 U12127 ( .A1(n12086), .A2(n12085), .B1(n12084), .B2(n12083), .ZN(
        n12087) );
  NOR2_X1 U12128 ( .A1(n12088), .A2(n12087), .ZN(n12097) );
  INV_X1 U12129 ( .A(n12089), .ZN(n12090) );
  NAND2_X1 U12130 ( .A1(n12091), .A2(n12090), .ZN(n12096) );
  INV_X1 U12131 ( .A(n12092), .ZN(n12093) );
  INV_X1 U12134 ( .A(n12099), .ZN(n12100) );
  AOI22_X1 U12135 ( .A1(pmp_addr_i[125]), .A2(n12102), .B1(n12101), .B2(n12100), .ZN(n12110) );
  NOR2_X1 U12136 ( .A1(n12104), .A2(n12103), .ZN(n12105) );
  NAND4_X1 U12137 ( .A1(n12108), .A2(n12107), .A3(n12106), .A4(n12105), .ZN(
        n12109) );
  OAI211_X1 U12138 ( .C1(n12112), .C2(n12111), .A(n12110), .B(n12109), .ZN(
        n12113) );
  NOR2_X1 U12139 ( .A1(n12114), .A2(n12113), .ZN(n12122) );
  AOI22_X1 U12140 ( .A1(pmp_addr_i[317]), .A2(n12116), .B1(n12115), .B2(
        pmp_addr_i[445]), .ZN(n12121) );
  NAND2_X1 U12141 ( .A1(n12117), .A2(pmp_addr_i[157]), .ZN(n12120) );
  NAND2_X1 U12142 ( .A1(n12118), .A2(pmp_addr_i[381]), .ZN(n12119) );
  NAND4_X1 U12143 ( .A1(n12122), .A2(n12121), .A3(n12120), .A4(n12119), .ZN(
        n12124) );
  MUX2_X1 U12144 ( .A(n12125), .B(n12124), .S(n12123), .Z(n12126) );
  NOR2_X1 U12145 ( .A1(n12127), .A2(n12126), .ZN(n12130) );
  INV_X1 U12146 ( .A(n12140), .ZN(n12128) );
  AND2_X1 U12147 ( .A1(n12128), .A2(data_req_i), .ZN(data_req_o) );
  INV_X1 U12148 ( .A(data_gnt_i), .ZN(n12129) );
  NOR2_X1 U12149 ( .A1(n12130), .A2(n12129), .ZN(data_gnt_o) );
  NOR2_X1 U12150 ( .A1(n12132), .A2(n12131), .ZN(n12138) );
  NOR2_X1 U12151 ( .A1(n12134), .A2(n12133), .ZN(n12136) );
  NAND4_X1 U12152 ( .A1(n12138), .A2(n12137), .A3(n12136), .A4(n12135), .ZN(
        n12139) );
  AND2_X1 U12153 ( .A1(n12139), .A2(instr_req_i), .ZN(instr_req_o) );
  NAND3_X1 U12154 ( .A1(data_req_i), .A2(n12140), .A3(data_err_o_BAR), .ZN(
        n12142) );
  NAND2_X1 U12155 ( .A1(data_err_ack_i_BAR), .A2(data_err_state_q), .ZN(n12141) );
  NAND2_X1 U12156 ( .A1(n12142), .A2(n12141), .ZN(n4177) );
  SDFFR_X1 data_err_state_q_reg ( .D(n4177), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(rst_n), .Q(data_err_state_q), .QN(data_err_o_BAR) );
  BUF_X1 U175 ( .A(data_addr_i[28]), .Z(n10747) );
  BUF_X1 U181 ( .A(data_addr_i[29]), .Z(data_addr_o_29_) );
  CLKBUF_X3 U154 ( .A(n2623), .Z(n6005) );
  CLKBUF_X3 U160 ( .A(n5240), .Z(n150) );
  BUF_X2 U928 ( .A(n5163), .Z(n5111) );
  BUF_X2 U998 ( .A(n687), .Z(n4234) );
  INV_X2 U1165 ( .A(n543), .ZN(instr_addr_o_9_) );
  BUF_X2 U430 ( .A(n5996), .Z(n155) );
  CLKBUF_X3 U429 ( .A(n5996), .Z(n154) );
  INV_X2 U66 ( .A(instr_addr_i[9]), .ZN(n3846) );
  INV_X2 U83 ( .A(n2424), .ZN(n12267) );
  INV_X2 U7272 ( .A(data_addr_i[18]), .ZN(n10297) );
  NOR2_X1 U52 ( .A1(n1748), .A2(n1645), .ZN(n5734) );
  INV_X1 U34 ( .A(n3475), .ZN(n1644) );
  CLKBUF_X1 U8 ( .A(n2949), .Z(n3050) );
  NOR2_X1 U207 ( .A1(n11769), .A2(n3923), .ZN(n4681) );
  NOR2_X1 U53 ( .A1(n11587), .A2(n1648), .ZN(n11583) );
  OR2_X2 U107 ( .A1(n3745), .A2(n8079), .ZN(n3758) );
  BUF_X2 U105 ( .A(data_addr_i[7]), .Z(n7816) );
  INV_X1 U106 ( .A(n10473), .ZN(n22) );
  BUF_X2 U103 ( .A(data_addr_i[11]), .Z(data_addr_o_11_) );
  BUF_X2 U98 ( .A(data_addr_i[25]), .Z(n10614) );
  BUF_X2 U7364 ( .A(data_addr_i[30]), .Z(n10919) );
  INV_X1 U10745 ( .A(n11014), .ZN(n10047) );
  BUF_X1 U33 ( .A(n2103), .Z(n999) );
  INV_X2 U992 ( .A(n17), .ZN(n6019) );
  BUF_X2 U1198 ( .A(n3288), .Z(n5192) );
  BUF_X1 U424 ( .A(n191), .Z(n147) );
  INV_X1 U4280 ( .A(n3000), .ZN(n4908) );
  BUF_X1 U419 ( .A(instr_addr_o_18__BAR), .Z(n2082) );
  OAI21_X1 U1912 ( .B1(n5603), .B2(n5530), .A(n5614), .ZN(n1238) );
  AOI211_X1 U4 ( .C1(n1241), .C2(n1240), .A(n1239), .B(n1238), .ZN(n1306) );
  INV_X1 U9 ( .A(n5662), .ZN(n6376) );
  NOR2_X1 U5286 ( .A1(n11807), .A2(n3948), .ZN(n11790) );
  OR2_X1 U484 ( .A1(n3539), .A2(n3574), .ZN(n3626) );
  BUF_X2 U7678 ( .A(data_addr_i[30]), .Z(data_addr_o_30_) );
  BUF_X2 U7081 ( .A(data_addr_i[28]), .Z(n10635) );
  BUF_X1 U7669 ( .A(data_addr_i[23]), .Z(data_addr_o_23_) );
  BUF_X1 U94 ( .A(n9549), .Z(n24) );
  BUF_X1 U7684 ( .A(data_addr_o_20_), .Z(n9935) );
  BUF_X1 U7353 ( .A(data_addr_o_20_), .Z(n10530) );
  INV_X1 U87 ( .A(n4135), .ZN(n4835) );
  BUF_X2 U25 ( .A(n679), .Z(n2733) );
  INV_X1 U5328 ( .A(n4135), .ZN(instr_addr_o_24_) );
  INV_X1 U2984 ( .A(instr_addr_o_4__BAR), .ZN(n5291) );
  INV_X2 U702 ( .A(n4200), .ZN(n5268) );
  INV_X1 U4328 ( .A(n3992), .ZN(n5365) );
  INV_X1 U4324 ( .A(n1026), .ZN(n4909) );
  INV_X1 U3967 ( .A(n2739), .ZN(n6001) );
  INV_X1 U521 ( .A(n2733), .ZN(instr_addr_o_12_) );
  INV_X1 U84 ( .A(n4000), .ZN(n4556) );
  AND3_X2 U57 ( .A1(n1191), .A2(n1189), .A3(n1190), .ZN(n1303) );
  NOR2_X2 U2924 ( .A1(n1921), .A2(n1920), .ZN(n1938) );
  OR2_X2 U2914 ( .A1(n1923), .A2(n5647), .ZN(n1921) );
  OR2_X2 U373 ( .A1(n3100), .A2(n11194), .ZN(n5646) );
  BUF_X1 U300 ( .A(n545), .Z(n2881) );
  BUF_X1 U581 ( .A(n372), .Z(n5163) );
  INV_X1 U3 ( .A(n1569), .ZN(n12170) );
  INV_X1 U10 ( .A(n179), .ZN(n12173) );
  OR2_X1 U11 ( .A1(n3228), .A2(pmp_addr_i[494]), .ZN(n4068) );
  OR2_X1 U12 ( .A1(n3559), .A2(n3558), .ZN(n12176) );
  INV_X1 U13 ( .A(n2881), .ZN(n12202) );
  CLKBUF_X2 U16 ( .A(n537), .Z(n5052) );
  BUF_X1 U18 ( .A(n12132), .Z(n6046) );
  BUF_X1 U26 ( .A(n12134), .Z(n12229) );
  NAND3_X1 U27 ( .A1(n12169), .A2(n7), .A3(n12185), .ZN(n2390) );
  NAND3_X1 U28 ( .A1(n1642), .A2(n338), .A3(n339), .ZN(n12169) );
  NAND3_X1 U29 ( .A1(n12171), .A2(n12170), .A3(n1605), .ZN(n248) );
  NAND2_X1 U30 ( .A1(n1570), .A2(n1594), .ZN(n12171) );
  NAND3_X1 U37 ( .A1(n4667), .A2(n4668), .A3(n162), .ZN(n5020) );
  AND3_X2 U38 ( .A1(n3812), .A2(n12173), .A3(n12172), .ZN(n3827) );
  NAND2_X1 U39 ( .A1(n183), .A2(n185), .ZN(n12172) );
  NOR3_X1 U42 ( .A1(n12176), .A2(n98), .A3(n12175), .ZN(n270) );
  NAND4_X1 U51 ( .A1(n12174), .A2(n12192), .A3(n8081), .A4(n3754), .ZN(n73) );
  NAND3_X1 U54 ( .A1(n3638), .A2(n3636), .A3(n3637), .ZN(n12174) );
  OR2_X2 U60 ( .A1(n3561), .A2(n3560), .ZN(n12175) );
  NAND3_X1 U62 ( .A1(n12177), .A2(n72), .A3(n226), .ZN(n1404) );
  NAND3_X1 U65 ( .A1(n230), .A2(n1401), .A3(n1402), .ZN(n12177) );
  BUF_X2 U75 ( .A(n466), .Z(n5023) );
  BUF_X2 U81 ( .A(n6001), .Z(n12181) );
  CLKBUF_X1 U82 ( .A(instr_addr_i[13]), .Z(n5240) );
  CLKBUF_X1 U85 ( .A(n5253), .Z(n12178) );
  CLKBUF_X3 U100 ( .A(n5253), .Z(n12179) );
  INV_X1 U110 ( .A(n207), .ZN(n5253) );
  BUF_X1 U124 ( .A(n6001), .Z(n12180) );
  BUF_X2 U128 ( .A(n811), .Z(n2424) );
  INV_X1 U147 ( .A(n12217), .ZN(n12203) );
  INV_X1 U155 ( .A(n2881), .ZN(instr_addr_o_10_) );
  INV_X2 U156 ( .A(instr_addr_o_4__BAR), .ZN(n5976) );
  BUF_X1 U164 ( .A(data_addr_i[26]), .Z(n10606) );
  INV_X1 U166 ( .A(n8089), .ZN(n9987) );
  INV_X1 U168 ( .A(n10466), .ZN(n10847) );
  INV_X2 U170 ( .A(n12260), .ZN(n12184) );
  AND2_X1 U178 ( .A1(n6050), .A2(instr_gnt_i), .ZN(instr_gnt_o) );
  AND3_X1 U195 ( .A1(n2213), .A2(n227), .A3(n2212), .ZN(n2292) );
  OAI211_X1 U210 ( .C1(n5208), .C2(n5207), .A(n5216), .B(n5206), .ZN(n5318) );
  OR2_X1 U259 ( .A1(pmp_addr_i[217]), .A2(n5094), .ZN(n12221) );
  BUF_X1 U262 ( .A(n5023), .Z(n2611) );
  INV_X1 U266 ( .A(instr_addr_i[4]), .ZN(n3876) );
  INV_X1 U279 ( .A(n11776), .ZN(n11759) );
  OR2_X1 U280 ( .A1(n6670), .A2(n6669), .ZN(n11776) );
  INV_X1 U282 ( .A(n6069), .ZN(n12220) );
  INV_X1 U285 ( .A(data_addr_o_10_), .ZN(n10701) );
  INV_X1 U291 ( .A(data_addr_i[13]), .ZN(n11006) );
  INV_X1 U308 ( .A(n7820), .ZN(data_addr_o_10_) );
  OAI21_X1 U310 ( .B1(n5587), .B2(n1153), .A(n11907), .ZN(n5567) );
  OR2_X1 U312 ( .A1(n6101), .A2(n6813), .ZN(n12218) );
  INV_X1 U325 ( .A(n7914), .ZN(n12251) );
  AND3_X1 U330 ( .A1(n7873), .A2(n7910), .A3(n12251), .ZN(n7917) );
  AND2_X1 U332 ( .A1(n7573), .A2(n7574), .ZN(n12236) );
  INV_X1 U346 ( .A(pmp_addr_i[423]), .ZN(n3549) );
  AND4_X1 U351 ( .A1(n12236), .A2(n7575), .A3(n7576), .A4(n12188), .ZN(n7602)
         );
  CLKBUF_X1 U352 ( .A(n4505), .Z(n12214) );
  AND2_X1 U358 ( .A1(n499), .A2(pmp_addr_i[367]), .ZN(n3110) );
  AND4_X1 U360 ( .A1(n6089), .A2(n6088), .A3(n6087), .A4(n6086), .ZN(n12230)
         );
  AND2_X1 U410 ( .A1(n3334), .A2(n3337), .ZN(n12240) );
  CLKBUF_X1 U411 ( .A(n3277), .Z(n12227) );
  CLKBUF_X1 U421 ( .A(n207), .Z(n4578) );
  OAI21_X1 U427 ( .B1(n3476), .B2(n3603), .A(n1488), .ZN(n8634) );
  OR2_X1 U428 ( .A1(pmp_addr_i[473]), .A2(n5094), .ZN(n12204) );
  AND2_X1 U518 ( .A1(n3301), .A2(n3287), .ZN(n2463) );
  OR2_X1 U532 ( .A1(n5437), .A2(n5456), .ZN(n12205) );
  INV_X1 U540 ( .A(n11577), .ZN(n11519) );
  INV_X1 U550 ( .A(n1314), .ZN(n12189) );
  CLKBUF_X1 U552 ( .A(n396), .Z(n12215) );
  AND3_X1 U558 ( .A1(n1987), .A2(n2005), .A3(n2014), .ZN(n9) );
  NOR3_X1 U560 ( .A1(n2465), .A2(n2466), .A3(n3268), .ZN(n2474) );
  AND2_X1 U574 ( .A1(n5430), .A2(n5429), .ZN(n12243) );
  INV_X1 U584 ( .A(n12230), .ZN(n11147) );
  AND2_X1 U586 ( .A1(n165), .A2(n5818), .ZN(n2) );
  AND2_X1 U590 ( .A1(n1644), .A2(pmp_cfg_i[98]), .ZN(n12185) );
  AND3_X1 U593 ( .A1(n12206), .A2(n5436), .A3(n12205), .ZN(n12186) );
  AND2_X1 U604 ( .A1(n699), .A2(n8358), .ZN(n12187) );
  AND2_X1 U609 ( .A1(n7580), .A2(n7579), .ZN(n12188) );
  NAND2_X1 U621 ( .A1(n12190), .A2(n12189), .ZN(n1329) );
  NAND2_X1 U640 ( .A1(n1316), .A2(n1315), .ZN(n12190) );
  NAND3_X1 U641 ( .A1(n12235), .A2(n2464), .A3(n2474), .ZN(n2479) );
  NAND4_X1 U644 ( .A1(n3494), .A2(n3493), .A3(n3496), .A4(n3495), .ZN(n12192)
         );
  NAND2_X1 U662 ( .A1(n12193), .A2(n1101), .ZN(n1145) );
  NAND2_X1 U677 ( .A1(n188), .A2(n189), .ZN(n12193) );
  NAND3_X1 U684 ( .A1(n12194), .A2(n496), .A3(n494), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n446), .A2(n493), .ZN(n12194) );
  NAND2_X1 U693 ( .A1(n253), .A2(n677), .ZN(n252) );
  INV_X2 U696 ( .A(n3819), .ZN(n5842) );
  INV_X1 U768 ( .A(instr_addr_i[4]), .ZN(instr_addr_o_4__BAR) );
  CLKBUF_X1 U785 ( .A(n12266), .Z(instr_addr_o_16_) );
  INV_X1 U793 ( .A(n3025), .ZN(n4907) );
  CLKBUF_X1 U795 ( .A(n12264), .Z(n12195) );
  BUF_X2 U798 ( .A(n12264), .Z(instr_addr_o_27_) );
  NOR2_X1 U803 ( .A1(n3798), .A2(n3787), .ZN(n12197) );
  INV_X1 U816 ( .A(n580), .ZN(n12264) );
  AND4_X1 U1005 ( .A1(n2390), .A2(n2388), .A3(n2389), .A4(n2387), .ZN(n12198)
         );
  AND4_X1 U1012 ( .A1(n2390), .A2(n2388), .A3(n2389), .A4(n2387), .ZN(n12137)
         );
  BUF_X1 U1059 ( .A(n5996), .Z(n153) );
  INV_X1 U1111 ( .A(n5115), .ZN(n12199) );
  CLKBUF_X3 U1123 ( .A(n1632), .Z(n5115) );
  INV_X1 U1160 ( .A(n616), .ZN(instr_addr_o_14_) );
  CLKBUF_X3 U1181 ( .A(n433), .Z(n2896) );
  BUF_X2 U1207 ( .A(n433), .Z(n3228) );
  NAND3_X1 U1372 ( .A1(n2596), .A2(n2603), .A3(n12204), .ZN(n2564) );
  NAND2_X1 U1494 ( .A1(instr_addr_o_28_), .A2(n2563), .ZN(n2596) );
  NAND3_X1 U1498 ( .A1(n5226), .A2(n6875), .A3(n11820), .ZN(n12206) );
  NAND2_X1 U1499 ( .A1(n708), .A2(n169), .ZN(n739) );
  AND2_X1 U1515 ( .A1(n2739), .A2(n7362), .ZN(n4245) );
  BUF_X1 U1920 ( .A(n4560), .Z(n12207) );
  BUF_X1 U2130 ( .A(n5313), .Z(n12208) );
  NAND3_X1 U2131 ( .A1(n12209), .A2(n12246), .A3(n2295), .ZN(n12249) );
  NAND3_X1 U2358 ( .A1(n2276), .A2(n2292), .A3(n2277), .ZN(n12209) );
  NAND3_X1 U2435 ( .A1(n12210), .A2(n1786), .A3(n1788), .ZN(n1894) );
  NAND3_X1 U2463 ( .A1(n1771), .A2(n1785), .A3(n84), .ZN(n12210) );
  BUF_X1 U2531 ( .A(n511), .Z(n12211) );
  OAI21_X1 U3409 ( .B1(n1536), .B2(n1535), .A(n12212), .ZN(n1553) );
  OR2_X1 U3410 ( .A1(n1533), .A2(n1534), .ZN(n12212) );
  NAND2_X1 U3418 ( .A1(n223), .A2(n1554), .ZN(n7) );
  BUF_X1 U3496 ( .A(n12157), .Z(n12213) );
  BUF_X1 U3538 ( .A(n2896), .Z(n12217) );
  NAND4_X1 U3571 ( .A1(n12220), .A2(n12219), .A3(n6073), .A4(n12218), .ZN(
        n6077) );
  INV_X1 U3615 ( .A(n6070), .ZN(n12219) );
  NAND3_X1 U3624 ( .A1(n868), .A2(n862), .A3(n12221), .ZN(n832) );
  NAND2_X1 U3658 ( .A1(n6018), .A2(n728), .ZN(n868) );
  NAND4_X1 U3750 ( .A1(n12222), .A2(n87), .A3(n607), .A4(n608), .ZN(n79) );
  NAND3_X1 U3753 ( .A1(n567), .A2(n534), .A3(n535), .ZN(n12222) );
  INV_X1 U4045 ( .A(n12112), .ZN(n12223) );
  NAND2_X1 U4404 ( .A1(n12111), .A2(n12223), .ZN(n12237) );
  CLKBUF_X3 U4453 ( .A(n499), .Z(n5048) );
  NAND2_X1 U4454 ( .A1(n5567), .A2(n9638), .ZN(n12224) );
  NAND2_X1 U4517 ( .A1(n5567), .A2(n9638), .ZN(n12225) );
  INV_X1 U4584 ( .A(n3992), .ZN(n12226) );
  INV_X1 U4585 ( .A(n2881), .ZN(n213) );
  AND2_X1 U4890 ( .A1(n12184), .A2(n8652), .ZN(n8564) );
  INV_X1 U5401 ( .A(n679), .ZN(n5245) );
  AND2_X1 U5923 ( .A1(n135), .A2(n8653), .ZN(n1482) );
  CLKBUF_X1 U6040 ( .A(n3992), .Z(n135) );
  INV_X1 U6236 ( .A(instr_addr_i[17]), .ZN(n12228) );
  INV_X2 U6409 ( .A(n5023), .ZN(n5277) );
  AND2_X1 U6601 ( .A1(n135), .A2(n7855), .ZN(n2485) );
  INV_X1 U6610 ( .A(instr_addr_i[31]), .ZN(n511) );
  BUF_X1 U6615 ( .A(n3295), .Z(n4005) );
  INV_X1 U6616 ( .A(n3295), .ZN(n5136) );
  INV_X1 U6617 ( .A(n511), .ZN(n5154) );
  INV_X2 U6953 ( .A(n8089), .ZN(n11014) );
  NOR2_X1 U6954 ( .A1(n1258), .A2(n1165), .ZN(n177) );
  AOI22_X1 U6985 ( .A1(n4603), .A2(n4616), .B1(n4602), .B2(pmp_addr_i[424]), 
        .ZN(n4618) );
  NAND4_X1 U7072 ( .A1(n12232), .A2(n12231), .A3(n5939), .A4(n5938), .ZN(n58)
         );
  NAND2_X1 U7077 ( .A1(n5936), .A2(n5935), .ZN(n12231) );
  NAND2_X1 U7094 ( .A1(n5934), .A2(n5942), .ZN(n12232) );
  NAND4_X1 U7099 ( .A1(n12234), .A2(n12233), .A3(n5888), .A4(n5887), .ZN(n5909) );
  INV_X1 U7100 ( .A(n5885), .ZN(n12233) );
  INV_X1 U7112 ( .A(n5884), .ZN(n12234) );
  OR2_X1 U7128 ( .A1(n3846), .A2(pmp_addr_i[167]), .ZN(n5038) );
  NAND3_X1 U7283 ( .A1(n12247), .A2(n2431), .A3(n12248), .ZN(n12235) );
  NAND4_X1 U7406 ( .A1(n12239), .A2(n12238), .A3(n11815), .A4(n12237), .ZN(
        n11818) );
  NAND2_X1 U7645 ( .A1(n12101), .A2(n12099), .ZN(n12238) );
  NAND2_X1 U7676 ( .A1(n12102), .A2(n11758), .ZN(n12239) );
  NAND4_X1 U7703 ( .A1(n3339), .A2(n3335), .A3(n3338), .A4(n12240), .ZN(n3348)
         );
  NAND3_X1 U7745 ( .A1(n8949), .A2(n8948), .A3(n156), .ZN(n15) );
  NAND2_X1 U7822 ( .A1(n3170), .A2(n3154), .ZN(n3172) );
  NAND2_X1 U7854 ( .A1(n4836), .A2(n3153), .ZN(n3170) );
  NAND3_X1 U7901 ( .A1(n3869), .A2(n12250), .A3(n3868), .ZN(n12134) );
  NAND3_X1 U8574 ( .A1(n12242), .A2(n877), .A3(n272), .ZN(n1406) );
  AOI21_X1 U8577 ( .B1(n12241), .B2(n842), .A(n840), .ZN(n876) );
  OAI211_X1 U8578 ( .C1(n830), .C2(n831), .A(n829), .B(n828), .ZN(n12241) );
  NAND2_X1 U8850 ( .A1(n783), .A2(n782), .ZN(n12242) );
  NAND3_X1 U8855 ( .A1(n63), .A2(n1938), .A3(n1936), .ZN(n1966) );
  NAND4_X1 U9094 ( .A1(n12245), .A2(n12244), .A3(n5432), .A4(n12243), .ZN(
        n5468) );
  NAND2_X1 U9298 ( .A1(n5419), .A2(n11849), .ZN(n12244) );
  NAND2_X1 U9416 ( .A1(n5418), .A2(n11824), .ZN(n12245) );
  NAND2_X1 U10151 ( .A1(n2292), .A2(n2291), .ZN(n12246) );
  INV_X2 U11294 ( .A(n376), .ZN(n4753) );
  INV_X1 U11350 ( .A(n2404), .ZN(n12247) );
  NAND2_X1 U11667 ( .A1(n2405), .A2(n2428), .ZN(n12248) );
  NAND3_X1 U11857 ( .A1(n5082), .A2(n5081), .A3(n5080), .ZN(n265) );
  NAND4_X1 U11886 ( .A1(n12249), .A2(n12253), .A3(n6935), .A4(pmp_cfg_i[74]), 
        .ZN(n2387) );
  NAND3_X1 U11887 ( .A1(n3205), .A2(n249), .A3(n254), .ZN(n12250) );
  NAND4_X1 U11888 ( .A1(n9340), .A2(n11027), .A3(n11028), .A4(n12252), .ZN(
        n12127) );
  AND2_X1 U11973 ( .A1(n9339), .A2(n9341), .ZN(n12252) );
  INV_X1 U11974 ( .A(n2338), .ZN(n244) );
  OAI21_X1 U12002 ( .B1(n2300), .B2(n2336), .A(n2299), .ZN(n2338) );
  NAND3_X1 U12132 ( .A1(n245), .A2(n2384), .A3(n2383), .ZN(n12253) );
  BUF_X2 U12133 ( .A(n687), .Z(n499) );
  NAND4_X1 U12157 ( .A1(n12254), .A2(n12097), .A3(n12096), .A4(n12098), .ZN(
        n12114) );
  NAND2_X1 U12158 ( .A1(n12094), .A2(n12093), .ZN(n12254) );
  NAND4_X1 U12159 ( .A1(n12255), .A2(n11580), .A3(n11579), .A4(n11581), .ZN(
        n11819) );
  NAND2_X1 U12160 ( .A1(n12094), .A2(n12092), .ZN(n12255) );
  NAND2_X1 U12161 ( .A1(n10646), .A2(n10647), .ZN(n11577) );
  NAND2_X1 U12162 ( .A1(n12256), .A2(n12257), .ZN(n95) );
  NAND4_X1 U12163 ( .A1(n4797), .A2(n4800), .A3(n4799), .A4(n4798), .ZN(n12256) );
  NAND2_X1 U12164 ( .A1(n4758), .A2(n4800), .ZN(n12257) );
  CLKBUF_X1 U12165 ( .A(n2739), .Z(n616) );
  INV_X1 U12166 ( .A(n1632), .ZN(n4560) );
endmodule



    module riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16 ( 
        clk, rst_n, core_id_i, cluster_id_i, mtvec_o, utvec_o, boot_addr_i, 
        csr_addr_i, csr_wdata_i, csr_op_i, csr_rdata_o, frm_o, fprec_o, 
        fflags_i, fflags_we_i, m_irq_enable_o, u_irq_enable_o, csr_irq_sec_i, 
        sec_lvl_o, mepc_o, uepc_o, debug_mode_i, debug_cause_i, 
        debug_csr_save_i, depc_o, debug_single_step_o, debug_ebreakm_o, 
        debug_ebreaku_o, pmp_addr_o, pmp_cfg_o, priv_lvl_o, pc_if_i, pc_id_i, 
        pc_ex_i, csr_save_if_i, csr_save_id_i, csr_restore_mret_i, 
        csr_restore_uret_i, csr_restore_dret_i, csr_save_cause_i, hwlp_start_i, 
        hwlp_end_i, hwlp_cnt_i, hwlp_data_o, hwlp_regid_o, hwlp_we_o, 
        id_valid_i, is_compressed_i, imiss_i, pc_set_i, jump_i, branch_i, 
        branch_taken_i, ld_stall_i, jr_stall_i, pipeline_stall_i, 
        apu_typeconflict_i, apu_contention_i, apu_dep_i, apu_wb_i, mem_load_i, 
        mem_store_i, ext_counters_i, csr_cause_i_5__BAR, csr_cause_i_4_, 
        csr_cause_i_3_, csr_cause_i_2_, csr_cause_i_0_, csr_save_ex_i_BAR, 
        csr_cause_i_1__BAR, is_decoding_i, csr_access_i_BAR );
  input [3:0] core_id_i;
  input [5:0] cluster_id_i;
  output [23:0] mtvec_o;
  output [23:0] utvec_o;
  input [30:0] boot_addr_i;
  input [11:0] csr_addr_i;
  input [31:0] csr_wdata_i;
  input [1:0] csr_op_i;
  output [31:0] csr_rdata_o;
  output [2:0] frm_o;
  output [4:0] fprec_o;
  input [4:0] fflags_i;
  output [31:0] mepc_o;
  output [31:0] uepc_o;
  input [2:0] debug_cause_i;
  output [31:0] depc_o;
  output [511:0] pmp_addr_o;
  output [127:0] pmp_cfg_o;
  output [1:0] priv_lvl_o;
  input [31:0] pc_if_i;
  input [31:0] pc_id_i;
  input [31:0] pc_ex_i;
  input [63:0] hwlp_start_i;
  input [63:0] hwlp_end_i;
  input [63:0] hwlp_cnt_i;
  output [31:0] hwlp_data_o;
  output [0:0] hwlp_regid_o;
  output [2:0] hwlp_we_o;
  input [1:2] ext_counters_i;
  input clk, rst_n, fflags_we_i, csr_irq_sec_i, debug_mode_i, debug_csr_save_i,
         csr_save_if_i, csr_save_id_i, csr_restore_mret_i, csr_restore_uret_i,
         csr_restore_dret_i, csr_save_cause_i, id_valid_i, is_compressed_i,
         imiss_i, pc_set_i, jump_i, branch_i, branch_taken_i, ld_stall_i,
         jr_stall_i, pipeline_stall_i, apu_typeconflict_i, apu_contention_i,
         apu_dep_i, apu_wb_i, mem_load_i, mem_store_i, csr_cause_i_5__BAR,
         csr_cause_i_4_, csr_cause_i_3_, csr_cause_i_2_, csr_cause_i_0_,
         csr_save_ex_i_BAR, csr_cause_i_1__BAR, is_decoding_i,
         csr_access_i_BAR;
  output m_irq_enable_o, u_irq_enable_o, sec_lvl_o, debug_single_step_o,
         debug_ebreakm_o, debug_ebreaku_o;
  wire   csr_access_i, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         \priv_lvl_o[0] , is_decoding_i_BAR, dcsr_q_xdebugver__30_,
         dcsr_q_zero2__27_, dcsr_q_zero2__26_, dcsr_q_zero2__25_,
         dcsr_q_zero2__24_, dcsr_q_zero2__23_, dcsr_q_zero2__22_,
         dcsr_q_zero2__21_, dcsr_q_zero2__20_, dcsr_q_zero2__19_,
         dcsr_q_zero2__18_, dcsr_q_zero2__17_, dcsr_q_zero2__16_,
         dcsr_q_zero1_, dcsr_q_ebreaks_, dcsr_q_stepie_, dcsr_q_cause__8_,
         dcsr_q_cause__7_, dcsr_q_cause__6_, dcsr_q_zero0_, dcsr_q_prv__1_,
         dcsr_q_prv__0_, N2756, id_valid_q, PCCR_inc_0_, PCCR_inc_q_0_, n2022,
         n2024, n2025, n2026, n2033, n2034, n2035, n2041, n2051, n2056, n2057,
         n2058, n2062, n2065, n2068, n2071, n2082, n2088, n2089, n2090, n2094,
         n2097, n2098, n2099, n2103, n2105, n2114, n2120, n2121, n2122, n2126,
         n2129, n2135, n2136, n2138, n2663, n2733, n2737, n2741, n2761, n2764,
         n2807, n4183, n1675, n55, n56, n57, n58, n60, n62, n63, n64, n65, n67,
         n68, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n168, n169, n170, n171, n174, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n195, n196, n197, n198, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n241, n243, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n387, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n594, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n821, n822, n823, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n886, n890,
         n893, n894, n897, n898, n901, n902, n905, n906, n909, n910, n911,
         n914, n919, n922, n923, n926, n928, n929, n931, n932, n4184, n935,
         n936, n937, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n964, n966, n967, n968, n969, n970, n971, n975, n979, n983,
         n984, n985, n986, n987, n989, n990, n995, n996, n998, n1000, n1002,
         n1004, n1006, n1007, n1009, n1011, n1012, n1018, n1020, n1022, n1024,
         n1028, n1029, n1031, n1037, n1038, n1039, n1041, n1042, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1054, n1056, n1057, n1059, n1061,
         n1065, n1067, n1069, n1070, n1072, n1074, n1076, n1078, n1079, n1081,
         n1085, n1087, n1088, n1089, n1090, n1091, n1092, n1094, n1096, n1098,
         n1100, n1102, n1106, n1107, n1109, n1113, n1115, n1118, n1119, n1122,
         n1123, n1124, n1125, n1126, n1127, n1129, n1130, n1132, n1134, n1136,
         n1140, n1141, n1142, n1144, n1148, n1154, n1155, n1157, n1159, n1161,
         n1163, n1164, n1165, n1166, n1167, n1168, n1170, n1172, n1174, n1178,
         n1181, n1182, n1183, n1185, n1198, n1199, n1209, n1212, n1221, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1379, n1380, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1414, n1415, n1416, n1418,
         n1419, n1421, n1422, n1423, n1424, n1426, n1427, n1428, n1429, n1434,
         n1437, n1438, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1449, n1450, n1452, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1505, n1520, n1544, n1553, n1579, n1580, n1584,
         n1607, n1622, n1677, n1678, n1681, n1682, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1702, n1704, n1705, n1706, n1714, n1715, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3913,
         n3914, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3944, n3946, n3948, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3960, n3961, n3962,
         n3964, n3966, n3967, n3969, n3970, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4099, n4100,
         n4101, n4103, n4105, n4106, n4107, n4109, n4110, n4112, n4113, n4114,
         n4115, n4116, n4117, n4119, n4120, n4121, n4122, n4123, n4125, n4127,
         n4128, n4130, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4147, n4148, n4149, n4151,
         n4153, n4155, n4157, n4159, n4161, n4163, n4165, n4167, n4169, n4171,
         n4173, n4175, n4176, n4178, n4180;
  wire   [6:0] mstatus_q;
  wire   [31:0] mscratch_q;
  wire   [5:0] mcause_q;
  wire   [31:0] dscratch0_q;
  wire   [31:0] dscratch1_q;
  wire   [5:0] ucause_q;
  wire   [31:0] mepc_n;
  wire   [31:0] uepc_n;
  wire   [31:0] depc_n;
  wire   [4:0] mstatus_n;
  wire   [11:0] PCER_q;
  wire   [1:0] PCMR_q;
  wire   [31:0] PCCR_q;
  wire   [30:0] PCCR_n;
  wire   [1:0] PCMR_n;
  wire   [11:0] PCER_n;
  assign csr_access_i = csr_access_i_BAR;
  assign sec_lvl_o = \priv_lvl_o[0] ;
  assign priv_lvl_o[0] = \priv_lvl_o[0] ;
  assign is_decoding_i_BAR = is_decoding_i;
  assign hwlp_data_o[13] = n501;
  assign hwlp_data_o[7] = n520;
  assign hwlp_data_o[2] = n564;
  assign hwlp_data_o[29] = n929;

  CLKBUF_X1 U11 ( .A(n990), .Z(n64) );
  CLKBUF_X2 U14 ( .A(n582), .Z(n65) );
  INV_X1 U16 ( .A(n1403), .ZN(n1440) );
  INV_X1 U18 ( .A(n241), .ZN(n864) );
  NOR4_X1 U20 ( .A1(csr_addr_i[4]), .A2(n106), .A3(n108), .A4(n133), .ZN(n121)
         );
  INV_X1 U21 ( .A(csr_op_i[1]), .ZN(n708) );
  NOR2_X1 U22 ( .A1(n811), .A2(n134), .ZN(n923) );
  NAND2_X1 U23 ( .A1(n3700), .A2(n1385), .ZN(n1198) );
  AOI21_X1 U24 ( .B1(csr_wdata_i[22]), .B2(n1257), .A(n292), .ZN(n1007) );
  AOI21_X1 U25 ( .B1(csr_wdata_i[5]), .B2(n1257), .A(n326), .ZN(n970) );
  AND2_X1 U26 ( .A1(csr_op_i[1]), .A2(csr_op_i[0]), .ZN(n1257) );
  OR2_X1 U30 ( .A1(n174), .A2(n1198), .ZN(n1446) );
  AND2_X1 U31 ( .A1(n958), .A2(n956), .ZN(n67) );
  NAND3_X1 U39 ( .A1(n1386), .A2(n1385), .A3(n1384), .ZN(n1438) );
  INV_X2 U40 ( .A(n551), .ZN(n767) );
  NAND3_X1 U42 ( .A1(n954), .A2(n955), .A3(n958), .ZN(n967) );
  NAND2_X2 U43 ( .A1(n790), .A2(n1385), .ZN(n1368) );
  INV_X1 U45 ( .A(csr_wdata_i[25]), .ZN(n193) );
  INV_X1 U46 ( .A(n1675), .ZN(n68) );
  INV_X4 U48 ( .A(n1257), .ZN(n1362) );
  AOI211_X2 U49 ( .C1(csr_addr_i[11]), .C2(n196), .A(n673), .B(n141), .ZN(n761) );
  OAI21_X1 U50 ( .B1(n384), .B2(csr_wdata_i[18]), .A(n383), .ZN(n1675) );
  AND4_X1 U51 ( .A1(n1396), .A2(n1376), .A3(n1375), .A4(n1374), .ZN(n70) );
  OR2_X1 U52 ( .A1(n118), .A2(n117), .ZN(n71) );
  NOR2_X1 U53 ( .A1(n133), .A2(n122), .ZN(n146) );
  NOR2_X1 U54 ( .A1(n98), .A2(n79), .ZN(n813) );
  NOR2_X1 U55 ( .A1(n353), .A2(n881), .ZN(n743) );
  OR2_X1 U56 ( .A1(\priv_lvl_o[0] ), .A2(priv_lvl_o[1]), .ZN(n846) );
  NOR2_X1 U57 ( .A1(n743), .A2(n742), .ZN(n826) );
  INV_X1 U58 ( .A(n708), .ZN(n814) );
  INV_X1 U59 ( .A(csr_wdata_i[6]), .ZN(n1256) );
  NOR2_X1 U60 ( .A1(n814), .A2(csr_op_i[0]), .ZN(n1394) );
  NOR2_X1 U61 ( .A1(n901), .A2(n353), .ZN(n1429) );
  NAND2_X1 U62 ( .A1(csr_wdata_i[27]), .A2(n1362), .ZN(n276) );
  NAND2_X1 U63 ( .A1(csr_wdata_i[20]), .A2(n1362), .ZN(n311) );
  NOR2_X1 U64 ( .A1(n171), .A2(n1198), .ZN(n241) );
  NOR2_X1 U65 ( .A1(n115), .A2(n114), .ZN(n1371) );
  INV_X1 U66 ( .A(n679), .ZN(n886) );
  OAI21_X1 U67 ( .B1(n131), .B2(csr_wdata_i[31]), .A(n130), .ZN(n935) );
  OAI21_X1 U68 ( .B1(n659), .B2(csr_wdata_i[30]), .A(n658), .ZN(n931) );
  OAI21_X1 U69 ( .B1(n636), .B2(csr_wdata_i[29]), .A(n635), .ZN(n929) );
  INV_X1 U70 ( .A(hwlp_data_o[28]), .ZN(n1422) );
  INV_X1 U71 ( .A(hwlp_data_o[27]), .ZN(n1421) );
  INV_X1 U72 ( .A(hwlp_data_o[24]), .ZN(n1416) );
  INV_X1 U73 ( .A(hwlp_data_o[20]), .ZN(n1412) );
  INV_X1 U74 ( .A(hwlp_data_o[19]), .ZN(n1411) );
  INV_X1 U81 ( .A(n1438), .ZN(n1437) );
  NAND2_X1 U82 ( .A1(priv_lvl_o[1]), .A2(\priv_lvl_o[0] ), .ZN(n940) );
  NOR2_X1 U83 ( .A1(debug_csr_save_i), .A2(n940), .ZN(n1042) );
  INV_X1 U84 ( .A(n846), .ZN(n1047) );
  NOR2_X1 U85 ( .A1(n1042), .A2(n1047), .ZN(n1039) );
  INV_X1 U86 ( .A(csr_restore_dret_i), .ZN(n72) );
  NOR3_X1 U87 ( .A1(csr_restore_mret_i), .A2(csr_save_cause_i), .A3(
        csr_restore_uret_i), .ZN(n830) );
  AOI22_X1 U88 ( .A1(n1039), .A2(csr_save_cause_i), .B1(n72), .B2(n830), .ZN(
        n76) );
  NOR2_X1 U89 ( .A1(mstatus_q[2]), .A2(mstatus_q[1]), .ZN(n834) );
  AOI21_X1 U90 ( .B1(mstatus_q[1]), .B2(mstatus_q[2]), .A(n834), .ZN(n943) );
  NAND2_X1 U91 ( .A1(csr_restore_mret_i), .A2(n943), .ZN(n73) );
  NAND2_X1 U92 ( .A1(n76), .A2(n73), .ZN(n823) );
  NOR2_X1 U93 ( .A1(csr_irq_sec_i), .A2(csr_cause_i_5__BAR), .ZN(n850) );
  NOR2_X1 U94 ( .A1(n850), .A2(n846), .ZN(n74) );
  INV_X1 U95 ( .A(csr_save_cause_i), .ZN(n1038) );
  AOI21_X1 U97 ( .B1(csr_save_cause_i), .B2(n74), .A(n942), .ZN(n1122) );
  INV_X1 U98 ( .A(csr_restore_mret_i), .ZN(n847) );
  NOR2_X1 U99 ( .A1(n834), .A2(n847), .ZN(n829) );
  INV_X1 U100 ( .A(n829), .ZN(n75) );
  NAND3_X1 U101 ( .A1(n76), .A2(n1122), .A3(n75), .ZN(n821) );
  AOI21_X1 U102 ( .B1(csr_restore_dret_i), .B2(dcsr_q_prv__0_), .A(n821), .ZN(
        n77) );
  AOI21_X1 U103 ( .B1(n1481), .B2(n823), .A(n77), .ZN(n78) );
  INV_X1 U104 ( .A(n78), .ZN(n1449) );
  NAND2_X1 U105 ( .A1(csr_wdata_i[0]), .A2(n1362), .ZN(n758) );
  INV_X1 U106 ( .A(csr_addr_i[5]), .ZN(n157) );
  INV_X1 U107 ( .A(csr_addr_i[6]), .ZN(n100) );
  AND2_X1 U108 ( .A1(csr_addr_i[7]), .A2(n100), .ZN(n80) );
  INV_X1 U109 ( .A(csr_addr_i[10]), .ZN(n98) );
  NAND2_X1 U110 ( .A1(csr_addr_i[9]), .A2(csr_addr_i[8]), .ZN(n79) );
  INV_X1 U111 ( .A(n813), .ZN(n196) );
  NOR2_X1 U112 ( .A1(n196), .A2(csr_addr_i[11]), .ZN(n154) );
  NAND4_X1 U113 ( .A1(n157), .A2(n80), .A3(n154), .A4(n1715), .ZN(n1240) );
  INV_X2 U114 ( .A(n1240), .ZN(n790) );
  INV_X2 U115 ( .A(n1394), .ZN(n1385) );
  NAND4_X1 U116 ( .A1(PCMR_q[1]), .A2(PCCR_q[1]), .A3(PCCR_q[8]), .A4(
        PCCR_q[15]), .ZN(n85) );
  NAND4_X1 U117 ( .A1(PCCR_q[11]), .A2(PCCR_q[12]), .A3(PCCR_q[13]), .A4(
        PCCR_q[14]), .ZN(n84) );
  NAND4_X1 U118 ( .A1(PCCR_q[7]), .A2(PCCR_q[4]), .A3(PCCR_q[6]), .A4(
        PCCR_q[5]), .ZN(n81) );
  NOR3_X1 U119 ( .A1(n1460), .A2(n1452), .A3(n81), .ZN(n82) );
  NAND4_X1 U120 ( .A1(PCCR_q[0]), .A2(PCCR_q[25]), .A3(PCCR_q[26]), .A4(n82), 
        .ZN(n83) );
  NOR3_X1 U121 ( .A1(n85), .A2(n84), .A3(n83), .ZN(n92) );
  NAND4_X1 U122 ( .A1(PCCR_q[31]), .A2(PCCR_q[17]), .A3(PCCR_q[18]), .A4(
        PCCR_q[24]), .ZN(n89) );
  NAND4_X1 U123 ( .A1(PCCR_q[27]), .A2(PCCR_q[28]), .A3(PCCR_q[29]), .A4(
        PCCR_q[30]), .ZN(n88) );
  NAND4_X1 U124 ( .A1(PCCR_q[9]), .A2(PCCR_q[10]), .A3(PCCR_q[16]), .A4(
        PCCR_q[23]), .ZN(n87) );
  NAND4_X1 U125 ( .A1(PCCR_q[22]), .A2(PCCR_q[19]), .A3(PCCR_q[20]), .A4(
        PCCR_q[21]), .ZN(n86) );
  NOR4_X1 U126 ( .A1(n89), .A2(n88), .A3(n87), .A4(n86), .ZN(n91) );
  NAND2_X1 U127 ( .A1(n1368), .A2(PCCR_inc_q_0_), .ZN(n90) );
  AOI21_X1 U128 ( .B1(n92), .B2(n91), .A(n90), .ZN(n1271) );
  AND3_X1 U129 ( .A1(n1257), .A2(csr_wdata_i[0]), .A3(n790), .ZN(n93) );
  NOR2_X1 U130 ( .A1(n1366), .A2(n93), .ZN(n95) );
  AOI21_X1 U131 ( .B1(n790), .B2(csr_op_i[0]), .A(n1271), .ZN(n1315) );
  CLKBUF_X1 U132 ( .A(n1315), .Z(n1298) );
  INV_X1 U133 ( .A(n1298), .ZN(n94) );
  MUX2_X1 U134 ( .A(n95), .B(n94), .S(PCCR_q[0]), .Z(n96) );
  OAI21_X1 U135 ( .B1(n758), .B2(n1368), .A(n96), .ZN(n97) );
  INV_X1 U136 ( .A(n97), .ZN(n1450) );
  NOR3_X1 U138 ( .A1(csr_addr_i[6]), .A2(csr_addr_i[7]), .A3(csr_addr_i[5]), 
        .ZN(n138) );
  INV_X1 U139 ( .A(csr_addr_i[4]), .ZN(n107) );
  NAND2_X1 U140 ( .A1(n138), .A2(n107), .ZN(n122) );
  OR3_X1 U141 ( .A1(csr_addr_i[10]), .A2(csr_addr_i[9]), .A3(csr_addr_i[8]), 
        .ZN(n139) );
  OR2_X1 U142 ( .A1(n122), .A2(n139), .ZN(n741) );
  INV_X1 U143 ( .A(csr_addr_i[1]), .ZN(n114) );
  NAND2_X1 U144 ( .A1(n114), .A2(csr_addr_i[0]), .ZN(n1224) );
  INV_X1 U145 ( .A(n1224), .ZN(n101) );
  INV_X1 U146 ( .A(csr_addr_i[2]), .ZN(n1372) );
  NOR2_X1 U147 ( .A1(n1372), .A2(csr_addr_i[3]), .ZN(n909) );
  NAND2_X1 U148 ( .A1(n101), .A2(n909), .ZN(n901) );
  NOR2_X1 U149 ( .A1(n741), .A2(n901), .ZN(n1398) );
  NAND2_X1 U150 ( .A1(n3700), .A2(n1398), .ZN(n647) );
  NOR2_X1 U151 ( .A1(csr_addr_i[2]), .A2(n1224), .ZN(n1046) );
  INV_X1 U152 ( .A(csr_addr_i[3]), .ZN(n811) );
  NAND2_X1 U153 ( .A1(n1046), .A2(n811), .ZN(n679) );
  NAND3_X1 U154 ( .A1(csr_addr_i[9]), .A2(csr_addr_i[8]), .A3(n98), .ZN(n133)
         );
  NOR2_X1 U155 ( .A1(csr_addr_i[7]), .A2(csr_addr_i[5]), .ZN(n99) );
  NAND3_X1 U156 ( .A1(csr_addr_i[6]), .A2(n99), .A3(n107), .ZN(n104) );
  NOR2_X1 U157 ( .A1(n133), .A2(n104), .ZN(n105) );
  NAND2_X1 U158 ( .A1(n886), .A2(n105), .ZN(n1130) );
  NOR2_X1 U159 ( .A1(csr_addr_i[11]), .A2(n1130), .ZN(n582) );
  AOI22_X1 U160 ( .A1(n790), .A2(PCCR_q[31]), .B1(n65), .B2(mepc_o[31]), .ZN(
        n103) );
  NAND3_X1 U161 ( .A1(csr_addr_i[7]), .A2(csr_addr_i[5]), .A3(n100), .ZN(n106)
         );
  NOR2_X1 U162 ( .A1(csr_addr_i[3]), .A2(csr_addr_i[2]), .ZN(n116) );
  INV_X1 U163 ( .A(n116), .ZN(n108) );
  NAND2_X1 U164 ( .A1(n121), .A2(n101), .ZN(n171) );
  NOR2_X1 U165 ( .A1(csr_addr_i[11]), .A2(n171), .ZN(n180) );
  CLKBUF_X1 U166 ( .A(n180), .Z(n800) );
  INV_X1 U167 ( .A(csr_addr_i[0]), .ZN(n115) );
  NAND2_X1 U168 ( .A1(n115), .A2(n114), .ZN(n1223) );
  INV_X1 U169 ( .A(n1223), .ZN(n119) );
  NAND2_X1 U170 ( .A1(n121), .A2(n119), .ZN(n387) );
  OR2_X1 U171 ( .A1(csr_addr_i[11]), .A2(n387), .ZN(n551) );
  AOI22_X1 U172 ( .A1(n800), .A2(n30), .B1(n767), .B2(n42), .ZN(n102) );
  OAI211_X1 U173 ( .C1(n647), .C2(n1469), .A(n103), .B(n102), .ZN(n129) );
  NAND3_X1 U174 ( .A1(csr_addr_i[6]), .A2(csr_addr_i[7]), .A3(n107), .ZN(n156)
         );
  NOR2_X1 U175 ( .A1(csr_addr_i[5]), .A2(n156), .ZN(n812) );
  NAND2_X1 U176 ( .A1(n154), .A2(n812), .ZN(n120) );
  NAND2_X1 U177 ( .A1(n115), .A2(csr_addr_i[1]), .ZN(n1226) );
  INV_X1 U178 ( .A(n1226), .ZN(n1370) );
  NAND2_X1 U179 ( .A1(n1370), .A2(n909), .ZN(n905) );
  NOR2_X1 U180 ( .A1(n120), .A2(n905), .ZN(n641) );
  CLKBUF_X1 U181 ( .A(n641), .Z(n690) );
  NOR2_X1 U182 ( .A1(n139), .A2(n104), .ZN(n109) );
  NAND2_X1 U183 ( .A1(n886), .A2(n109), .ZN(n950) );
  NOR2_X1 U184 ( .A1(csr_addr_i[11]), .A2(n950), .ZN(n548) );
  CLKBUF_X1 U185 ( .A(n548), .Z(n801) );
  AOI22_X1 U186 ( .A1(n690), .A2(hwlp_cnt_i[63]), .B1(n801), .B2(uepc_o[31]), 
        .ZN(n113) );
  NOR2_X1 U187 ( .A1(csr_addr_i[2]), .A2(n1223), .ZN(n914) );
  NAND2_X1 U188 ( .A1(n914), .A2(n811), .ZN(n881) );
  INV_X1 U189 ( .A(n105), .ZN(n118) );
  NOR2_X1 U192 ( .A1(csr_addr_i[11]), .A2(n1374), .ZN(n153) );
  NOR2_X1 U194 ( .A1(n120), .A2(n881), .ZN(n136) );
  CLKBUF_X1 U195 ( .A(n136), .Z(n696) );
  AOI22_X1 U196 ( .A1(n691), .A2(mscratch_q[31]), .B1(n696), .B2(
        hwlp_start_i[31]), .ZN(n112) );
  NOR2_X1 U197 ( .A1(n107), .A2(n106), .ZN(n132) );
  NAND2_X1 U198 ( .A1(n154), .A2(n132), .ZN(n152) );
  NOR2_X1 U199 ( .A1(n108), .A2(n1226), .ZN(n890) );
  INV_X1 U200 ( .A(n890), .ZN(n117) );
  NOR2_X1 U201 ( .A1(n152), .A2(n117), .ZN(n410) );
  CLKBUF_X1 U202 ( .A(n410), .Z(n695) );
  NOR2_X1 U203 ( .A1(n679), .A2(n152), .ZN(n715) );
  CLKBUF_X1 U204 ( .A(n715), .Z(n701) );
  AOI22_X1 U205 ( .A1(n695), .A2(dscratch0_q[31]), .B1(n701), .B2(depc_o[31]), 
        .ZN(n111) );
  NOR2_X1 U206 ( .A1(n120), .A2(n679), .ZN(n716) );
  NAND2_X1 U207 ( .A1(n890), .A2(n109), .ZN(n1199) );
  NOR2_X1 U208 ( .A1(csr_addr_i[11]), .A2(n1199), .ZN(n789) );
  AOI22_X1 U209 ( .A1(n716), .A2(hwlp_end_i[31]), .B1(n789), .B2(ucause_q[5]), 
        .ZN(n110) );
  NAND4_X1 U210 ( .A1(n113), .A2(n112), .A3(n111), .A4(n110), .ZN(n128) );
  NOR2_X1 U211 ( .A1(n901), .A2(n120), .ZN(n798) );
  CLKBUF_X1 U212 ( .A(n798), .Z(n766) );
  NOR2_X1 U213 ( .A1(n120), .A2(n117), .ZN(n545) );
  AOI22_X1 U214 ( .A1(n766), .A2(hwlp_end_i[63]), .B1(n545), .B2(
        hwlp_cnt_i[31]), .ZN(n126) );
  NAND2_X1 U215 ( .A1(n116), .A2(n1371), .ZN(n893) );
  NOR2_X1 U216 ( .A1(n152), .A2(n893), .ZN(n279) );
  CLKBUF_X1 U217 ( .A(n279), .Z(n783) );
  NOR2_X1 U218 ( .A1(csr_addr_i[11]), .A2(n71), .ZN(n1029) );
  AOI22_X1 U219 ( .A1(n783), .A2(dscratch1_q[31]), .B1(n1029), .B2(mcause_q[5]), .ZN(n125) );
  NAND2_X1 U220 ( .A1(n121), .A2(n1370), .ZN(n243) );
  NOR2_X1 U221 ( .A1(csr_addr_i[11]), .A2(n243), .ZN(n179) );
  CLKBUF_X1 U222 ( .A(n179), .Z(n748) );
  NAND2_X1 U223 ( .A1(n119), .A2(n909), .ZN(n897) );
  NOR2_X1 U224 ( .A1(n120), .A2(n897), .ZN(n137) );
  CLKBUF_X1 U225 ( .A(n137), .Z(n799) );
  AOI22_X1 U226 ( .A1(n748), .A2(n18), .B1(n799), .B2(hwlp_start_i[63]), .ZN(
        n124) );
  NAND2_X1 U227 ( .A1(n121), .A2(n1371), .ZN(n174) );
  NOR2_X1 U228 ( .A1(csr_addr_i[11]), .A2(n174), .ZN(n181) );
  CLKBUF_X1 U229 ( .A(n181), .Z(n642) );
  INV_X1 U230 ( .A(n146), .ZN(n353) );
  INV_X1 U231 ( .A(n1429), .ZN(n1375) );
  NOR2_X1 U232 ( .A1(csr_addr_i[11]), .A2(n1375), .ZN(n350) );
  INV_X1 U233 ( .A(n350), .ZN(n714) );
  AOI22_X1 U235 ( .A1(n642), .A2(n6), .B1(n734), .B2(mtvec_o[23]), .ZN(n123)
         );
  NAND4_X1 U236 ( .A1(n126), .A2(n125), .A3(n124), .A4(n123), .ZN(n127) );
  OR3_X1 U237 ( .A1(n129), .A2(n128), .A3(n127), .ZN(csr_rdata_o[31]) );
  NAND2_X1 U238 ( .A1(csr_op_i[1]), .A2(csr_rdata_o[31]), .ZN(n131) );
  NAND2_X1 U239 ( .A1(csr_wdata_i[31]), .A2(n1362), .ZN(n130) );
  INV_X1 U242 ( .A(n132), .ZN(n195) );
  INV_X1 U244 ( .A(n911), .ZN(n134) );
  CLKBUF_X1 U247 ( .A(n716), .Z(n782) );
  AOI22_X1 U248 ( .A1(n782), .A2(hwlp_end_i[8]), .B1(n715), .B2(depc_o[8]), 
        .ZN(n145) );
  AOI22_X1 U249 ( .A1(n65), .A2(mepc_o[8]), .B1(n696), .B2(hwlp_start_i[8]), 
        .ZN(n144) );
  AOI22_X1 U250 ( .A1(n783), .A2(dscratch1_q[8]), .B1(n695), .B2(
        dscratch0_q[8]), .ZN(n143) );
  NAND2_X1 U251 ( .A1(csr_addr_i[4]), .A2(n138), .ZN(n673) );
  AOI21_X1 U252 ( .B1(n3700), .B2(n139), .A(n897), .ZN(n140) );
  INV_X1 U253 ( .A(n140), .ZN(n141) );
  AOI22_X1 U254 ( .A1(n799), .A2(hwlp_start_i[40]), .B1(n761), .B2(
        cluster_id_i[3]), .ZN(n142) );
  INV_X2 U256 ( .A(n647), .ZN(n1380) );
  AOI22_X1 U257 ( .A1(n766), .A2(hwlp_end_i[40]), .B1(n801), .B2(uepc_o[8]), 
        .ZN(n147) );
  NAND3_X1 U258 ( .A1(n146), .A2(n886), .A3(n3700), .ZN(n643) );
  OAI211_X1 U259 ( .C1(n1240), .C2(n1463), .A(n147), .B(n643), .ZN(n148) );
  AOI21_X1 U260 ( .B1(n1380), .B2(utvec_o[0]), .A(n148), .ZN(n165) );
  AOI22_X1 U261 ( .A1(n642), .A2(pmp_cfg_o[104]), .B1(n350), .B2(mtvec_o[0]), 
        .ZN(n151) );
  AOI22_X1 U262 ( .A1(n690), .A2(hwlp_cnt_i[40]), .B1(n760), .B2(hwlp_cnt_i[8]), .ZN(n150) );
  NAND2_X1 U263 ( .A1(n748), .A2(pmp_cfg_o[72]), .ZN(n149) );
  AND3_X1 U264 ( .A1(n151), .A2(n150), .A3(n149), .ZN(n164) );
  NOR2_X1 U265 ( .A1(n152), .A2(n881), .ZN(n609) );
  CLKBUF_X1 U266 ( .A(n609), .Z(n735) );
  AOI22_X1 U267 ( .A1(n735), .A2(dcsr_q_cause__8_), .B1(n691), .B2(
        mscratch_q[8]), .ZN(n163) );
  INV_X1 U268 ( .A(n154), .ZN(n158) );
  NOR2_X1 U269 ( .A1(csr_addr_i[9]), .A2(csr_addr_i[8]), .ZN(n155) );
  NAND3_X1 U270 ( .A1(csr_addr_i[11]), .A2(csr_addr_i[10]), .A3(n155), .ZN(
        n672) );
  AOI221_X1 U271 ( .B1(csr_addr_i[5]), .B2(n158), .C1(n157), .C2(n672), .A(
        n156), .ZN(n159) );
  NAND2_X1 U272 ( .A1(n1715), .A2(n159), .ZN(n678) );
  NOR2_X2 U273 ( .A1(n881), .A2(n678), .ZN(n788) );
  NAND2_X1 U274 ( .A1(n800), .A2(pmp_cfg_o[40]), .ZN(n160) );
  OAI21_X1 U275 ( .B1(n551), .B2(n1607), .A(n160), .ZN(n161) );
  AOI21_X1 U276 ( .B1(n788), .B2(PCER_q[8]), .A(n161), .ZN(n162) );
  INV_X1 U279 ( .A(csr_wdata_i[8]), .ZN(n170) );
  NOR2_X1 U280 ( .A1(n708), .A2(csr_wdata_i[8]), .ZN(n168) );
  NAND2_X1 U281 ( .A1(csr_rdata_o[8]), .A2(n168), .ZN(n169) );
  OAI21_X1 U282 ( .B1(n170), .B2(n1257), .A(n169), .ZN(hwlp_data_o[8]) );
  AOI22_X1 U290 ( .A1(n783), .A2(dscratch1_q[25]), .B1(n548), .B2(uepc_o[25]), 
        .ZN(n178) );
  AOI22_X1 U291 ( .A1(n799), .A2(hwlp_start_i[57]), .B1(n410), .B2(
        dscratch0_q[25]), .ZN(n177) );
  AOI22_X1 U292 ( .A1(n782), .A2(hwlp_end_i[25]), .B1(n696), .B2(
        hwlp_start_i[25]), .ZN(n176) );
  AND3_X1 U293 ( .A1(n178), .A2(n177), .A3(n176), .ZN(n185) );
  AOI22_X1 U294 ( .A1(n1380), .A2(utvec_o[17]), .B1(n734), .B2(mtvec_o[17]), 
        .ZN(n184) );
  AOI22_X1 U295 ( .A1(n748), .A2(pmp_cfg_o[89]), .B1(n800), .B2(pmp_cfg_o[57]), 
        .ZN(n183) );
  AOI22_X1 U296 ( .A1(n181), .A2(pmp_cfg_o[121]), .B1(n767), .B2(pmp_cfg_o[25]), .ZN(n182) );
  AND4_X1 U297 ( .A1(n185), .A2(n184), .A3(n183), .A4(n182), .ZN(n191) );
  AOI22_X1 U298 ( .A1(n790), .A2(PCCR_q[25]), .B1(n735), .B2(dcsr_q_zero2__25_), .ZN(n189) );
  AOI22_X1 U299 ( .A1(n691), .A2(mscratch_q[25]), .B1(n690), .B2(
        hwlp_cnt_i[57]), .ZN(n188) );
  AOI22_X1 U300 ( .A1(n766), .A2(hwlp_end_i[57]), .B1(n701), .B2(depc_o[25]), 
        .ZN(n187) );
  AOI22_X1 U301 ( .A1(n582), .A2(mepc_o[25]), .B1(n760), .B2(hwlp_cnt_i[25]), 
        .ZN(n186) );
  AND4_X1 U302 ( .A1(n189), .A2(n188), .A3(n187), .A4(n186), .ZN(n190) );
  NAND2_X1 U303 ( .A1(n191), .A2(n190), .ZN(csr_rdata_o[25]) );
  NAND3_X1 U304 ( .A1(csr_rdata_o[25]), .A2(csr_op_i[1]), .A3(n193), .ZN(n192)
         );
  OAI21_X2 U305 ( .B1(n193), .B2(n1257), .A(n192), .ZN(hwlp_data_o[25]) );
  NOR3_X1 U308 ( .A1(csr_addr_i[3]), .A2(n196), .A3(n195), .ZN(n1373) );
  NAND2_X1 U309 ( .A1(n914), .A2(n1373), .ZN(n197) );
  NOR2_X1 U310 ( .A1(n1198), .A2(n197), .ZN(n198) );
  AOI22_X1 U313 ( .A1(n279), .A2(dscratch1_q[24]), .B1(n548), .B2(uepc_o[24]), 
        .ZN(n203) );
  AOI22_X1 U314 ( .A1(n179), .A2(pmp_cfg_o[88]), .B1(n1380), .B2(utvec_o[16]), 
        .ZN(n202) );
  AOI22_X1 U315 ( .A1(n181), .A2(pmp_cfg_o[120]), .B1(n180), .B2(pmp_cfg_o[56]), .ZN(n201) );
  NAND2_X1 U316 ( .A1(n350), .A2(mtvec_o[16]), .ZN(n200) );
  AND4_X1 U317 ( .A1(n203), .A2(n202), .A3(n201), .A4(n200), .ZN(n213) );
  AOI22_X1 U318 ( .A1(n790), .A2(PCCR_q[24]), .B1(n760), .B2(hwlp_cnt_i[24]), 
        .ZN(n207) );
  AOI22_X1 U319 ( .A1(n690), .A2(hwlp_cnt_i[56]), .B1(n766), .B2(
        hwlp_end_i[56]), .ZN(n206) );
  AOI22_X1 U320 ( .A1(n799), .A2(hwlp_start_i[56]), .B1(n696), .B2(
        hwlp_start_i[24]), .ZN(n205) );
  AOI22_X1 U321 ( .A1(n782), .A2(hwlp_end_i[24]), .B1(n701), .B2(depc_o[24]), 
        .ZN(n204) );
  AND4_X1 U322 ( .A1(n207), .A2(n206), .A3(n205), .A4(n204), .ZN(n212) );
  AOI22_X1 U323 ( .A1(n691), .A2(mscratch_q[24]), .B1(n65), .B2(mepc_o[24]), 
        .ZN(n211) );
  AOI22_X1 U324 ( .A1(n609), .A2(dcsr_q_zero2__24_), .B1(n695), .B2(
        dscratch0_q[24]), .ZN(n209) );
  NAND2_X1 U325 ( .A1(n767), .A2(pmp_cfg_o[24]), .ZN(n208) );
  AND2_X1 U326 ( .A1(n209), .A2(n208), .ZN(n210) );
  NAND4_X1 U327 ( .A1(n213), .A2(n212), .A3(n211), .A4(n210), .ZN(
        csr_rdata_o[24]) );
  INV_X1 U328 ( .A(csr_wdata_i[24]), .ZN(n214) );
  NAND3_X1 U329 ( .A1(csr_rdata_o[24]), .A2(csr_op_i[1]), .A3(n214), .ZN(n216)
         );
  NAND2_X1 U330 ( .A1(csr_wdata_i[24]), .A2(n1362), .ZN(n215) );
  NAND2_X1 U331 ( .A1(n216), .A2(n215), .ZN(hwlp_data_o[24]) );
  NAND2_X1 U336 ( .A1(csr_addr_i[2]), .A2(n923), .ZN(n936) );
  NOR2_X1 U337 ( .A1(n1224), .A2(n936), .ZN(n928) );
  NOR2_X1 U342 ( .A1(n1223), .A2(n936), .ZN(n926) );
  NOR2_X1 U347 ( .A1(n1226), .A2(n936), .ZN(n932) );
  AOI22_X1 U352 ( .A1(n790), .A2(PCCR_q[10]), .B1(n782), .B2(hwlp_end_i[10]), 
        .ZN(n226) );
  AOI22_X1 U353 ( .A1(n642), .A2(pmp_cfg_o[106]), .B1(n800), .B2(pmp_cfg_o[42]), .ZN(n225) );
  OAI211_X1 U354 ( .C1(n551), .C2(n1478), .A(n226), .B(n225), .ZN(n237) );
  AOI22_X1 U355 ( .A1(n548), .A2(uepc_o[10]), .B1(n761), .B2(cluster_id_i[5]), 
        .ZN(n230) );
  AOI22_X1 U356 ( .A1(n65), .A2(mepc_o[10]), .B1(n783), .B2(dscratch1_q[10]), 
        .ZN(n229) );
  AOI22_X1 U357 ( .A1(n691), .A2(mscratch_q[10]), .B1(n798), .B2(
        hwlp_end_i[42]), .ZN(n228) );
  CLKBUF_X1 U358 ( .A(n545), .Z(n760) );
  AOI22_X1 U359 ( .A1(n696), .A2(hwlp_start_i[10]), .B1(n760), .B2(
        hwlp_cnt_i[10]), .ZN(n227) );
  NAND4_X1 U360 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(n236) );
  AOI22_X1 U361 ( .A1(n799), .A2(hwlp_start_i[42]), .B1(n641), .B2(
        hwlp_cnt_i[42]), .ZN(n234) );
  AOI22_X1 U362 ( .A1(n695), .A2(dscratch0_q[10]), .B1(n701), .B2(depc_o[10]), 
        .ZN(n233) );
  AOI22_X1 U363 ( .A1(n748), .A2(pmp_cfg_o[74]), .B1(n788), .B2(PCER_q[10]), 
        .ZN(n232) );
  AOI22_X1 U364 ( .A1(n1380), .A2(utvec_o[2]), .B1(n350), .B2(mtvec_o[2]), 
        .ZN(n231) );
  NAND4_X1 U365 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(n235) );
  OR3_X1 U366 ( .A1(n237), .A2(n236), .A3(n235), .ZN(csr_rdata_o[10]) );
  NAND2_X1 U367 ( .A1(n814), .A2(csr_rdata_o[10]), .ZN(n239) );
  NAND2_X1 U368 ( .A1(csr_wdata_i[10]), .A2(n1362), .ZN(n238) );
  OAI21_X2 U369 ( .B1(n239), .B2(csr_wdata_i[10]), .A(n238), .ZN(
        hwlp_data_o[10]) );
  OR2_X1 U374 ( .A1(n243), .A2(n1198), .ZN(n865) );
  AOI22_X1 U378 ( .A1(n790), .A2(PCCR_q[19]), .B1(n690), .B2(hwlp_cnt_i[51]), 
        .ZN(n248) );
  AOI22_X1 U379 ( .A1(n609), .A2(dcsr_q_zero2__19_), .B1(n799), .B2(
        hwlp_start_i[51]), .ZN(n247) );
  AOI22_X1 U380 ( .A1(n783), .A2(dscratch1_q[19]), .B1(n715), .B2(depc_o[19]), 
        .ZN(n246) );
  AOI22_X1 U381 ( .A1(n691), .A2(mscratch_q[19]), .B1(n801), .B2(uepc_o[19]), 
        .ZN(n245) );
  AND4_X1 U382 ( .A1(n248), .A2(n247), .A3(n246), .A4(n245), .ZN(n258) );
  AOI22_X1 U383 ( .A1(n642), .A2(pmp_cfg_o[115]), .B1(n800), .B2(pmp_cfg_o[51]), .ZN(n257) );
  AOI22_X1 U384 ( .A1(n782), .A2(hwlp_end_i[19]), .B1(n695), .B2(
        dscratch0_q[19]), .ZN(n250) );
  NAND2_X1 U385 ( .A1(n767), .A2(pmp_cfg_o[19]), .ZN(n249) );
  AND2_X1 U386 ( .A1(n250), .A2(n249), .ZN(n256) );
  AOI22_X1 U387 ( .A1(n582), .A2(mepc_o[19]), .B1(n766), .B2(hwlp_end_i[51]), 
        .ZN(n254) );
  AOI22_X1 U388 ( .A1(n696), .A2(hwlp_start_i[19]), .B1(n760), .B2(
        hwlp_cnt_i[19]), .ZN(n253) );
  NAND2_X1 U389 ( .A1(n734), .A2(mtvec_o[11]), .ZN(n252) );
  AOI22_X1 U390 ( .A1(n179), .A2(pmp_cfg_o[83]), .B1(n1380), .B2(utvec_o[11]), 
        .ZN(n251) );
  AND4_X1 U391 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(n255) );
  NAND4_X1 U392 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(
        csr_rdata_o[19]) );
  INV_X1 U393 ( .A(csr_wdata_i[19]), .ZN(n259) );
  NAND3_X1 U394 ( .A1(csr_rdata_o[19]), .A2(csr_op_i[1]), .A3(n259), .ZN(n261)
         );
  NAND2_X1 U395 ( .A1(csr_wdata_i[19]), .A2(n1362), .ZN(n260) );
  NAND2_X1 U396 ( .A1(n261), .A2(n260), .ZN(hwlp_data_o[19]) );
  AOI22_X1 U399 ( .A1(n790), .A2(PCCR_q[27]), .B1(n766), .B2(hwlp_end_i[59]), 
        .ZN(n266) );
  AOI22_X1 U400 ( .A1(n695), .A2(dscratch0_q[27]), .B1(n548), .B2(uepc_o[27]), 
        .ZN(n265) );
  AOI22_X1 U401 ( .A1(n783), .A2(dscratch1_q[27]), .B1(n799), .B2(
        hwlp_start_i[59]), .ZN(n264) );
  AOI22_X1 U402 ( .A1(n782), .A2(hwlp_end_i[27]), .B1(n701), .B2(depc_o[27]), 
        .ZN(n263) );
  AND4_X1 U403 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(n274) );
  AOI22_X1 U404 ( .A1(n609), .A2(dcsr_q_zero2__27_), .B1(n65), .B2(mepc_o[27]), 
        .ZN(n270) );
  AOI22_X1 U405 ( .A1(n696), .A2(hwlp_start_i[27]), .B1(n690), .B2(
        hwlp_cnt_i[59]), .ZN(n269) );
  AOI22_X1 U406 ( .A1(n179), .A2(pmp_cfg_o[91]), .B1(n1380), .B2(utvec_o[19]), 
        .ZN(n268) );
  AOI22_X1 U407 ( .A1(n181), .A2(pmp_cfg_o[123]), .B1(n180), .B2(pmp_cfg_o[59]), .ZN(n267) );
  AND4_X1 U408 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(n273) );
  AOI22_X1 U409 ( .A1(n691), .A2(mscratch_q[27]), .B1(n760), .B2(
        hwlp_cnt_i[27]), .ZN(n272) );
  AOI22_X1 U410 ( .A1(n734), .A2(mtvec_o[19]), .B1(n767), .B2(pmp_cfg_o[27]), 
        .ZN(n271) );
  NAND4_X1 U411 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(
        csr_rdata_o[27]) );
  INV_X1 U412 ( .A(csr_wdata_i[27]), .ZN(n275) );
  NAND3_X1 U413 ( .A1(csr_rdata_o[27]), .A2(csr_op_i[1]), .A3(n275), .ZN(n277)
         );
  NAND2_X1 U414 ( .A1(n277), .A2(n276), .ZN(hwlp_data_o[27]) );
  AOI22_X1 U417 ( .A1(n767), .A2(n46), .B1(n734), .B2(mtvec_o[14]), .ZN(n291)
         );
  AOI22_X1 U418 ( .A1(n748), .A2(n22), .B1(n1380), .B2(utvec_o[14]), .ZN(n290)
         );
  AOI22_X1 U419 ( .A1(n790), .A2(PCCR_q[22]), .B1(n641), .B2(hwlp_cnt_i[54]), 
        .ZN(n283) );
  AOI22_X1 U420 ( .A1(n695), .A2(dscratch0_q[22]), .B1(n798), .B2(
        hwlp_end_i[54]), .ZN(n282) );
  AOI22_X1 U421 ( .A1(n582), .A2(mepc_o[22]), .B1(n799), .B2(hwlp_start_i[54]), 
        .ZN(n281) );
  AOI22_X1 U422 ( .A1(n716), .A2(hwlp_end_i[22]), .B1(n279), .B2(
        dscratch1_q[22]), .ZN(n280) );
  AND4_X1 U423 ( .A1(n283), .A2(n282), .A3(n281), .A4(n280), .ZN(n289) );
  AOI22_X1 U424 ( .A1(n735), .A2(dcsr_q_zero2__22_), .B1(n701), .B2(depc_o[22]), .ZN(n287) );
  AOI22_X1 U425 ( .A1(n696), .A2(hwlp_start_i[22]), .B1(n760), .B2(
        hwlp_cnt_i[22]), .ZN(n286) );
  AOI22_X1 U426 ( .A1(n691), .A2(mscratch_q[22]), .B1(n548), .B2(uepc_o[22]), 
        .ZN(n285) );
  AOI22_X1 U427 ( .A1(n642), .A2(n10), .B1(n800), .B2(n34), .ZN(n284) );
  AND4_X1 U428 ( .A1(n287), .A2(n286), .A3(n285), .A4(n284), .ZN(n288) );
  NAND4_X1 U429 ( .A1(n291), .A2(n290), .A3(n289), .A4(n288), .ZN(
        csr_rdata_o[22]) );
  AOI21_X1 U430 ( .B1(csr_op_i[1]), .B2(csr_rdata_o[22]), .A(csr_wdata_i[22]), 
        .ZN(n292) );
  OAI22_X1 U431 ( .A1(n865), .A2(n1007), .B1(n22), .B2(n3966), .ZN(n293) );
  INV_X1 U432 ( .A(n293), .ZN(n2068) );
  AOI22_X1 U435 ( .A1(n701), .A2(depc_o[20]), .B1(n801), .B2(uepc_o[20]), .ZN(
        n298) );
  AOI22_X1 U436 ( .A1(n690), .A2(hwlp_cnt_i[52]), .B1(n798), .B2(
        hwlp_end_i[52]), .ZN(n297) );
  AOI22_X1 U437 ( .A1(n609), .A2(dcsr_q_zero2__20_), .B1(n691), .B2(
        mscratch_q[20]), .ZN(n296) );
  AOI22_X1 U438 ( .A1(n783), .A2(dscratch1_q[20]), .B1(n695), .B2(
        dscratch0_q[20]), .ZN(n295) );
  NAND4_X1 U439 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(n303) );
  AOI22_X1 U440 ( .A1(n179), .A2(pmp_cfg_o[84]), .B1(n767), .B2(pmp_cfg_o[20]), 
        .ZN(n301) );
  AOI22_X1 U441 ( .A1(n716), .A2(hwlp_end_i[20]), .B1(n760), .B2(
        hwlp_cnt_i[20]), .ZN(n300) );
  NAND2_X1 U442 ( .A1(n734), .A2(mtvec_o[12]), .ZN(n299) );
  NAND3_X1 U443 ( .A1(n301), .A2(n300), .A3(n299), .ZN(n302) );
  NOR2_X1 U444 ( .A1(n303), .A2(n302), .ZN(n309) );
  AOI22_X1 U445 ( .A1(n799), .A2(hwlp_start_i[52]), .B1(n696), .B2(
        hwlp_start_i[20]), .ZN(n308) );
  AOI22_X1 U446 ( .A1(n800), .A2(pmp_cfg_o[52]), .B1(pmp_cfg_o[116]), .B2(n642), .ZN(n307) );
  AOI22_X1 U447 ( .A1(n1380), .A2(utvec_o[12]), .B1(n65), .B2(mepc_o[20]), 
        .ZN(n304) );
  OAI211_X1 U448 ( .C1(n1240), .C2(n1464), .A(n304), .B(n643), .ZN(n305) );
  INV_X1 U449 ( .A(n305), .ZN(n306) );
  NAND4_X1 U450 ( .A1(n309), .A2(n308), .A3(n307), .A4(n306), .ZN(
        csr_rdata_o[20]) );
  INV_X1 U451 ( .A(csr_wdata_i[20]), .ZN(n310) );
  NAND3_X1 U452 ( .A1(csr_rdata_o[20]), .A2(csr_op_i[1]), .A3(n310), .ZN(n312)
         );
  NAND2_X1 U453 ( .A1(n312), .A2(n311), .ZN(hwlp_data_o[20]) );
  AOI22_X1 U456 ( .A1(n642), .A2(n17), .B1(n767), .B2(n53), .ZN(n325) );
  AOI22_X1 U457 ( .A1(n800), .A2(n41), .B1(n788), .B2(PCER_q[5]), .ZN(n324) );
  AOI22_X1 U458 ( .A1(n790), .A2(PCCR_q[5]), .B1(n761), .B2(cluster_id_i[0]), 
        .ZN(n317) );
  AOI22_X1 U459 ( .A1(n137), .A2(hwlp_start_i[37]), .B1(n715), .B2(depc_o[5]), 
        .ZN(n316) );
  AOI22_X1 U460 ( .A1(n782), .A2(hwlp_end_i[5]), .B1(n783), .B2(dscratch1_q[5]), .ZN(n315) );
  AOI22_X1 U461 ( .A1(n153), .A2(mscratch_q[5]), .B1(n798), .B2(hwlp_end_i[37]), .ZN(n314) );
  AND4_X1 U462 ( .A1(n317), .A2(n316), .A3(n315), .A4(n314), .ZN(n323) );
  AOI22_X1 U463 ( .A1(n65), .A2(mepc_o[5]), .B1(n641), .B2(hwlp_cnt_i[37]), 
        .ZN(n321) );
  AOI22_X1 U464 ( .A1(n695), .A2(dscratch0_q[5]), .B1(n545), .B2(hwlp_cnt_i[5]), .ZN(n320) );
  AOI22_X1 U465 ( .A1(n735), .A2(dcsr_q_zero0_), .B1(n801), .B2(uepc_o[5]), 
        .ZN(n319) );
  AOI22_X1 U466 ( .A1(n748), .A2(n29), .B1(n136), .B2(hwlp_start_i[5]), .ZN(
        n318) );
  AND4_X1 U467 ( .A1(n321), .A2(n320), .A3(n319), .A4(n318), .ZN(n322) );
  NAND4_X1 U468 ( .A1(n325), .A2(n324), .A3(n323), .A4(n322), .ZN(
        csr_rdata_o[5]) );
  AOI21_X1 U469 ( .B1(csr_op_i[1]), .B2(csr_rdata_o[5]), .A(csr_wdata_i[5]), 
        .ZN(n326) );
  OAI22_X1 U472 ( .A1(n1446), .A2(n970), .B1(n17), .B2(n3969), .ZN(n328) );
  INV_X1 U473 ( .A(n328), .ZN(n2051) );
  AOI22_X1 U474 ( .A1(n734), .A2(mtvec_o[8]), .B1(n767), .B2(pmp_cfg_o[16]), 
        .ZN(n331) );
  AOI22_X1 U475 ( .A1(n799), .A2(hwlp_start_i[48]), .B1(n641), .B2(
        hwlp_cnt_i[48]), .ZN(n330) );
  AOI22_X1 U476 ( .A1(n582), .A2(mepc_o[16]), .B1(n783), .B2(dscratch1_q[16]), 
        .ZN(n329) );
  AND3_X1 U477 ( .A1(n331), .A2(n330), .A3(n329), .ZN(n341) );
  AOI22_X1 U478 ( .A1(n790), .A2(PCCR_q[16]), .B1(n782), .B2(hwlp_end_i[16]), 
        .ZN(n335) );
  AOI22_X1 U479 ( .A1(n609), .A2(dcsr_q_zero2__16_), .B1(n695), .B2(
        dscratch0_q[16]), .ZN(n334) );
  AOI22_X1 U480 ( .A1(n766), .A2(hwlp_end_i[48]), .B1(n715), .B2(depc_o[16]), 
        .ZN(n333) );
  AOI22_X1 U481 ( .A1(n696), .A2(hwlp_start_i[16]), .B1(n760), .B2(
        hwlp_cnt_i[16]), .ZN(n332) );
  AND4_X1 U482 ( .A1(n335), .A2(n334), .A3(n333), .A4(n332), .ZN(n340) );
  AOI22_X1 U483 ( .A1(n691), .A2(mscratch_q[16]), .B1(n801), .B2(uepc_o[16]), 
        .ZN(n339) );
  AOI22_X1 U484 ( .A1(n181), .A2(pmp_cfg_o[112]), .B1(n180), .B2(pmp_cfg_o[48]), .ZN(n337) );
  AOI22_X1 U485 ( .A1(n179), .A2(pmp_cfg_o[80]), .B1(n1380), .B2(utvec_o[8]), 
        .ZN(n336) );
  AND2_X1 U486 ( .A1(n337), .A2(n336), .ZN(n338) );
  NAND4_X1 U487 ( .A1(n341), .A2(n340), .A3(n339), .A4(n338), .ZN(
        csr_rdata_o[16]) );
  INV_X1 U488 ( .A(csr_wdata_i[16]), .ZN(n342) );
  NAND3_X1 U489 ( .A1(csr_rdata_o[16]), .A2(csr_op_i[1]), .A3(n342), .ZN(n344)
         );
  NAND2_X1 U490 ( .A1(csr_wdata_i[16]), .A2(n1362), .ZN(n343) );
  AND2_X1 U491 ( .A1(n344), .A2(n343), .ZN(n1409) );
  AOI22_X1 U495 ( .A1(n696), .A2(hwlp_start_i[12]), .B1(n801), .B2(uepc_o[12]), 
        .ZN(n349) );
  AOI22_X1 U496 ( .A1(n735), .A2(debug_ebreaku_o), .B1(n279), .B2(
        dscratch1_q[12]), .ZN(n348) );
  AOI22_X1 U497 ( .A1(n799), .A2(hwlp_start_i[44]), .B1(n690), .B2(
        hwlp_cnt_i[44]), .ZN(n347) );
  AOI22_X1 U498 ( .A1(n716), .A2(hwlp_end_i[12]), .B1(n695), .B2(
        dscratch0_q[12]), .ZN(n346) );
  AND4_X1 U499 ( .A1(n349), .A2(n348), .A3(n347), .A4(n346), .ZN(n365) );
  AOI22_X1 U500 ( .A1(n65), .A2(mepc_o[12]), .B1(n798), .B2(hwlp_end_i[44]), 
        .ZN(n352) );
  NAND2_X1 U501 ( .A1(n350), .A2(mtvec_o[4]), .ZN(n351) );
  NAND2_X1 U502 ( .A1(n352), .A2(n351), .ZN(n359) );
  NAND2_X1 U503 ( .A1(n743), .A2(n3700), .ZN(n506) );
  INV_X1 U504 ( .A(n506), .ZN(n770) );
  AOI22_X1 U505 ( .A1(n770), .A2(mstatus_q[2]), .B1(n1380), .B2(utvec_o[4]), 
        .ZN(n357) );
  NAND2_X1 U506 ( .A1(n179), .A2(pmp_cfg_o[76]), .ZN(n356) );
  NAND2_X1 U507 ( .A1(n800), .A2(pmp_cfg_o[44]), .ZN(n355) );
  NAND2_X1 U508 ( .A1(n642), .A2(pmp_cfg_o[108]), .ZN(n354) );
  NAND4_X1 U509 ( .A1(n357), .A2(n356), .A3(n355), .A4(n354), .ZN(n358) );
  NOR2_X1 U510 ( .A1(n359), .A2(n358), .ZN(n364) );
  AOI22_X1 U511 ( .A1(n701), .A2(depc_o[12]), .B1(n545), .B2(hwlp_cnt_i[12]), 
        .ZN(n360) );
  OAI211_X1 U512 ( .C1(n1240), .C2(n1462), .A(n360), .B(n643), .ZN(n361) );
  INV_X1 U513 ( .A(n361), .ZN(n363) );
  AOI22_X1 U514 ( .A1(n691), .A2(mscratch_q[12]), .B1(n767), .B2(pmp_cfg_o[12]), .ZN(n362) );
  NAND4_X1 U515 ( .A1(n365), .A2(n364), .A3(n363), .A4(n362), .ZN(
        csr_rdata_o[12]) );
  NOR2_X1 U516 ( .A1(n708), .A2(csr_wdata_i[12]), .ZN(n366) );
  NAND2_X1 U517 ( .A1(csr_rdata_o[12]), .A2(n366), .ZN(n368) );
  NAND2_X1 U518 ( .A1(csr_wdata_i[12]), .A2(n1362), .ZN(n367) );
  AND2_X1 U519 ( .A1(n368), .A2(n367), .ZN(n1405) );
  AOI22_X1 U525 ( .A1(n642), .A2(pmp_cfg_o[114]), .B1(n1380), .B2(utvec_o[10]), 
        .ZN(n382) );
  AOI22_X1 U526 ( .A1(n800), .A2(pmp_cfg_o[50]), .B1(n734), .B2(mtvec_o[10]), 
        .ZN(n381) );
  AOI22_X1 U527 ( .A1(n790), .A2(PCCR_q[18]), .B1(n65), .B2(mepc_o[18]), .ZN(
        n374) );
  AOI22_X1 U528 ( .A1(n766), .A2(hwlp_end_i[50]), .B1(n715), .B2(depc_o[18]), 
        .ZN(n373) );
  AOI22_X1 U529 ( .A1(n735), .A2(dcsr_q_zero2__18_), .B1(n799), .B2(
        hwlp_start_i[50]), .ZN(n372) );
  AOI22_X1 U530 ( .A1(n782), .A2(hwlp_end_i[18]), .B1(n801), .B2(uepc_o[18]), 
        .ZN(n371) );
  AND4_X1 U531 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(n380) );
  AOI22_X1 U532 ( .A1(n691), .A2(mscratch_q[18]), .B1(n696), .B2(
        hwlp_start_i[18]), .ZN(n378) );
  AOI22_X1 U533 ( .A1(n695), .A2(dscratch0_q[18]), .B1(n690), .B2(
        hwlp_cnt_i[50]), .ZN(n377) );
  AOI22_X1 U534 ( .A1(n783), .A2(dscratch1_q[18]), .B1(n760), .B2(
        hwlp_cnt_i[18]), .ZN(n376) );
  AOI22_X1 U535 ( .A1(n767), .A2(pmp_cfg_o[18]), .B1(n748), .B2(pmp_cfg_o[82]), 
        .ZN(n375) );
  AND4_X1 U536 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(n379) );
  NAND4_X1 U537 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(
        csr_rdata_o[18]) );
  NAND2_X1 U538 ( .A1(n814), .A2(csr_rdata_o[18]), .ZN(n384) );
  NAND2_X1 U539 ( .A1(csr_wdata_i[18]), .A2(n1362), .ZN(n383) );
  OR2_X1 U544 ( .A1(n387), .A2(n1198), .ZN(n1443) );
  INV_X1 U545 ( .A(n1443), .ZN(n1445) );
  AOI22_X1 U550 ( .A1(n800), .A2(pmp_cfg_o[58]), .B1(n748), .B2(pmp_cfg_o[90]), 
        .ZN(n401) );
  AOI22_X1 U551 ( .A1(n642), .A2(pmp_cfg_o[122]), .B1(n767), .B2(pmp_cfg_o[26]), .ZN(n400) );
  AOI22_X1 U552 ( .A1(n790), .A2(PCCR_q[26]), .B1(n782), .B2(hwlp_end_i[26]), 
        .ZN(n393) );
  AOI22_X1 U553 ( .A1(n609), .A2(dcsr_q_zero2__26_), .B1(n701), .B2(depc_o[26]), .ZN(n392) );
  AOI22_X1 U554 ( .A1(n766), .A2(hwlp_end_i[58]), .B1(n801), .B2(uepc_o[26]), 
        .ZN(n391) );
  AOI22_X1 U555 ( .A1(n799), .A2(hwlp_start_i[58]), .B1(n410), .B2(
        dscratch0_q[26]), .ZN(n390) );
  AND4_X1 U556 ( .A1(n393), .A2(n392), .A3(n391), .A4(n390), .ZN(n399) );
  AOI22_X1 U557 ( .A1(n690), .A2(hwlp_cnt_i[58]), .B1(n760), .B2(
        hwlp_cnt_i[26]), .ZN(n397) );
  AOI22_X1 U558 ( .A1(n582), .A2(mepc_o[26]), .B1(n696), .B2(hwlp_start_i[26]), 
        .ZN(n396) );
  AOI22_X1 U559 ( .A1(n691), .A2(mscratch_q[26]), .B1(n279), .B2(
        dscratch1_q[26]), .ZN(n395) );
  AOI22_X1 U560 ( .A1(n1380), .A2(utvec_o[18]), .B1(n734), .B2(mtvec_o[18]), 
        .ZN(n394) );
  AND4_X1 U561 ( .A1(n397), .A2(n396), .A3(n395), .A4(n394), .ZN(n398) );
  NAND4_X1 U562 ( .A1(n401), .A2(n400), .A3(n399), .A4(n398), .ZN(
        csr_rdata_o[26]) );
  NAND2_X1 U563 ( .A1(n814), .A2(csr_rdata_o[26]), .ZN(n403) );
  NAND2_X1 U564 ( .A1(csr_wdata_i[26]), .A2(n1362), .ZN(n402) );
  OAI22_X1 U566 ( .A1(n864), .A2(n3955), .B1(pmp_cfg_o[58]), .B2(n241), .ZN(
        n404) );
  INV_X1 U567 ( .A(n404), .ZN(n2088) );
  OAI22_X1 U568 ( .A1(n865), .A2(n3955), .B1(pmp_cfg_o[90]), .B2(n3966), .ZN(
        n405) );
  INV_X1 U569 ( .A(n405), .ZN(n2056) );
  OAI22_X1 U570 ( .A1(n1443), .A2(n3955), .B1(pmp_cfg_o[26]), .B2(n1445), .ZN(
        n406) );
  INV_X1 U571 ( .A(n406), .ZN(n2120) );
  OAI22_X1 U572 ( .A1(n1446), .A2(n3955), .B1(pmp_cfg_o[122]), .B2(n3969), 
        .ZN(n407) );
  INV_X1 U573 ( .A(n407), .ZN(n2024) );
  AOI22_X1 U578 ( .A1(n642), .A2(n11), .B1(n800), .B2(n35), .ZN(n422) );
  AOI22_X1 U579 ( .A1(n1380), .A2(utvec_o[13]), .B1(n734), .B2(mtvec_o[13]), 
        .ZN(n421) );
  AOI22_X1 U580 ( .A1(n790), .A2(PCCR_q[21]), .B1(n735), .B2(dcsr_q_zero2__21_), .ZN(n414) );
  AOI22_X1 U581 ( .A1(n799), .A2(hwlp_start_i[53]), .B1(n701), .B2(depc_o[21]), 
        .ZN(n413) );
  AOI22_X1 U582 ( .A1(n691), .A2(mscratch_q[21]), .B1(n410), .B2(
        dscratch0_q[21]), .ZN(n412) );
  AOI22_X1 U583 ( .A1(n696), .A2(hwlp_start_i[21]), .B1(n641), .B2(
        hwlp_cnt_i[53]), .ZN(n411) );
  AND4_X1 U584 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(n420) );
  AOI22_X1 U585 ( .A1(n783), .A2(dscratch1_q[21]), .B1(n760), .B2(
        hwlp_cnt_i[21]), .ZN(n418) );
  AOI22_X1 U586 ( .A1(n766), .A2(hwlp_end_i[53]), .B1(n801), .B2(uepc_o[21]), 
        .ZN(n417) );
  AOI22_X1 U587 ( .A1(n782), .A2(hwlp_end_i[21]), .B1(n65), .B2(mepc_o[21]), 
        .ZN(n416) );
  AOI22_X1 U588 ( .A1(n767), .A2(n47), .B1(n748), .B2(n23), .ZN(n415) );
  AND4_X1 U589 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(n419) );
  NAND4_X1 U590 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(
        csr_rdata_o[21]) );
  NAND2_X1 U591 ( .A1(n814), .A2(csr_rdata_o[21]), .ZN(n424) );
  NAND2_X1 U592 ( .A1(csr_wdata_i[21]), .A2(n1362), .ZN(n423) );
  OAI22_X1 U598 ( .A1(n864), .A2(hwlp_data_o[21]), .B1(n35), .B2(n241), .ZN(
        n427) );
  INV_X1 U599 ( .A(n427), .ZN(n2099) );
  OAI22_X1 U600 ( .A1(n1446), .A2(hwlp_data_o[21]), .B1(n11), .B2(n3969), .ZN(
        n428) );
  INV_X1 U601 ( .A(n428), .ZN(n2035) );
  AOI22_X1 U602 ( .A1(n642), .A2(n13), .B1(n734), .B2(mtvec_o[6]), .ZN(n440)
         );
  AOI22_X1 U603 ( .A1(n800), .A2(n37), .B1(n767), .B2(n49), .ZN(n439) );
  AOI22_X1 U604 ( .A1(n790), .A2(PCCR_q[14]), .B1(n690), .B2(hwlp_cnt_i[46]), 
        .ZN(n432) );
  AOI22_X1 U605 ( .A1(n609), .A2(dcsr_q_zero1_), .B1(n701), .B2(depc_o[14]), 
        .ZN(n431) );
  AOI22_X1 U606 ( .A1(n582), .A2(mepc_o[14]), .B1(n801), .B2(uepc_o[14]), .ZN(
        n430) );
  AOI22_X1 U607 ( .A1(n153), .A2(mscratch_q[14]), .B1(n136), .B2(
        hwlp_start_i[14]), .ZN(n429) );
  AND4_X1 U608 ( .A1(n432), .A2(n431), .A3(n430), .A4(n429), .ZN(n438) );
  AOI22_X1 U609 ( .A1(n410), .A2(dscratch0_q[14]), .B1(n766), .B2(
        hwlp_end_i[46]), .ZN(n436) );
  AOI22_X1 U610 ( .A1(n783), .A2(dscratch1_q[14]), .B1(n137), .B2(
        hwlp_start_i[46]), .ZN(n435) );
  AOI22_X1 U611 ( .A1(n782), .A2(hwlp_end_i[14]), .B1(n760), .B2(
        hwlp_cnt_i[14]), .ZN(n434) );
  AOI22_X1 U612 ( .A1(n748), .A2(n25), .B1(n1380), .B2(utvec_o[6]), .ZN(n433)
         );
  AND4_X1 U613 ( .A1(n436), .A2(n435), .A3(n434), .A4(n433), .ZN(n437) );
  NAND4_X1 U614 ( .A1(n440), .A2(n439), .A3(n438), .A4(n437), .ZN(
        csr_rdata_o[14]) );
  NAND2_X1 U615 ( .A1(n814), .A2(csr_rdata_o[14]), .ZN(n442) );
  NAND2_X1 U616 ( .A1(csr_wdata_i[14]), .A2(n1362), .ZN(n441) );
  OAI21_X1 U617 ( .B1(n442), .B2(csr_wdata_i[14]), .A(n441), .ZN(n443) );
  INV_X1 U618 ( .A(n443), .ZN(n1407) );
  AOI22_X1 U631 ( .A1(n137), .A2(hwlp_start_i[43]), .B1(n696), .B2(
        hwlp_start_i[11]), .ZN(n453) );
  AOI22_X1 U632 ( .A1(n766), .A2(hwlp_end_i[43]), .B1(n545), .B2(
        hwlp_cnt_i[11]), .ZN(n452) );
  AOI22_X1 U633 ( .A1(n782), .A2(hwlp_end_i[11]), .B1(n609), .B2(
        dcsr_q_stepie_), .ZN(n451) );
  AOI22_X1 U634 ( .A1(n691), .A2(mscratch_q[11]), .B1(n410), .B2(
        dscratch0_q[11]), .ZN(n450) );
  NAND4_X1 U635 ( .A1(n453), .A2(n452), .A3(n451), .A4(n450), .ZN(n458) );
  AOI22_X1 U636 ( .A1(n734), .A2(mtvec_o[3]), .B1(mstatus_q[1]), .B2(n770), 
        .ZN(n456) );
  AOI22_X1 U637 ( .A1(n65), .A2(mepc_o[11]), .B1(n690), .B2(hwlp_cnt_i[43]), 
        .ZN(n455) );
  AOI22_X1 U638 ( .A1(n179), .A2(pmp_cfg_o[75]), .B1(utvec_o[3]), .B2(n1380), 
        .ZN(n454) );
  NAND3_X1 U639 ( .A1(n456), .A2(n455), .A3(n454), .ZN(n457) );
  NOR2_X1 U640 ( .A1(n458), .A2(n457), .ZN(n465) );
  AOI22_X1 U641 ( .A1(n783), .A2(dscratch1_q[11]), .B1(n548), .B2(uepc_o[11]), 
        .ZN(n464) );
  AOI22_X1 U642 ( .A1(n181), .A2(pmp_cfg_o[107]), .B1(n180), .B2(pmp_cfg_o[43]), .ZN(n463) );
  AOI22_X1 U643 ( .A1(n790), .A2(PCCR_q[11]), .B1(n701), .B2(depc_o[11]), .ZN(
        n460) );
  NAND2_X1 U644 ( .A1(n767), .A2(pmp_cfg_o[11]), .ZN(n459) );
  NAND2_X1 U645 ( .A1(n460), .A2(n459), .ZN(n461) );
  AOI21_X1 U646 ( .B1(n788), .B2(PCER_q[11]), .A(n461), .ZN(n462) );
  NAND4_X1 U647 ( .A1(n465), .A2(n464), .A3(n463), .A4(n462), .ZN(
        csr_rdata_o[11]) );
  INV_X1 U648 ( .A(csr_wdata_i[11]), .ZN(n466) );
  NAND3_X1 U649 ( .A1(csr_rdata_o[11]), .A2(csr_op_i[1]), .A3(n466), .ZN(n468)
         );
  NAND2_X1 U650 ( .A1(csr_wdata_i[11]), .A2(n1362), .ZN(n467) );
  AND2_X1 U651 ( .A1(n468), .A2(n467), .ZN(n1404) );
  AOI22_X1 U655 ( .A1(n767), .A2(n52), .B1(n788), .B2(PCER_q[6]), .ZN(n481) );
  AOI22_X1 U656 ( .A1(n642), .A2(n16), .B1(n800), .B2(n40), .ZN(n480) );
  AOI22_X1 U657 ( .A1(n790), .A2(PCCR_q[6]), .B1(n701), .B2(depc_o[6]), .ZN(
        n473) );
  AOI22_X1 U658 ( .A1(n153), .A2(mscratch_q[6]), .B1(n137), .B2(
        hwlp_start_i[38]), .ZN(n472) );
  AOI22_X1 U659 ( .A1(n690), .A2(hwlp_cnt_i[38]), .B1(n766), .B2(
        hwlp_end_i[38]), .ZN(n471) );
  AOI22_X1 U660 ( .A1(n735), .A2(dcsr_q_cause__6_), .B1(n783), .B2(
        dscratch1_q[6]), .ZN(n470) );
  AND4_X1 U661 ( .A1(n473), .A2(n472), .A3(n471), .A4(n470), .ZN(n479) );
  AOI22_X1 U662 ( .A1(n548), .A2(uepc_o[6]), .B1(n760), .B2(hwlp_cnt_i[6]), 
        .ZN(n477) );
  AOI22_X1 U663 ( .A1(n695), .A2(dscratch0_q[6]), .B1(n136), .B2(
        hwlp_start_i[6]), .ZN(n476) );
  AOI22_X1 U664 ( .A1(n716), .A2(hwlp_end_i[6]), .B1(n761), .B2(
        cluster_id_i[1]), .ZN(n475) );
  AOI22_X1 U665 ( .A1(n748), .A2(n28), .B1(n65), .B2(mepc_o[6]), .ZN(n474) );
  AND4_X1 U666 ( .A1(n477), .A2(n476), .A3(n475), .A4(n474), .ZN(n478) );
  NAND4_X1 U667 ( .A1(n481), .A2(n480), .A3(n479), .A4(n478), .ZN(
        csr_rdata_o[6]) );
  NAND3_X1 U668 ( .A1(csr_op_i[1]), .A2(csr_rdata_o[6]), .A3(n1256), .ZN(n482)
         );
  OAI21_X1 U669 ( .B1(n1256), .B2(n1257), .A(n482), .ZN(n483) );
  INV_X1 U670 ( .A(n483), .ZN(n1392) );
  AOI22_X1 U678 ( .A1(n642), .A2(n14), .B1(n734), .B2(mtvec_o[5]), .ZN(n498)
         );
  AOI22_X1 U679 ( .A1(n800), .A2(n38), .B1(n748), .B2(n26), .ZN(n497) );
  AOI22_X1 U680 ( .A1(n790), .A2(PCCR_q[13]), .B1(n782), .B2(hwlp_end_i[13]), 
        .ZN(n490) );
  AOI22_X1 U681 ( .A1(n153), .A2(mscratch_q[13]), .B1(n801), .B2(uepc_o[13]), 
        .ZN(n489) );
  AOI22_X1 U682 ( .A1(n735), .A2(dcsr_q_ebreaks_), .B1(n701), .B2(depc_o[13]), 
        .ZN(n488) );
  AOI22_X1 U683 ( .A1(n137), .A2(hwlp_start_i[45]), .B1(n410), .B2(
        dscratch0_q[13]), .ZN(n487) );
  AND4_X1 U684 ( .A1(n490), .A2(n489), .A3(n488), .A4(n487), .ZN(n496) );
  AOI22_X1 U685 ( .A1(n582), .A2(mepc_o[13]), .B1(n783), .B2(dscratch1_q[13]), 
        .ZN(n494) );
  AOI22_X1 U686 ( .A1(n690), .A2(hwlp_cnt_i[45]), .B1(n766), .B2(
        hwlp_end_i[45]), .ZN(n493) );
  AOI22_X1 U687 ( .A1(n136), .A2(hwlp_start_i[13]), .B1(n760), .B2(
        hwlp_cnt_i[13]), .ZN(n492) );
  AOI22_X1 U688 ( .A1(n767), .A2(n50), .B1(n1380), .B2(utvec_o[5]), .ZN(n491)
         );
  AND4_X1 U689 ( .A1(n494), .A2(n493), .A3(n492), .A4(n491), .ZN(n495) );
  NAND4_X1 U690 ( .A1(n498), .A2(n497), .A3(n496), .A4(n495), .ZN(
        csr_rdata_o[13]) );
  NAND2_X1 U691 ( .A1(n814), .A2(csr_rdata_o[13]), .ZN(n500) );
  NAND2_X1 U692 ( .A1(csr_wdata_i[13]), .A2(n1362), .ZN(n499) );
  OAI21_X1 U693 ( .B1(n500), .B2(csr_wdata_i[13]), .A(n499), .ZN(n501) );
  INV_X1 U694 ( .A(n501), .ZN(n1406) );
  AOI22_X1 U699 ( .A1(n790), .A2(PCCR_q[7]), .B1(n801), .B2(uepc_o[7]), .ZN(
        n505) );
  AOI22_X1 U700 ( .A1(n767), .A2(n51), .B1(n788), .B2(PCER_q[7]), .ZN(n504) );
  OAI211_X1 U701 ( .C1(n1461), .C2(n506), .A(n505), .B(n504), .ZN(n517) );
  AOI22_X1 U702 ( .A1(n691), .A2(mscratch_q[7]), .B1(n766), .B2(hwlp_end_i[39]), .ZN(n510) );
  AOI22_X1 U703 ( .A1(n136), .A2(hwlp_start_i[7]), .B1(n715), .B2(depc_o[7]), 
        .ZN(n509) );
  AOI22_X1 U704 ( .A1(n65), .A2(mepc_o[7]), .B1(n545), .B2(hwlp_cnt_i[7]), 
        .ZN(n508) );
  AOI22_X1 U705 ( .A1(n735), .A2(dcsr_q_cause__7_), .B1(n695), .B2(
        dscratch0_q[7]), .ZN(n507) );
  NAND4_X1 U706 ( .A1(n510), .A2(n509), .A3(n508), .A4(n507), .ZN(n516) );
  AOI22_X1 U707 ( .A1(n799), .A2(hwlp_start_i[39]), .B1(n761), .B2(
        cluster_id_i[2]), .ZN(n514) );
  AOI22_X1 U708 ( .A1(n782), .A2(hwlp_end_i[7]), .B1(n279), .B2(dscratch1_q[7]), .ZN(n513) );
  AOI22_X1 U709 ( .A1(n642), .A2(n15), .B1(n641), .B2(hwlp_cnt_i[39]), .ZN(
        n512) );
  AOI22_X1 U710 ( .A1(n800), .A2(n39), .B1(n748), .B2(n27), .ZN(n511) );
  NAND4_X1 U711 ( .A1(n514), .A2(n513), .A3(n512), .A4(n511), .ZN(n515) );
  OR3_X1 U712 ( .A1(n517), .A2(n516), .A3(n515), .ZN(csr_rdata_o[7]) );
  NAND2_X1 U713 ( .A1(csr_op_i[1]), .A2(csr_rdata_o[7]), .ZN(n519) );
  NAND2_X1 U714 ( .A1(csr_wdata_i[7]), .A2(n1362), .ZN(n518) );
  OAI21_X1 U715 ( .B1(n519), .B2(csr_wdata_i[7]), .A(n518), .ZN(n520) );
  INV_X1 U716 ( .A(n520), .ZN(n1393) );
  AOI22_X1 U733 ( .A1(n767), .A2(n48), .B1(n1380), .B2(utvec_o[7]), .ZN(n540)
         );
  AOI22_X1 U734 ( .A1(n800), .A2(n36), .B1(n748), .B2(n24), .ZN(n539) );
  AOI22_X1 U735 ( .A1(n790), .A2(PCCR_q[15]), .B1(n783), .B2(dscratch1_q[15]), 
        .ZN(n532) );
  AOI22_X1 U736 ( .A1(n695), .A2(dscratch0_q[15]), .B1(n690), .B2(
        hwlp_cnt_i[47]), .ZN(n531) );
  AOI22_X1 U737 ( .A1(n716), .A2(hwlp_end_i[15]), .B1(n801), .B2(uepc_o[15]), 
        .ZN(n530) );
  AOI22_X1 U738 ( .A1(n691), .A2(mscratch_q[15]), .B1(n136), .B2(
        hwlp_start_i[15]), .ZN(n529) );
  AND4_X1 U739 ( .A1(n532), .A2(n531), .A3(n530), .A4(n529), .ZN(n538) );
  AOI22_X1 U740 ( .A1(n137), .A2(hwlp_start_i[47]), .B1(n798), .B2(
        hwlp_end_i[47]), .ZN(n536) );
  AOI22_X1 U741 ( .A1(n609), .A2(debug_ebreakm_o), .B1(n760), .B2(
        hwlp_cnt_i[15]), .ZN(n535) );
  AOI22_X1 U742 ( .A1(n65), .A2(mepc_o[15]), .B1(n715), .B2(depc_o[15]), .ZN(
        n534) );
  AOI22_X1 U743 ( .A1(n642), .A2(n12), .B1(n734), .B2(mtvec_o[7]), .ZN(n533)
         );
  AND4_X1 U744 ( .A1(n536), .A2(n535), .A3(n534), .A4(n533), .ZN(n537) );
  NAND4_X1 U745 ( .A1(n540), .A2(n539), .A3(n538), .A4(n537), .ZN(
        csr_rdata_o[15]) );
  NAND2_X1 U746 ( .A1(n814), .A2(csr_rdata_o[15]), .ZN(n542) );
  NAND2_X1 U747 ( .A1(csr_wdata_i[15]), .A2(n1362), .ZN(n541) );
  OAI21_X1 U748 ( .B1(n542), .B2(csr_wdata_i[15]), .A(n541), .ZN(n543) );
  INV_X1 U749 ( .A(n543), .ZN(n1408) );
  AOI22_X1 U752 ( .A1(n782), .A2(hwlp_end_i[2]), .B1(n545), .B2(hwlp_cnt_i[2]), 
        .ZN(n561) );
  AOI22_X1 U753 ( .A1(n735), .A2(debug_single_step_o), .B1(n789), .B2(
        ucause_q[2]), .ZN(n560) );
  AOI22_X1 U754 ( .A1(n748), .A2(pmp_cfg_o[66]), .B1(n788), .B2(PCER_q[2]), 
        .ZN(n546) );
  OAI211_X1 U755 ( .C1(n1240), .C2(n1452), .A(n546), .B(n643), .ZN(n547) );
  AOI21_X1 U756 ( .B1(n800), .B2(pmp_cfg_o[34]), .A(n547), .ZN(n559) );
  AOI22_X1 U757 ( .A1(n696), .A2(hwlp_start_i[2]), .B1(n690), .B2(
        hwlp_cnt_i[34]), .ZN(n550) );
  AOI22_X1 U758 ( .A1(n695), .A2(dscratch0_q[2]), .B1(n548), .B2(uepc_o[2]), 
        .ZN(n549) );
  OAI211_X1 U759 ( .C1(n551), .C2(n1470), .A(n550), .B(n549), .ZN(n557) );
  AOI22_X1 U760 ( .A1(n65), .A2(mepc_o[2]), .B1(n799), .B2(hwlp_start_i[34]), 
        .ZN(n555) );
  AOI22_X1 U761 ( .A1(n153), .A2(mscratch_q[2]), .B1(n279), .B2(dscratch1_q[2]), .ZN(n554) );
  AOI22_X1 U762 ( .A1(n766), .A2(hwlp_end_i[34]), .B1(n701), .B2(depc_o[2]), 
        .ZN(n553) );
  AOI22_X1 U763 ( .A1(n1029), .A2(mcause_q[2]), .B1(n761), .B2(core_id_i[2]), 
        .ZN(n552) );
  NAND4_X1 U764 ( .A1(n555), .A2(n554), .A3(n553), .A4(n552), .ZN(n556) );
  AOI211_X1 U765 ( .C1(n642), .C2(pmp_cfg_o[98]), .A(n557), .B(n556), .ZN(n558) );
  NAND4_X1 U766 ( .A1(n561), .A2(n560), .A3(n559), .A4(n558), .ZN(
        csr_rdata_o[2]) );
  NAND2_X1 U767 ( .A1(csr_op_i[1]), .A2(csr_rdata_o[2]), .ZN(n563) );
  NAND2_X1 U768 ( .A1(csr_wdata_i[2]), .A2(n1362), .ZN(n562) );
  OAI21_X1 U769 ( .B1(n563), .B2(csr_wdata_i[2]), .A(n562), .ZN(n564) );
  INV_X1 U770 ( .A(n564), .ZN(n1442) );
  AOI22_X1 U787 ( .A1(n691), .A2(mscratch_q[17]), .B1(n760), .B2(
        hwlp_cnt_i[17]), .ZN(n576) );
  AOI22_X1 U788 ( .A1(n716), .A2(hwlp_end_i[17]), .B1(n801), .B2(uepc_o[17]), 
        .ZN(n575) );
  AOI22_X1 U789 ( .A1(n690), .A2(hwlp_cnt_i[49]), .B1(n798), .B2(
        hwlp_end_i[49]), .ZN(n574) );
  AOI22_X1 U790 ( .A1(n783), .A2(dscratch1_q[17]), .B1(n410), .B2(
        dscratch0_q[17]), .ZN(n573) );
  NAND4_X1 U791 ( .A1(n576), .A2(n575), .A3(n574), .A4(n573), .ZN(n581) );
  AOI22_X1 U792 ( .A1(n179), .A2(pmp_cfg_o[81]), .B1(n767), .B2(pmp_cfg_o[17]), 
        .ZN(n579) );
  AOI22_X1 U793 ( .A1(n790), .A2(PCCR_q[17]), .B1(n735), .B2(dcsr_q_zero2__17_), .ZN(n578) );
  AOI22_X1 U794 ( .A1(n137), .A2(hwlp_start_i[49]), .B1(n136), .B2(
        hwlp_start_i[17]), .ZN(n577) );
  NAND3_X1 U795 ( .A1(n579), .A2(n578), .A3(n577), .ZN(n580) );
  NOR2_X1 U796 ( .A1(n581), .A2(n580), .ZN(n589) );
  AOI22_X1 U797 ( .A1(n1380), .A2(utvec_o[9]), .B1(n734), .B2(mtvec_o[9]), 
        .ZN(n588) );
  AOI22_X1 U798 ( .A1(n582), .A2(mepc_o[17]), .B1(n701), .B2(depc_o[17]), .ZN(
        n587) );
  NAND2_X1 U799 ( .A1(mstatus_q[0]), .A2(n770), .ZN(n584) );
  NAND2_X1 U800 ( .A1(pmp_cfg_o[113]), .A2(n642), .ZN(n583) );
  NAND2_X1 U801 ( .A1(n584), .A2(n583), .ZN(n585) );
  AOI21_X1 U802 ( .B1(n800), .B2(pmp_cfg_o[49]), .A(n585), .ZN(n586) );
  NAND4_X1 U803 ( .A1(n589), .A2(n588), .A3(n587), .A4(n586), .ZN(
        csr_rdata_o[17]) );
  INV_X1 U804 ( .A(csr_wdata_i[17]), .ZN(n590) );
  NAND3_X1 U805 ( .A1(csr_rdata_o[17]), .A2(csr_op_i[1]), .A3(n590), .ZN(n592)
         );
  NAND2_X1 U806 ( .A1(csr_wdata_i[17]), .A2(n1362), .ZN(n591) );
  AND2_X1 U807 ( .A1(n592), .A2(n591), .ZN(n1410) );
  INV_X1 U811 ( .A(n1198), .ZN(n954) );
  NAND2_X1 U812 ( .A1(n743), .A2(n954), .ZN(n946) );
  INV_X1 U813 ( .A(n946), .ZN(n945) );
  AOI22_X1 U814 ( .A1(n946), .A2(mstatus_q[0]), .B1(hwlp_data_o[17]), .B2(n945), .ZN(n594) );
  INV_X1 U815 ( .A(n594), .ZN(N2756) );
  CLKBUF_X1 U818 ( .A(n1007), .Z(hwlp_data_o[22]) );
  AOI22_X1 U832 ( .A1(n734), .A2(mtvec_o[15]), .B1(n799), .B2(hwlp_start_i[55]), .ZN(n602) );
  OAI211_X1 U833 ( .C1(n1240), .C2(n1465), .A(n602), .B(n643), .ZN(n608) );
  AOI22_X1 U834 ( .A1(n695), .A2(dscratch0_q[23]), .B1(n701), .B2(depc_o[23]), 
        .ZN(n606) );
  AOI22_X1 U835 ( .A1(n716), .A2(hwlp_end_i[23]), .B1(n760), .B2(
        hwlp_cnt_i[23]), .ZN(n605) );
  AOI22_X1 U836 ( .A1(n691), .A2(mscratch_q[23]), .B1(n548), .B2(uepc_o[23]), 
        .ZN(n604) );
  AOI22_X1 U837 ( .A1(n65), .A2(mepc_o[23]), .B1(n696), .B2(hwlp_start_i[23]), 
        .ZN(n603) );
  NAND4_X1 U838 ( .A1(n606), .A2(n605), .A3(n604), .A4(n603), .ZN(n607) );
  AOI211_X1 U839 ( .C1(n1380), .C2(utvec_o[15]), .A(n608), .B(n607), .ZN(n615)
         );
  AOI22_X1 U840 ( .A1(n609), .A2(dcsr_q_zero2__23_), .B1(n279), .B2(
        dscratch1_q[23]), .ZN(n613) );
  AOI22_X1 U841 ( .A1(n690), .A2(hwlp_cnt_i[55]), .B1(n766), .B2(
        hwlp_end_i[55]), .ZN(n612) );
  AOI22_X1 U842 ( .A1(n642), .A2(n9), .B1(n800), .B2(n33), .ZN(n611) );
  AOI22_X1 U843 ( .A1(n767), .A2(n45), .B1(n748), .B2(n21), .ZN(n610) );
  AND4_X1 U844 ( .A1(n613), .A2(n612), .A3(n611), .A4(n610), .ZN(n614) );
  NAND2_X1 U845 ( .A1(n615), .A2(n614), .ZN(csr_rdata_o[23]) );
  NAND2_X1 U846 ( .A1(n814), .A2(csr_rdata_o[23]), .ZN(n617) );
  NAND2_X1 U847 ( .A1(csr_wdata_i[23]), .A2(n1362), .ZN(n616) );
  OAI21_X2 U848 ( .B1(n617), .B2(csr_wdata_i[23]), .A(n616), .ZN(
        hwlp_data_o[23]) );
  AOI22_X1 U859 ( .A1(n783), .A2(dscratch1_q[29]), .B1(n696), .B2(
        hwlp_start_i[29]), .ZN(n634) );
  AOI22_X1 U860 ( .A1(n799), .A2(hwlp_start_i[61]), .B1(n695), .B2(
        dscratch0_q[29]), .ZN(n633) );
  AOI22_X1 U861 ( .A1(n790), .A2(PCCR_q[29]), .B1(n798), .B2(hwlp_end_i[61]), 
        .ZN(n625) );
  AOI22_X1 U862 ( .A1(n65), .A2(mepc_o[29]), .B1(n545), .B2(hwlp_cnt_i[29]), 
        .ZN(n624) );
  AOI22_X1 U863 ( .A1(n716), .A2(hwlp_end_i[29]), .B1(n548), .B2(uepc_o[29]), 
        .ZN(n623) );
  NAND3_X1 U864 ( .A1(n625), .A2(n624), .A3(n623), .ZN(n631) );
  AOI22_X1 U865 ( .A1(n691), .A2(mscratch_q[29]), .B1(n690), .B2(
        hwlp_cnt_i[61]), .ZN(n629) );
  AOI22_X1 U866 ( .A1(n748), .A2(n20), .B1(n701), .B2(depc_o[29]), .ZN(n628)
         );
  AOI22_X1 U867 ( .A1(n642), .A2(n8), .B1(n734), .B2(mtvec_o[21]), .ZN(n627)
         );
  AOI22_X1 U868 ( .A1(n767), .A2(n44), .B1(n1380), .B2(utvec_o[21]), .ZN(n626)
         );
  NAND4_X1 U869 ( .A1(n629), .A2(n628), .A3(n627), .A4(n626), .ZN(n630) );
  AOI211_X1 U870 ( .C1(n180), .C2(n32), .A(n631), .B(n630), .ZN(n632) );
  NAND3_X1 U871 ( .A1(n634), .A2(n633), .A3(n632), .ZN(csr_rdata_o[29]) );
  NAND2_X1 U872 ( .A1(n814), .A2(csr_rdata_o[29]), .ZN(n636) );
  NAND2_X1 U873 ( .A1(csr_wdata_i[29]), .A2(n1362), .ZN(n635) );
  INV_X1 U874 ( .A(n929), .ZN(n1423) );
  AOI22_X1 U884 ( .A1(n695), .A2(dscratch0_q[30]), .B1(n701), .B2(depc_o[30]), 
        .ZN(n657) );
  AOI22_X1 U885 ( .A1(n696), .A2(hwlp_start_i[30]), .B1(n641), .B2(
        hwlp_cnt_i[62]), .ZN(n656) );
  AOI22_X1 U886 ( .A1(n642), .A2(n7), .B1(n782), .B2(hwlp_end_i[30]), .ZN(n644) );
  OAI211_X1 U887 ( .C1(n1240), .C2(n1466), .A(n644), .B(n643), .ZN(n645) );
  AOI21_X1 U888 ( .B1(n179), .B2(n19), .A(n645), .ZN(n655) );
  AOI22_X1 U889 ( .A1(n767), .A2(n43), .B1(n734), .B2(mtvec_o[22]), .ZN(n646)
         );
  OAI21_X1 U890 ( .B1(n647), .B2(n1467), .A(n646), .ZN(n653) );
  AOI22_X1 U891 ( .A1(n783), .A2(dscratch1_q[30]), .B1(n801), .B2(uepc_o[30]), 
        .ZN(n651) );
  AOI22_X1 U892 ( .A1(n735), .A2(dcsr_q_xdebugver__30_), .B1(n65), .B2(
        mepc_o[30]), .ZN(n650) );
  AOI22_X1 U893 ( .A1(n137), .A2(hwlp_start_i[62]), .B1(n766), .B2(
        hwlp_end_i[62]), .ZN(n649) );
  AOI22_X1 U894 ( .A1(n691), .A2(mscratch_q[30]), .B1(n545), .B2(
        hwlp_cnt_i[30]), .ZN(n648) );
  NAND4_X1 U895 ( .A1(n651), .A2(n650), .A3(n649), .A4(n648), .ZN(n652) );
  AOI211_X1 U896 ( .C1(n180), .C2(n31), .A(n653), .B(n652), .ZN(n654) );
  NAND4_X1 U897 ( .A1(n657), .A2(n656), .A3(n655), .A4(n654), .ZN(
        csr_rdata_o[30]) );
  NAND2_X1 U898 ( .A1(n814), .A2(csr_rdata_o[30]), .ZN(n659) );
  NAND2_X1 U899 ( .A1(csr_wdata_i[30]), .A2(n1362), .ZN(n658) );
  INV_X1 U900 ( .A(n931), .ZN(n1426) );
  AOI22_X1 U918 ( .A1(n790), .A2(PCCR_q[1]), .B1(n641), .B2(hwlp_cnt_i[33]), 
        .ZN(n671) );
  AOI22_X1 U919 ( .A1(n766), .A2(hwlp_end_i[33]), .B1(n701), .B2(depc_o[1]), 
        .ZN(n670) );
  AOI22_X1 U920 ( .A1(n153), .A2(mscratch_q[1]), .B1(n801), .B2(uepc_o[1]), 
        .ZN(n669) );
  AOI22_X1 U921 ( .A1(n137), .A2(hwlp_start_i[33]), .B1(n136), .B2(
        hwlp_start_i[1]), .ZN(n668) );
  NAND4_X1 U922 ( .A1(n671), .A2(n670), .A3(n669), .A4(n668), .ZN(n687) );
  AOI22_X1 U923 ( .A1(n1029), .A2(mcause_q[1]), .B1(n761), .B2(core_id_i[1]), 
        .ZN(n677) );
  AOI22_X1 U924 ( .A1(n782), .A2(hwlp_end_i[1]), .B1(n65), .B2(mepc_o[1]), 
        .ZN(n676) );
  AOI22_X1 U925 ( .A1(n783), .A2(dscratch1_q[1]), .B1(n545), .B2(hwlp_cnt_i[1]), .ZN(n675) );
  NOR3_X1 U926 ( .A1(n881), .A2(n673), .A3(n672), .ZN(n747) );
  AOI22_X1 U927 ( .A1(n789), .A2(ucause_q[1]), .B1(priv_lvl_o[1]), .B2(n747), 
        .ZN(n674) );
  NAND4_X1 U928 ( .A1(n677), .A2(n676), .A3(n675), .A4(n674), .ZN(n686) );
  NOR2_X1 U929 ( .A1(n679), .A2(n678), .ZN(n730) );
  INV_X1 U930 ( .A(n730), .ZN(n1235) );
  INV_X1 U931 ( .A(n788), .ZN(n857) );
  AOI22_X1 U932 ( .A1(n735), .A2(dcsr_q_prv__1_), .B1(n410), .B2(
        dscratch0_q[1]), .ZN(n681) );
  AOI22_X1 U933 ( .A1(n748), .A2(pmp_cfg_o[65]), .B1(n800), .B2(pmp_cfg_o[33]), 
        .ZN(n680) );
  OAI211_X1 U934 ( .C1(n857), .C2(n1458), .A(n681), .B(n680), .ZN(n682) );
  INV_X1 U935 ( .A(n682), .ZN(n684) );
  AOI22_X1 U936 ( .A1(n181), .A2(pmp_cfg_o[97]), .B1(n767), .B2(pmp_cfg_o[1]), 
        .ZN(n683) );
  OAI211_X1 U937 ( .C1(n1235), .C2(n1584), .A(n684), .B(n683), .ZN(n685) );
  OR3_X1 U938 ( .A1(n687), .A2(n686), .A3(n685), .ZN(csr_rdata_o[1]) );
  AOI21_X1 U939 ( .B1(csr_op_i[1]), .B2(csr_rdata_o[1]), .A(csr_wdata_i[1]), 
        .ZN(n688) );
  AOI21_X1 U940 ( .B1(csr_wdata_i[1]), .B2(n1257), .A(n688), .ZN(n1031) );
  AOI22_X1 U944 ( .A1(n790), .A2(PCCR_q[28]), .B1(n799), .B2(hwlp_start_i[60]), 
        .ZN(n694) );
  AOI22_X1 U945 ( .A1(n766), .A2(hwlp_end_i[60]), .B1(n760), .B2(
        hwlp_cnt_i[28]), .ZN(n693) );
  AOI22_X1 U946 ( .A1(n691), .A2(mscratch_q[28]), .B1(n690), .B2(
        hwlp_cnt_i[60]), .ZN(n692) );
  AND3_X1 U947 ( .A1(n694), .A2(n693), .A3(n692), .ZN(n707) );
  AOI22_X1 U948 ( .A1(n695), .A2(dscratch0_q[28]), .B1(n801), .B2(uepc_o[28]), 
        .ZN(n700) );
  AOI22_X1 U949 ( .A1(n65), .A2(mepc_o[28]), .B1(n696), .B2(hwlp_start_i[28]), 
        .ZN(n699) );
  AOI22_X1 U950 ( .A1(n748), .A2(pmp_cfg_o[92]), .B1(n1380), .B2(utvec_o[20]), 
        .ZN(n698) );
  AOI22_X1 U951 ( .A1(n181), .A2(pmp_cfg_o[124]), .B1(n180), .B2(pmp_cfg_o[60]), .ZN(n697) );
  AND4_X1 U952 ( .A1(n700), .A2(n699), .A3(n698), .A4(n697), .ZN(n706) );
  AOI22_X1 U953 ( .A1(n734), .A2(mtvec_o[20]), .B1(n279), .B2(dscratch1_q[28]), 
        .ZN(n705) );
  AOI22_X1 U954 ( .A1(n782), .A2(hwlp_end_i[28]), .B1(n701), .B2(depc_o[28]), 
        .ZN(n703) );
  NAND2_X1 U955 ( .A1(n767), .A2(pmp_cfg_o[28]), .ZN(n702) );
  AND2_X1 U956 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND4_X1 U957 ( .A1(n707), .A2(n706), .A3(n705), .A4(n704), .ZN(
        csr_rdata_o[28]) );
  NOR2_X1 U958 ( .A1(n708), .A2(csr_wdata_i[28]), .ZN(n709) );
  NAND2_X1 U959 ( .A1(csr_rdata_o[28]), .A2(n709), .ZN(n711) );
  NAND2_X1 U960 ( .A1(csr_wdata_i[28]), .A2(n1362), .ZN(n710) );
  NAND2_X1 U961 ( .A1(n711), .A2(n710), .ZN(hwlp_data_o[28]) );
  AOI22_X1 U962 ( .A1(n180), .A2(pmp_cfg_o[41]), .B1(pmp_cfg_o[105]), .B2(n181), .ZN(n713) );
  AOI22_X1 U963 ( .A1(n790), .A2(PCCR_q[9]), .B1(n695), .B2(dscratch0_q[9]), 
        .ZN(n712) );
  OAI211_X1 U964 ( .C1(n714), .C2(n1553), .A(n713), .B(n712), .ZN(n727) );
  AOI22_X1 U965 ( .A1(n783), .A2(dscratch1_q[9]), .B1(n715), .B2(depc_o[9]), 
        .ZN(n720) );
  AOI22_X1 U966 ( .A1(n761), .A2(cluster_id_i[4]), .B1(n760), .B2(
        hwlp_cnt_i[9]), .ZN(n719) );
  AOI22_X1 U967 ( .A1(n716), .A2(hwlp_end_i[9]), .B1(n690), .B2(hwlp_cnt_i[41]), .ZN(n718) );
  AOI22_X1 U968 ( .A1(n799), .A2(hwlp_start_i[41]), .B1(n801), .B2(uepc_o[9]), 
        .ZN(n717) );
  NAND4_X1 U969 ( .A1(n720), .A2(n719), .A3(n718), .A4(n717), .ZN(n726) );
  AOI22_X1 U970 ( .A1(n1380), .A2(utvec_o[1]), .B1(n788), .B2(PCER_q[9]), .ZN(
        n724) );
  AOI22_X1 U971 ( .A1(n153), .A2(mscratch_q[9]), .B1(n696), .B2(
        hwlp_start_i[9]), .ZN(n723) );
  AOI22_X1 U972 ( .A1(n65), .A2(mepc_o[9]), .B1(n798), .B2(hwlp_end_i[41]), 
        .ZN(n722) );
  AOI22_X1 U973 ( .A1(n767), .A2(pmp_cfg_o[9]), .B1(n748), .B2(pmp_cfg_o[73]), 
        .ZN(n721) );
  NAND4_X1 U974 ( .A1(n724), .A2(n723), .A3(n722), .A4(n721), .ZN(n725) );
  OR3_X1 U975 ( .A1(n727), .A2(n726), .A3(n725), .ZN(csr_rdata_o[9]) );
  NAND2_X1 U976 ( .A1(csr_op_i[1]), .A2(csr_rdata_o[9]), .ZN(n729) );
  NAND2_X1 U977 ( .A1(csr_wdata_i[9]), .A2(n1362), .ZN(n728) );
  OAI21_X2 U978 ( .B1(n729), .B2(csr_wdata_i[9]), .A(n728), .ZN(hwlp_data_o[9]) );
  AOI22_X1 U979 ( .A1(n789), .A2(ucause_q[0]), .B1(n801), .B2(n4), .ZN(n733)
         );
  AOI22_X1 U980 ( .A1(n761), .A2(core_id_i[0]), .B1(n760), .B2(hwlp_cnt_i[0]), 
        .ZN(n732) );
  AOI22_X1 U981 ( .A1(n788), .A2(PCER_q[0]), .B1(n730), .B2(PCMR_q[0]), .ZN(
        n731) );
  NAND3_X1 U982 ( .A1(n733), .A2(n732), .A3(n731), .ZN(n756) );
  AOI21_X1 U983 ( .B1(n782), .B2(hwlp_end_i[0]), .A(n734), .ZN(n738) );
  AOI22_X1 U984 ( .A1(dcsr_q_prv__0_), .A2(n735), .B1(n153), .B2(mscratch_q[0]), .ZN(n737) );
  AOI22_X1 U985 ( .A1(n65), .A2(n3), .B1(n279), .B2(dscratch1_q[0]), .ZN(n736)
         );
  NAND3_X1 U986 ( .A1(n738), .A2(n737), .A3(n736), .ZN(n739) );
  AOI211_X1 U987 ( .C1(n790), .C2(PCCR_q[0]), .A(n1380), .B(n739), .ZN(n740)
         );
  INV_X1 U988 ( .A(n740), .ZN(n755) );
  NOR2_X1 U989 ( .A1(n741), .A2(n881), .ZN(n742) );
  NOR2_X1 U990 ( .A1(csr_addr_i[11]), .A2(n826), .ZN(n791) );
  AOI22_X1 U991 ( .A1(mstatus_q[6]), .A2(n791), .B1(n767), .B2(pmp_cfg_o[0]), 
        .ZN(n746) );
  AOI22_X1 U992 ( .A1(n136), .A2(hwlp_start_i[0]), .B1(n641), .B2(
        hwlp_cnt_i[32]), .ZN(n745) );
  AOI22_X1 U993 ( .A1(n137), .A2(hwlp_start_i[32]), .B1(n410), .B2(
        dscratch0_q[0]), .ZN(n744) );
  NAND3_X1 U994 ( .A1(n746), .A2(n745), .A3(n744), .ZN(n754) );
  AOI22_X1 U995 ( .A1(n766), .A2(hwlp_end_i[32]), .B1(n715), .B2(n5), .ZN(n752) );
  AOI22_X1 U996 ( .A1(n180), .A2(pmp_cfg_o[32]), .B1(\priv_lvl_o[0] ), .B2(
        n747), .ZN(n751) );
  AOI22_X1 U997 ( .A1(n642), .A2(pmp_cfg_o[96]), .B1(n748), .B2(pmp_cfg_o[64]), 
        .ZN(n750) );
  NAND2_X1 U998 ( .A1(n1029), .A2(mcause_q[0]), .ZN(n749) );
  NAND4_X1 U999 ( .A1(n752), .A2(n751), .A3(n750), .A4(n749), .ZN(n753) );
  OR4_X1 U1000 ( .A1(n756), .A2(n755), .A3(n754), .A4(n753), .ZN(
        csr_rdata_o[0]) );
  INV_X1 U1001 ( .A(csr_wdata_i[0]), .ZN(n757) );
  NAND3_X1 U1002 ( .A1(csr_rdata_o[0]), .A2(csr_op_i[1]), .A3(n757), .ZN(n759)
         );
  AND2_X1 U1003 ( .A1(n759), .A2(n758), .ZN(n1387) );
  AOI22_X1 U1005 ( .A1(n783), .A2(dscratch1_q[3]), .B1(n760), .B2(
        hwlp_cnt_i[3]), .ZN(n765) );
  AOI22_X1 U1006 ( .A1(n136), .A2(hwlp_start_i[3]), .B1(n641), .B2(
        hwlp_cnt_i[35]), .ZN(n764) );
  AOI22_X1 U1007 ( .A1(n153), .A2(mscratch_q[3]), .B1(n789), .B2(ucause_q[3]), 
        .ZN(n763) );
  AOI22_X1 U1008 ( .A1(n1029), .A2(mcause_q[3]), .B1(n761), .B2(core_id_i[3]), 
        .ZN(n762) );
  NAND4_X1 U1009 ( .A1(n765), .A2(n764), .A3(n763), .A4(n762), .ZN(n781) );
  AOI22_X1 U1010 ( .A1(n766), .A2(hwlp_end_i[35]), .B1(n801), .B2(uepc_o[3]), 
        .ZN(n774) );
  AOI22_X1 U1011 ( .A1(n782), .A2(hwlp_end_i[3]), .B1(n410), .B2(
        dscratch0_q[3]), .ZN(n769) );
  NAND2_X1 U1012 ( .A1(n767), .A2(pmp_cfg_o[3]), .ZN(n768) );
  AND2_X1 U1013 ( .A1(n769), .A2(n768), .ZN(n773) );
  AOI22_X1 U1014 ( .A1(n179), .A2(pmp_cfg_o[67]), .B1(mstatus_q[5]), .B2(n770), 
        .ZN(n772) );
  AOI22_X1 U1015 ( .A1(pmp_cfg_o[99]), .A2(n181), .B1(n180), .B2(pmp_cfg_o[35]), .ZN(n771) );
  NAND4_X1 U1016 ( .A1(n774), .A2(n773), .A3(n772), .A4(n771), .ZN(n779) );
  NAND2_X1 U1017 ( .A1(n788), .A2(PCER_q[3]), .ZN(n777) );
  AOI22_X1 U1018 ( .A1(n790), .A2(PCCR_q[3]), .B1(n715), .B2(depc_o[3]), .ZN(
        n776) );
  AOI22_X1 U1019 ( .A1(n65), .A2(mepc_o[3]), .B1(n799), .B2(hwlp_start_i[35]), 
        .ZN(n775) );
  NAND3_X1 U1020 ( .A1(n777), .A2(n776), .A3(n775), .ZN(n778) );
  OR2_X1 U1021 ( .A1(n779), .A2(n778), .ZN(n780) );
  OR2_X1 U1022 ( .A1(n781), .A2(n780), .ZN(csr_rdata_o[3]) );
  AOI22_X1 U1023 ( .A1(n696), .A2(hwlp_start_i[4]), .B1(n690), .B2(
        hwlp_cnt_i[36]), .ZN(n787) );
  AOI22_X1 U1024 ( .A1(n153), .A2(mscratch_q[4]), .B1(n65), .B2(mepc_o[4]), 
        .ZN(n786) );
  AOI22_X1 U1025 ( .A1(n782), .A2(hwlp_end_i[4]), .B1(n701), .B2(depc_o[4]), 
        .ZN(n785) );
  AOI22_X1 U1026 ( .A1(n783), .A2(dscratch1_q[4]), .B1(n545), .B2(
        hwlp_cnt_i[4]), .ZN(n784) );
  NAND4_X1 U1027 ( .A1(n787), .A2(n786), .A3(n785), .A4(n784), .ZN(n797) );
  NAND2_X1 U1028 ( .A1(n788), .A2(PCER_q[4]), .ZN(n795) );
  AOI22_X1 U1029 ( .A1(n790), .A2(PCCR_q[4]), .B1(n789), .B2(ucause_q[4]), 
        .ZN(n794) );
  NAND2_X1 U1030 ( .A1(n791), .A2(mstatus_q[4]), .ZN(n793) );
  NAND2_X1 U1031 ( .A1(n695), .A2(dscratch0_q[4]), .ZN(n792) );
  NAND4_X1 U1032 ( .A1(n795), .A2(n794), .A3(n793), .A4(n792), .ZN(n796) );
  NOR2_X1 U1033 ( .A1(n797), .A2(n796), .ZN(n807) );
  AOI22_X1 U1034 ( .A1(n799), .A2(hwlp_start_i[36]), .B1(n798), .B2(
        hwlp_end_i[36]), .ZN(n806) );
  AOI22_X1 U1035 ( .A1(n748), .A2(pmp_cfg_o[68]), .B1(n800), .B2(pmp_cfg_o[36]), .ZN(n805) );
  AOI22_X1 U1036 ( .A1(n1029), .A2(mcause_q[4]), .B1(n801), .B2(uepc_o[4]), 
        .ZN(n803) );
  AOI22_X1 U1037 ( .A1(n181), .A2(pmp_cfg_o[100]), .B1(n767), .B2(pmp_cfg_o[4]), .ZN(n802) );
  AND2_X1 U1038 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND4_X1 U1039 ( .A1(n807), .A2(n806), .A3(n805), .A4(n804), .ZN(
        csr_rdata_o[4]) );
  INV_X1 U1040 ( .A(csr_wdata_i[4]), .ZN(n808) );
  NAND3_X1 U1041 ( .A1(csr_rdata_o[4]), .A2(csr_op_i[1]), .A3(n808), .ZN(n810)
         );
  NAND2_X1 U1042 ( .A1(csr_wdata_i[4]), .A2(n1362), .ZN(n809) );
  AND2_X1 U1043 ( .A1(n810), .A2(n809), .ZN(n1390) );
  NAND4_X1 U1045 ( .A1(n813), .A2(n812), .A3(n954), .A4(n811), .ZN(n1225) );
  NOR3_X1 U1046 ( .A1(n1371), .A2(n1372), .A3(n1225), .ZN(hwlp_regid_o[0]) );
  INV_X1 U1048 ( .A(csr_rdata_o[3]), .ZN(n818) );
  INV_X1 U1049 ( .A(csr_wdata_i[3]), .ZN(n815) );
  NAND2_X1 U1050 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U1051 ( .A1(csr_wdata_i[3]), .A2(n1362), .ZN(n816) );
  OAI21_X1 U1052 ( .B1(n818), .B2(n817), .A(n816), .ZN(n4184) );
  INV_X1 U1055 ( .A(csr_op_i[0]), .ZN(n855) );
  NOR2_X2 U1056 ( .A1(n855), .A2(n857), .ZN(n1233) );
  NOR2_X1 U1057 ( .A1(n1394), .A2(n857), .ZN(n1231) );
  OAI211_X1 U1058 ( .C1(n1362), .C2(n1479), .A(n1231), .B(csr_wdata_i[11]), 
        .ZN(n819) );
  OAI21_X1 U1059 ( .B1(n1233), .B2(n1479), .A(n819), .ZN(PCER_n[11]) );
  MUX2_X1 U1060 ( .A(hwlp_data_o[11]), .B(pmp_cfg_o[107]), .S(n1446), .Z(n2041) );
  MUX2_X1 U1061 ( .A(hwlp_data_o[11]), .B(pmp_cfg_o[43]), .S(n864), .Z(n2105)
         );
  NAND2_X1 U1063 ( .A1(debug_csr_save_i), .A2(n942), .ZN(n1221) );
  AOI21_X1 U1066 ( .B1(csr_restore_dret_i), .B2(dcsr_q_prv__1_), .A(n821), 
        .ZN(n822) );
  AOI21_X1 U1067 ( .B1(n1459), .B2(n823), .A(n822), .ZN(n2022) );
  MUX2_X1 U1070 ( .A(hwlp_data_o[12]), .B(pmp_cfg_o[12]), .S(n1443), .Z(n2138)
         );
  OAI211_X1 U1079 ( .C1(n1362), .C2(n1457), .A(csr_wdata_i[4]), .B(n1231), 
        .ZN(n825) );
  OAI21_X1 U1080 ( .B1(n1233), .B2(n1457), .A(n825), .ZN(PCER_n[4]) );
  MUX2_X1 U1082 ( .A(hwlp_data_o[4]), .B(pmp_cfg_o[36]), .S(n864), .Z(n2114)
         );
  MUX2_X1 U1083 ( .A(hwlp_data_o[4]), .B(pmp_cfg_o[68]), .S(n865), .Z(n2082)
         );
  NOR2_X1 U1084 ( .A1(n826), .A2(n1198), .ZN(n833) );
  INV_X1 U1085 ( .A(n833), .ZN(n832) );
  AOI22_X1 U1086 ( .A1(hwlp_data_o[4]), .A2(n833), .B1(n832), .B2(mstatus_q[4]), .ZN(n828) );
  NAND2_X1 U1087 ( .A1(n850), .A2(n1047), .ZN(n831) );
  INV_X1 U1088 ( .A(n1212), .ZN(n1209) );
  INV_X1 U1089 ( .A(csr_restore_uret_i), .ZN(n839) );
  NAND2_X1 U1090 ( .A1(n1209), .A2(mstatus_q[6]), .ZN(n827) );
  OAI211_X1 U1091 ( .C1(n828), .C2(n1209), .A(n839), .B(n827), .ZN(n2807) );
  AOI211_X1 U1092 ( .C1(csr_save_cause_i), .C2(n831), .A(n830), .B(n829), .ZN(
        n838) );
  AOI22_X1 U1093 ( .A1(hwlp_data_o[0]), .A2(n833), .B1(mstatus_q[6]), .B2(n832), .ZN(n837) );
  NAND3_X1 U1094 ( .A1(csr_restore_mret_i), .A2(mstatus_q[3]), .A3(n834), .ZN(
        n836) );
  NAND2_X1 U1095 ( .A1(csr_restore_uret_i), .A2(mstatus_q[4]), .ZN(n835) );
  OAI211_X1 U1096 ( .C1(n838), .C2(n837), .A(n836), .B(n835), .ZN(mstatus_n[4]) );
  OAI21_X1 U1101 ( .B1(csr_save_cause_i), .B2(n847), .A(n1122), .ZN(n840) );
  NAND2_X1 U1102 ( .A1(n840), .A2(n839), .ZN(n941) );
  NOR2_X1 U1104 ( .A1(n941), .A2(n3925), .ZN(n841) );
  NAND3_X1 U1105 ( .A1(n841), .A2(mstatus_q[2]), .A3(mstatus_q[1]), .ZN(n843)
         );
  NAND2_X1 U1106 ( .A1(n841), .A2(n847), .ZN(n848) );
  OAI22_X1 U1107 ( .A1(n1702), .A2(n946), .B1(n945), .B2(n1454), .ZN(n842) );
  NAND3_X1 U1108 ( .A1(n843), .A2(n848), .A3(n842), .ZN(n845) );
  NAND4_X1 U1109 ( .A1(csr_restore_mret_i), .A2(mstatus_q[2]), .A3(
        mstatus_q[1]), .A4(mstatus_q[3]), .ZN(n844) );
  NAND2_X1 U1110 ( .A1(n845), .A2(n844), .ZN(mstatus_n[3]) );
  NOR2_X1 U1111 ( .A1(n846), .A2(n1455), .ZN(u_irq_enable_o) );
  INV_X1 U1112 ( .A(debug_csr_save_i), .ZN(n951) );
  NAND2_X1 U1113 ( .A1(n942), .A2(n951), .ZN(n948) );
  OAI222_X1 U1114 ( .A1(n1461), .A2(n945), .B1(n946), .B2(n1393), .C1(n847), 
        .C2(n943), .ZN(n849) );
  NAND2_X1 U1115 ( .A1(n849), .A2(n848), .ZN(n853) );
  INV_X1 U1116 ( .A(n850), .ZN(n851) );
  NAND3_X1 U1117 ( .A1(csr_save_cause_i), .A2(u_irq_enable_o), .A3(n851), .ZN(
        n852) );
  OAI211_X1 U1118 ( .C1(n1454), .C2(n948), .A(n853), .B(n852), .ZN(
        mstatus_n[2]) );
  OAI211_X1 U1119 ( .C1(n1362), .C2(n1468), .A(n1385), .B(csr_wdata_i[0]), 
        .ZN(n854) );
  OAI22_X1 U1120 ( .A1(n1233), .A2(n1468), .B1(n857), .B2(n854), .ZN(PCER_n[0]) );
  NOR2_X1 U1121 ( .A1(n855), .A2(n1235), .ZN(n1236) );
  OAI211_X1 U1122 ( .C1(n1362), .C2(n1456), .A(n1385), .B(csr_wdata_i[0]), 
        .ZN(n856) );
  OAI22_X1 U1123 ( .A1(n1236), .A2(n1456), .B1(n1235), .B2(n856), .ZN(
        PCMR_n[0]) );
  OAI211_X1 U1125 ( .C1(n1362), .C2(n1458), .A(csr_wdata_i[1]), .B(n1385), 
        .ZN(n858) );
  OAI22_X1 U1126 ( .A1(n1233), .A2(n1458), .B1(n858), .B2(n857), .ZN(PCER_n[1]) );
  OAI211_X1 U1129 ( .C1(n1362), .C2(n1471), .A(n1231), .B(csr_wdata_i[5]), 
        .ZN(n859) );
  OAI21_X1 U1130 ( .B1(n1233), .B2(n1471), .A(n859), .ZN(PCER_n[5]) );
  OAI211_X1 U1131 ( .C1(n1362), .C2(n1472), .A(n1231), .B(csr_wdata_i[6]), 
        .ZN(n860) );
  OAI21_X1 U1132 ( .B1(n1233), .B2(n1472), .A(n860), .ZN(PCER_n[6]) );
  MUX2_X1 U1135 ( .A(hwlp_data_o[9]), .B(pmp_cfg_o[41]), .S(n864), .Z(n2103)
         );
  MUX2_X1 U1136 ( .A(hwlp_data_o[9]), .B(pmp_cfg_o[9]), .S(n1443), .Z(n2135)
         );
  MUX2_X1 U1137 ( .A(hwlp_data_o[9]), .B(pmp_cfg_o[73]), .S(n865), .Z(n2071)
         );
  OAI211_X1 U1138 ( .C1(n1362), .C2(n1480), .A(csr_wdata_i[10]), .B(n1231), 
        .ZN(n861) );
  OAI21_X1 U1139 ( .B1(n1233), .B2(n1480), .A(n861), .ZN(PCER_n[10]) );
  MUX2_X1 U1146 ( .A(hwlp_data_o[19]), .B(pmp_cfg_o[19]), .S(n1443), .Z(n2129)
         );
  MUX2_X1 U1147 ( .A(hwlp_data_o[19]), .B(pmp_cfg_o[115]), .S(n1446), .Z(n2033) );
  MUX2_X1 U1148 ( .A(hwlp_data_o[19]), .B(pmp_cfg_o[51]), .S(n864), .Z(n2097)
         );
  MUX2_X1 U1149 ( .A(hwlp_data_o[19]), .B(pmp_cfg_o[83]), .S(n865), .Z(n2065)
         );
  MUX2_X1 U1151 ( .A(hwlp_data_o[20]), .B(pmp_cfg_o[52]), .S(n864), .Z(n2098)
         );
  MUX2_X1 U1153 ( .A(hwlp_data_o[20]), .B(pmp_cfg_o[116]), .S(n1446), .Z(n2034) );
  MUX2_X1 U1154 ( .A(hwlp_data_o[24]), .B(pmp_cfg_o[24]), .S(n1443), .Z(n2126)
         );
  MUX2_X1 U1155 ( .A(hwlp_data_o[24]), .B(pmp_cfg_o[56]), .S(n864), .Z(n2094)
         );
  MUX2_X1 U1156 ( .A(hwlp_data_o[24]), .B(pmp_cfg_o[88]), .S(n865), .Z(n2062)
         );
  MUX2_X1 U1160 ( .A(hwlp_data_o[27]), .B(pmp_cfg_o[27]), .S(n1443), .Z(n2121)
         );
  MUX2_X1 U1161 ( .A(hwlp_data_o[27]), .B(pmp_cfg_o[123]), .S(n1446), .Z(n2025) );
  MUX2_X1 U1162 ( .A(hwlp_data_o[27]), .B(pmp_cfg_o[59]), .S(n864), .Z(n2089)
         );
  MUX2_X1 U1163 ( .A(hwlp_data_o[27]), .B(pmp_cfg_o[91]), .S(n865), .Z(n2057)
         );
  MUX2_X1 U1164 ( .A(hwlp_data_o[28]), .B(pmp_cfg_o[28]), .S(n1443), .Z(n2122)
         );
  MUX2_X1 U1165 ( .A(hwlp_data_o[28]), .B(pmp_cfg_o[124]), .S(n1446), .Z(n2026) );
  MUX2_X1 U1166 ( .A(hwlp_data_o[28]), .B(pmp_cfg_o[60]), .S(n864), .Z(n2090)
         );
  MUX2_X1 U1167 ( .A(hwlp_data_o[28]), .B(pmp_cfg_o[92]), .S(n865), .Z(n2058)
         );
  AND2_X1 U1168 ( .A1(PCER_q[10]), .A2(is_compressed_i), .ZN(n866) );
  OAI211_X1 U1169 ( .C1(PCER_q[1]), .C2(n866), .A(id_valid_i), .B(
        is_decoding_i_BAR), .ZN(n880) );
  NAND2_X1 U1170 ( .A1(jump_i), .A2(PCER_q[7]), .ZN(n871) );
  AOI21_X1 U1171 ( .B1(branch_taken_i), .B2(PCER_q[9]), .A(PCER_q[8]), .ZN(
        n867) );
  INV_X1 U1172 ( .A(n867), .ZN(n868) );
  AOI22_X1 U1173 ( .A1(jr_stall_i), .A2(PCER_q[3]), .B1(branch_i), .B2(n868), 
        .ZN(n870) );
  NAND2_X1 U1174 ( .A1(ld_stall_i), .A2(PCER_q[2]), .ZN(n869) );
  NAND3_X1 U1175 ( .A1(n871), .A2(n870), .A3(n869), .ZN(n878) );
  NOR2_X1 U1176 ( .A1(pc_set_i), .A2(n1457), .ZN(n872) );
  NAND2_X1 U1177 ( .A1(imiss_i), .A2(n872), .ZN(n876) );
  AOI21_X1 U1178 ( .B1(pipeline_stall_i), .B2(PCER_q[11]), .A(PCER_q[0]), .ZN(
        n875) );
  NAND2_X1 U1179 ( .A1(mem_load_i), .A2(PCER_q[5]), .ZN(n874) );
  NAND2_X1 U1180 ( .A1(mem_store_i), .A2(PCER_q[6]), .ZN(n873) );
  NAND4_X1 U1181 ( .A1(n876), .A2(n875), .A3(n874), .A4(n873), .ZN(n877) );
  AOI21_X1 U1182 ( .B1(id_valid_q), .B2(n878), .A(n877), .ZN(n879) );
  AOI21_X1 U1183 ( .B1(n880), .B2(n879), .A(n1456), .ZN(PCCR_inc_0_) );
  INV_X1 U1184 ( .A(n881), .ZN(n882) );
  INV_X1 U1288 ( .A(n893), .ZN(n894) );
  INV_X1 U1322 ( .A(n897), .ZN(n898) );
  INV_X1 U1356 ( .A(n901), .ZN(n902) );
  INV_X1 U1390 ( .A(n905), .ZN(n906) );
  AND2_X1 U1424 ( .A1(n1371), .A2(n909), .ZN(n910) );
  NOR2_X1 U1523 ( .A1(n1226), .A2(csr_addr_i[2]), .ZN(n919) );
  AND2_X1 U1557 ( .A1(n1371), .A2(n1372), .ZN(n922) );
  INV_X1 U1684 ( .A(n936), .ZN(n937) );
  NOR2_X1 U1719 ( .A1(n940), .A2(n1454), .ZN(m_irq_enable_o) );
  AOI22_X1 U1720 ( .A1(mstatus_q[1]), .A2(n946), .B1(n945), .B2(
        hwlp_data_o[11]), .ZN(n944) );
  AOI211_X1 U1721 ( .C1(csr_restore_mret_i), .C2(n943), .A(n942), .B(n941), 
        .ZN(n947) );
  AOI21_X1 U1722 ( .B1(n944), .B2(n948), .A(n947), .ZN(mstatus_n[0]) );
  AOI22_X1 U1723 ( .A1(mstatus_q[2]), .A2(n946), .B1(n945), .B2(
        hwlp_data_o[12]), .ZN(n949) );
  AOI21_X1 U1724 ( .B1(n949), .B2(n948), .A(n947), .ZN(mstatus_n[1]) );
  INV_X1 U1725 ( .A(n950), .ZN(n955) );
  NOR2_X1 U1727 ( .A1(csr_save_ex_i_BAR), .A2(n958), .ZN(n971) );
  INV_X1 U1728 ( .A(csr_save_if_i), .ZN(n952) );
  NOR2_X1 U1729 ( .A1(n952), .A2(csr_save_id_i), .ZN(n957) );
  INV_X1 U1730 ( .A(n957), .ZN(n953) );
  NAND2_X1 U1731 ( .A1(csr_save_ex_i_BAR), .A2(n953), .ZN(n1126) );
  NOR2_X1 U1732 ( .A1(n958), .A2(n1126), .ZN(n1012) );
  AOI22_X1 U1733 ( .A1(pc_ex_i[0]), .A2(n63), .B1(pc_id_i[0]), .B2(n62), .ZN(
        n960) );
  NAND2_X1 U1734 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1735 ( .A1(n957), .A2(csr_save_ex_i_BAR), .ZN(n1124) );
  NOR2_X1 U1736 ( .A1(n958), .A2(n1124), .ZN(n990) );
  AOI22_X1 U1737 ( .A1(n4), .A2(n67), .B1(pc_if_i[0]), .B2(n64), .ZN(n959) );
  OAI211_X1 U1738 ( .C1(n1387), .C2(n967), .A(n960), .B(n959), .ZN(uepc_n[0])
         );
  INV_X1 U1739 ( .A(n1031), .ZN(n1388) );
  AOI22_X1 U1743 ( .A1(n63), .A2(pc_ex_i[2]), .B1(n62), .B2(pc_id_i[2]), .ZN(
        n964) );
  AOI22_X1 U1746 ( .A1(n63), .A2(pc_ex_i[3]), .B1(n62), .B2(pc_id_i[3]), .ZN(
        n966) );
  AOI22_X1 U1749 ( .A1(n63), .A2(pc_ex_i[4]), .B1(n62), .B2(pc_id_i[4]), .ZN(
        n969) );
  AOI22_X1 U1750 ( .A1(uepc_o[4]), .A2(n67), .B1(n64), .B2(pc_if_i[4]), .ZN(
        n968) );
  OAI211_X1 U1751 ( .C1(n1390), .C2(n967), .A(n969), .B(n968), .ZN(uepc_n[4])
         );
  INV_X1 U1752 ( .A(n970), .ZN(n1391) );
  AOI22_X1 U1756 ( .A1(n63), .A2(pc_ex_i[6]), .B1(n62), .B2(pc_id_i[6]), .ZN(
        n975) );
  AOI22_X1 U1762 ( .A1(n64), .A2(pc_if_i[8]), .B1(n62), .B2(pc_id_i[8]), .ZN(
        n979) );
  INV_X1 U1765 ( .A(hwlp_data_o[9]), .ZN(n1447) );
  INV_X1 U1769 ( .A(hwlp_data_o[10]), .ZN(n1444) );
  AOI22_X1 U1770 ( .A1(n63), .A2(pc_ex_i[10]), .B1(n62), .B2(pc_id_i[10]), 
        .ZN(n983) );
  AOI22_X1 U1773 ( .A1(n63), .A2(pc_ex_i[11]), .B1(n62), .B2(pc_id_i[11]), 
        .ZN(n985) );
  AOI22_X1 U1774 ( .A1(uepc_o[11]), .A2(n67), .B1(n64), .B2(pc_if_i[11]), .ZN(
        n984) );
  OAI211_X1 U1775 ( .C1(n1404), .C2(n967), .A(n985), .B(n984), .ZN(uepc_n[11])
         );
  AOI22_X1 U1776 ( .A1(n990), .A2(pc_if_i[12]), .B1(n63), .B2(pc_ex_i[12]), 
        .ZN(n987) );
  AOI22_X1 U1777 ( .A1(uepc_o[12]), .A2(n67), .B1(n62), .B2(pc_id_i[12]), .ZN(
        n986) );
  OAI211_X1 U1778 ( .C1(n1405), .C2(n967), .A(n987), .B(n986), .ZN(uepc_n[12])
         );
  AOI22_X1 U1779 ( .A1(n63), .A2(pc_ex_i[13]), .B1(n62), .B2(pc_id_i[13]), 
        .ZN(n989) );
  AOI22_X1 U1788 ( .A1(n64), .A2(pc_if_i[16]), .B1(n62), .B2(pc_id_i[16]), 
        .ZN(n996) );
  AOI22_X1 U1789 ( .A1(n67), .A2(uepc_o[16]), .B1(n971), .B2(pc_ex_i[16]), 
        .ZN(n995) );
  OAI211_X1 U1790 ( .C1(n1409), .C2(n967), .A(n996), .B(n995), .ZN(uepc_n[16])
         );
  AOI22_X1 U1791 ( .A1(n63), .A2(pc_ex_i[17]), .B1(n62), .B2(pc_id_i[17]), 
        .ZN(n998) );
  AOI22_X1 U1794 ( .A1(n64), .A2(pc_if_i[18]), .B1(n62), .B2(pc_id_i[18]), 
        .ZN(n1000) );
  AOI22_X1 U1797 ( .A1(n64), .A2(pc_if_i[19]), .B1(n63), .B2(pc_ex_i[19]), 
        .ZN(n1002) );
  AOI22_X1 U1800 ( .A1(n64), .A2(pc_if_i[20]), .B1(n62), .B2(pc_id_i[20]), 
        .ZN(n1004) );
  AOI22_X1 U1804 ( .A1(n63), .A2(pc_ex_i[21]), .B1(n62), .B2(pc_id_i[21]), 
        .ZN(n1006) );
  INV_X1 U1807 ( .A(n1007), .ZN(n1414) );
  AOI22_X1 U1808 ( .A1(n63), .A2(pc_ex_i[22]), .B1(n62), .B2(pc_id_i[22]), 
        .ZN(n1009) );
  INV_X1 U1811 ( .A(hwlp_data_o[23]), .ZN(n1415) );
  AOI22_X1 U1812 ( .A1(n64), .A2(pc_if_i[23]), .B1(n62), .B2(pc_id_i[23]), 
        .ZN(n1011) );
  INV_X1 U1818 ( .A(hwlp_data_o[25]), .ZN(n1418) );
  AOI22_X1 U1823 ( .A1(n64), .A2(pc_if_i[26]), .B1(n63), .B2(pc_ex_i[26]), 
        .ZN(n1018) );
  AOI22_X1 U1826 ( .A1(n64), .A2(pc_if_i[27]), .B1(n62), .B2(pc_id_i[27]), 
        .ZN(n1020) );
  AOI22_X1 U1829 ( .A1(n64), .A2(pc_if_i[28]), .B1(n62), .B2(pc_id_i[28]), 
        .ZN(n1022) );
  AOI22_X1 U1832 ( .A1(n64), .A2(pc_if_i[29]), .B1(n63), .B2(pc_ex_i[29]), 
        .ZN(n1024) );
  AOI22_X1 U1838 ( .A1(n64), .A2(pc_if_i[31]), .B1(n63), .B2(pc_ex_i[31]), 
        .ZN(n1028) );
  NOR2_X1 U1841 ( .A1(n1122), .A2(n1039), .ZN(n1037) );
  AND2_X1 U1843 ( .A1(n1385), .A2(n1029), .ZN(n1041) );
  NOR2_X1 U1859 ( .A1(n1039), .A2(n1038), .ZN(n1045) );
  NOR2_X1 U1864 ( .A1(n1394), .A2(n1054), .ZN(n1049) );
  AND2_X1 U1865 ( .A1(debug_csr_save_i), .A2(n1047), .ZN(n1048) );
  AOI21_X1 U1868 ( .B1(n1049), .B2(n3700), .A(n1677), .ZN(n1090) );
  NOR2_X1 U1869 ( .A1(n1050), .A2(n1124), .ZN(n1057) );
  NOR2_X1 U1871 ( .A1(csr_save_ex_i_BAR), .A2(n1050), .ZN(n1070) );
  NOR2_X1 U1872 ( .A1(n1050), .A2(n1126), .ZN(n1079) );
  AOI22_X1 U1873 ( .A1(pc_ex_i[0]), .A2(n55), .B1(pc_id_i[0]), .B2(n57), .ZN(
        n1051) );
  OR3_X1 U1875 ( .A1(n1198), .A2(n1054), .A3(n1677), .ZN(n1107) );
  AOI22_X1 U1876 ( .A1(pc_id_i[1]), .A2(n57), .B1(pc_if_i[1]), .B2(n56), .ZN(
        n1056) );
  AOI22_X1 U1879 ( .A1(n55), .A2(pc_ex_i[2]), .B1(n56), .B2(pc_if_i[2]), .ZN(
        n1059) );
  AOI22_X1 U1882 ( .A1(n55), .A2(pc_ex_i[3]), .B1(n56), .B2(pc_if_i[3]), .ZN(
        n1061) );
  AOI22_X1 U1888 ( .A1(pc_id_i[5]), .A2(n57), .B1(pc_if_i[5]), .B2(n56), .ZN(
        n1065) );
  AOI22_X1 U1891 ( .A1(n55), .A2(pc_ex_i[6]), .B1(n56), .B2(pc_if_i[6]), .ZN(
        n1067) );
  AOI22_X1 U1894 ( .A1(n55), .A2(pc_ex_i[7]), .B1(n57), .B2(pc_id_i[7]), .ZN(
        n1069) );
  AOI22_X1 U1897 ( .A1(n56), .A2(pc_if_i[8]), .B1(n57), .B2(pc_id_i[8]), .ZN(
        n1072) );
  AOI22_X1 U1900 ( .A1(n56), .A2(pc_if_i[9]), .B1(n57), .B2(pc_id_i[9]), .ZN(
        n1074) );
  AOI22_X1 U1903 ( .A1(n56), .A2(pc_if_i[10]), .B1(n57), .B2(pc_id_i[10]), 
        .ZN(n1076) );
  AOI22_X1 U1906 ( .A1(n55), .A2(pc_ex_i[11]), .B1(n57), .B2(pc_id_i[11]), 
        .ZN(n1078) );
  AOI22_X1 U1909 ( .A1(n55), .A2(pc_ex_i[12]), .B1(n57), .B2(pc_id_i[12]), 
        .ZN(n1081) );
  AOI22_X1 U1915 ( .A1(n55), .A2(pc_ex_i[14]), .B1(n57), .B2(pc_id_i[14]), 
        .ZN(n1085) );
  AOI22_X1 U1918 ( .A1(n55), .A2(pc_ex_i[15]), .B1(n57), .B2(pc_id_i[15]), 
        .ZN(n1087) );
  AOI22_X1 U1921 ( .A1(n55), .A2(pc_ex_i[16]), .B1(n57), .B2(pc_id_i[16]), 
        .ZN(n1089) );
  AOI22_X1 U1922 ( .A1(n1090), .A2(depc_o[16]), .B1(n56), .B2(pc_if_i[16]), 
        .ZN(n1088) );
  OAI211_X1 U1923 ( .C1(n1409), .C2(n1107), .A(n1089), .B(n1088), .ZN(
        depc_n[16]) );
  AOI22_X1 U1924 ( .A1(n55), .A2(pc_ex_i[17]), .B1(n1079), .B2(pc_id_i[17]), 
        .ZN(n1092) );
  AOI22_X1 U1925 ( .A1(n1090), .A2(depc_o[17]), .B1(n56), .B2(pc_if_i[17]), 
        .ZN(n1091) );
  OAI211_X1 U1926 ( .C1(n1410), .C2(n1107), .A(n1092), .B(n1091), .ZN(
        depc_n[17]) );
  AOI22_X1 U1927 ( .A1(n56), .A2(pc_if_i[18]), .B1(n57), .B2(pc_id_i[18]), 
        .ZN(n1094) );
  AOI22_X1 U1930 ( .A1(n56), .A2(pc_if_i[19]), .B1(n57), .B2(pc_id_i[19]), 
        .ZN(n1096) );
  AOI22_X1 U1933 ( .A1(n56), .A2(pc_if_i[20]), .B1(n57), .B2(pc_id_i[20]), 
        .ZN(n1098) );
  AOI22_X1 U1936 ( .A1(n55), .A2(pc_ex_i[21]), .B1(n56), .B2(pc_if_i[21]), 
        .ZN(n1100) );
  AOI22_X1 U1939 ( .A1(pc_if_i[22]), .A2(n56), .B1(pc_id_i[22]), .B2(n57), 
        .ZN(n1102) );
  AOI22_X1 U1945 ( .A1(n56), .A2(pc_if_i[24]), .B1(n57), .B2(pc_id_i[24]), 
        .ZN(n1106) );
  AOI22_X1 U1948 ( .A1(pc_id_i[25]), .A2(n57), .B1(pc_ex_i[25]), .B2(n55), 
        .ZN(n1109) );
  AOI22_X1 U1954 ( .A1(n56), .A2(pc_if_i[27]), .B1(n57), .B2(pc_id_i[27]), 
        .ZN(n1113) );
  AOI22_X1 U1957 ( .A1(n55), .A2(pc_ex_i[28]), .B1(n57), .B2(pc_id_i[28]), 
        .ZN(n1115) );
  AOI22_X1 U1963 ( .A1(n55), .A2(pc_ex_i[30]), .B1(n1057), .B2(pc_if_i[30]), 
        .ZN(n1119) );
  AOI22_X1 U1964 ( .A1(n1090), .A2(depc_o[30]), .B1(n57), .B2(pc_id_i[30]), 
        .ZN(n1118) );
  OAI211_X1 U1965 ( .C1(n1426), .C2(n1107), .A(n1119), .B(n1118), .ZN(
        depc_n[30]) );
  NOR2_X1 U1969 ( .A1(n1130), .A2(n1198), .ZN(n1123) );
  NOR2_X1 U1971 ( .A1(n1123), .A2(n1129), .ZN(n1166) );
  NOR2_X1 U1973 ( .A1(n1124), .A2(n1125), .ZN(n1142) );
  NOR2_X1 U1976 ( .A1(n1126), .A2(n1125), .ZN(n1155) );
  AOI22_X1 U1977 ( .A1(pc_ex_i[0]), .A2(n1141), .B1(pc_id_i[0]), .B2(n60), 
        .ZN(n1127) );
  OR3_X1 U1979 ( .A1(n1198), .A2(n1130), .A3(n1129), .ZN(n1183) );
  AOI22_X1 U1980 ( .A1(pc_id_i[1]), .A2(n60), .B1(pc_if_i[1]), .B2(n58), .ZN(
        n1132) );
  AOI22_X1 U1983 ( .A1(n58), .A2(pc_if_i[2]), .B1(n60), .B2(pc_id_i[2]), .ZN(
        n1134) );
  AOI22_X1 U1986 ( .A1(n58), .A2(pc_if_i[3]), .B1(n60), .B2(pc_id_i[3]), .ZN(
        n1136) );
  AOI22_X1 U1992 ( .A1(pc_if_i[5]), .A2(n58), .B1(pc_ex_i[5]), .B2(n1141), 
        .ZN(n1140) );
  AOI22_X1 U1995 ( .A1(n1141), .A2(pc_ex_i[6]), .B1(n60), .B2(pc_id_i[6]), 
        .ZN(n1144) );
  AOI22_X1 U2001 ( .A1(n1141), .A2(pc_ex_i[8]), .B1(n60), .B2(pc_id_i[8]), 
        .ZN(n1148) );
  AOI22_X1 U2010 ( .A1(n58), .A2(pc_if_i[11]), .B1(n60), .B2(pc_id_i[11]), 
        .ZN(n1154) );
  AOI22_X1 U2013 ( .A1(n58), .A2(pc_if_i[12]), .B1(n60), .B2(pc_id_i[12]), 
        .ZN(n1157) );
  AOI22_X1 U2016 ( .A1(n58), .A2(pc_if_i[13]), .B1(n60), .B2(pc_id_i[13]), 
        .ZN(n1159) );
  AOI22_X1 U2019 ( .A1(n1141), .A2(pc_ex_i[14]), .B1(n58), .B2(pc_if_i[14]), 
        .ZN(n1161) );
  AOI22_X1 U2022 ( .A1(n1141), .A2(pc_ex_i[15]), .B1(n60), .B2(pc_id_i[15]), 
        .ZN(n1163) );
  AOI22_X1 U2025 ( .A1(n1141), .A2(pc_ex_i[16]), .B1(n60), .B2(pc_id_i[16]), 
        .ZN(n1165) );
  AOI22_X1 U2026 ( .A1(n1166), .A2(mepc_o[16]), .B1(n58), .B2(pc_if_i[16]), 
        .ZN(n1164) );
  OAI211_X1 U2027 ( .C1(n1409), .C2(n1183), .A(n1165), .B(n1164), .ZN(
        mepc_n[16]) );
  AOI22_X1 U2028 ( .A1(n1141), .A2(pc_ex_i[17]), .B1(n1155), .B2(pc_id_i[17]), 
        .ZN(n1168) );
  AOI22_X1 U2029 ( .A1(n1166), .A2(mepc_o[17]), .B1(n58), .B2(pc_if_i[17]), 
        .ZN(n1167) );
  OAI211_X1 U2030 ( .C1(n1410), .C2(n1183), .A(n1168), .B(n1167), .ZN(
        mepc_n[17]) );
  AOI22_X1 U2031 ( .A1(n1141), .A2(pc_ex_i[18]), .B1(n60), .B2(pc_id_i[18]), 
        .ZN(n1170) );
  AOI22_X1 U2034 ( .A1(n58), .A2(pc_if_i[19]), .B1(n60), .B2(pc_id_i[19]), 
        .ZN(n1172) );
  AOI22_X1 U2037 ( .A1(n1141), .A2(pc_ex_i[20]), .B1(n58), .B2(pc_if_i[20]), 
        .ZN(n1174) );
  AOI22_X1 U2043 ( .A1(pc_ex_i[22]), .A2(n1141), .B1(pc_id_i[22]), .B2(n60), 
        .ZN(n1178) );
  AOI22_X1 U2049 ( .A1(n58), .A2(pc_if_i[24]), .B1(n60), .B2(pc_id_i[24]), 
        .ZN(n1182) );
  AOI22_X1 U2050 ( .A1(n1166), .A2(mepc_o[24]), .B1(n1141), .B2(pc_ex_i[24]), 
        .ZN(n1181) );
  OAI211_X1 U2051 ( .C1(n1416), .C2(n1183), .A(n1182), .B(n1181), .ZN(
        mepc_n[24]) );
  AOI22_X1 U2052 ( .A1(pc_id_i[25]), .A2(n60), .B1(pc_ex_i[25]), .B2(n1141), 
        .ZN(n1185) );
  NOR2_X1 U2095 ( .A1(n1223), .A2(n1225), .ZN(hwlp_we_o[0]) );
  NOR2_X1 U2096 ( .A1(n1224), .A2(n1225), .ZN(hwlp_we_o[1]) );
  NOR2_X1 U2097 ( .A1(n1226), .A2(n1225), .ZN(hwlp_we_o[2]) );
  OAI211_X1 U2098 ( .C1(n1362), .C2(n1473), .A(csr_wdata_i[2]), .B(n1231), 
        .ZN(n1227) );
  OAI21_X1 U2099 ( .B1(n1233), .B2(n1473), .A(n1227), .ZN(PCER_n[2]) );
  OAI211_X1 U2100 ( .C1(n1362), .C2(n1475), .A(csr_wdata_i[3]), .B(n1231), 
        .ZN(n1228) );
  OAI21_X1 U2101 ( .B1(n1233), .B2(n1475), .A(n1228), .ZN(PCER_n[3]) );
  OAI211_X1 U2102 ( .C1(n1362), .C2(n1474), .A(csr_wdata_i[7]), .B(n1231), 
        .ZN(n1229) );
  OAI21_X1 U2103 ( .B1(n1233), .B2(n1474), .A(n1229), .ZN(PCER_n[7]) );
  OAI211_X1 U2104 ( .C1(n1362), .C2(n1476), .A(csr_wdata_i[8]), .B(n1231), 
        .ZN(n1230) );
  OAI21_X1 U2105 ( .B1(n1233), .B2(n1476), .A(n1230), .ZN(PCER_n[8]) );
  OAI211_X1 U2106 ( .C1(n1362), .C2(n1477), .A(csr_wdata_i[9]), .B(n1231), 
        .ZN(n1232) );
  OAI21_X1 U2107 ( .B1(n1233), .B2(n1477), .A(n1232), .ZN(PCER_n[9]) );
  OAI211_X1 U2108 ( .C1(n1362), .C2(n1584), .A(csr_wdata_i[1]), .B(n1385), 
        .ZN(n1234) );
  OAI22_X1 U2109 ( .A1(n1236), .A2(n1584), .B1(n1235), .B2(n1234), .ZN(
        PCMR_n[1]) );
  OAI211_X1 U2110 ( .C1(n1362), .C2(n1498), .A(csr_wdata_i[1]), .B(n1385), 
        .ZN(n1239) );
  AOI22_X1 U2111 ( .A1(PCCR_q[1]), .A2(n1298), .B1(n1271), .B2(n1237), .ZN(
        n1238) );
  OAI21_X1 U2112 ( .B1(n1240), .B2(n1239), .A(n1238), .ZN(PCCR_n[0]) );
  OAI21_X1 U2113 ( .B1(n1362), .B2(n1452), .A(csr_wdata_i[2]), .ZN(n1243) );
  HA_X1 U2114 ( .A(PCCR_q[0]), .B(PCCR_q[1]), .CO(n1244), .S(n1237) );
  AOI22_X1 U2115 ( .A1(PCCR_q[2]), .A2(n1298), .B1(n1271), .B2(n1241), .ZN(
        n1242) );
  OAI21_X1 U2116 ( .B1(n1243), .B2(n1368), .A(n1242), .ZN(PCCR_n[1]) );
  OAI21_X1 U2117 ( .B1(n1362), .B2(n1460), .A(csr_wdata_i[3]), .ZN(n1247) );
  HA_X1 U2118 ( .A(n1244), .B(PCCR_q[2]), .CO(n1248), .S(n1241) );
  AOI22_X1 U2119 ( .A1(PCCR_q[3]), .A2(n1298), .B1(n1271), .B2(n1245), .ZN(
        n1246) );
  OAI21_X1 U2120 ( .B1(n1247), .B2(n1368), .A(n1246), .ZN(PCCR_n[2]) );
  OAI21_X1 U2121 ( .B1(n1362), .B2(n1492), .A(csr_wdata_i[4]), .ZN(n1251) );
  HA_X1 U2122 ( .A(n1248), .B(PCCR_q[3]), .CO(n1252), .S(n1245) );
  AOI22_X1 U2123 ( .A1(PCCR_q[4]), .A2(n1298), .B1(n1271), .B2(n1249), .ZN(
        n1250) );
  OAI21_X1 U2124 ( .B1(n1251), .B2(n1368), .A(n1250), .ZN(PCCR_n[3]) );
  OAI21_X1 U2125 ( .B1(n1362), .B2(n1482), .A(csr_wdata_i[5]), .ZN(n1255) );
  HA_X1 U2126 ( .A(n1252), .B(PCCR_q[4]), .CO(n1259), .S(n1249) );
  AOI22_X1 U2127 ( .A1(PCCR_q[5]), .A2(n1298), .B1(n1271), .B2(n1253), .ZN(
        n1254) );
  OAI21_X1 U2128 ( .B1(n1368), .B2(n1255), .A(n1254), .ZN(PCCR_n[4]) );
  AOI21_X1 U2129 ( .B1(n1257), .B2(PCCR_q[6]), .A(n1256), .ZN(n1258) );
  INV_X1 U2130 ( .A(n1258), .ZN(n1262) );
  HA_X1 U2131 ( .A(n1259), .B(PCCR_q[5]), .CO(n1263), .S(n1253) );
  AOI22_X1 U2132 ( .A1(PCCR_q[6]), .A2(n1298), .B1(n1271), .B2(n1260), .ZN(
        n1261) );
  OAI21_X1 U2133 ( .B1(n1262), .B2(n1368), .A(n1261), .ZN(PCCR_n[5]) );
  OAI21_X1 U2134 ( .B1(n1362), .B2(n1499), .A(csr_wdata_i[7]), .ZN(n1266) );
  HA_X1 U2135 ( .A(n1263), .B(PCCR_q[6]), .CO(n1267), .S(n1260) );
  AOI22_X1 U2136 ( .A1(PCCR_q[7]), .A2(n1298), .B1(n1271), .B2(n1264), .ZN(
        n1265) );
  OAI21_X1 U2137 ( .B1(n1266), .B2(n1368), .A(n1265), .ZN(PCCR_n[6]) );
  OAI21_X1 U2138 ( .B1(n1362), .B2(n1463), .A(csr_wdata_i[8]), .ZN(n1270) );
  HA_X1 U2139 ( .A(n1267), .B(PCCR_q[7]), .CO(n1272), .S(n1264) );
  AOI22_X1 U2140 ( .A1(PCCR_q[8]), .A2(n1298), .B1(n1366), .B2(n1268), .ZN(
        n1269) );
  OAI21_X1 U2141 ( .B1(n1270), .B2(n1368), .A(n1269), .ZN(PCCR_n[7]) );
  OAI21_X1 U2142 ( .B1(n1362), .B2(n1500), .A(csr_wdata_i[9]), .ZN(n1275) );
  CLKBUF_X1 U2143 ( .A(n1271), .Z(n1366) );
  HA_X1 U2144 ( .A(n1272), .B(PCCR_q[8]), .CO(n1276), .S(n1268) );
  AOI22_X1 U2145 ( .A1(PCCR_q[9]), .A2(n1315), .B1(n1366), .B2(n1273), .ZN(
        n1274) );
  OAI21_X1 U2146 ( .B1(n1275), .B2(n1368), .A(n1274), .ZN(PCCR_n[8]) );
  OAI21_X1 U2147 ( .B1(n1362), .B2(n1493), .A(csr_wdata_i[10]), .ZN(n1279) );
  HA_X1 U2148 ( .A(n1276), .B(PCCR_q[9]), .CO(n1280), .S(n1273) );
  AOI22_X1 U2149 ( .A1(PCCR_q[10]), .A2(n1298), .B1(n1366), .B2(n1277), .ZN(
        n1278) );
  OAI21_X1 U2150 ( .B1(n1279), .B2(n1368), .A(n1278), .ZN(PCCR_n[9]) );
  OAI21_X1 U2151 ( .B1(n1362), .B2(n1501), .A(csr_wdata_i[11]), .ZN(n1283) );
  HA_X1 U2152 ( .A(n1280), .B(PCCR_q[10]), .CO(n1284), .S(n1277) );
  AOI22_X1 U2153 ( .A1(PCCR_q[11]), .A2(n1298), .B1(n1366), .B2(n1281), .ZN(
        n1282) );
  OAI21_X1 U2154 ( .B1(n1283), .B2(n1368), .A(n1282), .ZN(PCCR_n[10]) );
  OAI21_X1 U2155 ( .B1(n1362), .B2(n1462), .A(csr_wdata_i[12]), .ZN(n1287) );
  HA_X1 U2156 ( .A(n1284), .B(PCCR_q[11]), .CO(n1288), .S(n1281) );
  AOI22_X1 U2157 ( .A1(PCCR_q[12]), .A2(n1298), .B1(n1366), .B2(n1285), .ZN(
        n1286) );
  OAI21_X1 U2158 ( .B1(n1287), .B2(n1368), .A(n1286), .ZN(PCCR_n[11]) );
  OAI21_X1 U2159 ( .B1(n1362), .B2(n1487), .A(csr_wdata_i[13]), .ZN(n1291) );
  HA_X1 U2160 ( .A(n1288), .B(PCCR_q[12]), .CO(n1292), .S(n1285) );
  AOI22_X1 U2161 ( .A1(PCCR_q[13]), .A2(n1298), .B1(n1366), .B2(n1289), .ZN(
        n1290) );
  OAI21_X1 U2162 ( .B1(n1291), .B2(n1368), .A(n1290), .ZN(PCCR_n[12]) );
  OAI21_X1 U2163 ( .B1(n1362), .B2(n1483), .A(csr_wdata_i[14]), .ZN(n1295) );
  HA_X1 U2164 ( .A(n1292), .B(PCCR_q[13]), .CO(n1296), .S(n1289) );
  AOI22_X1 U2165 ( .A1(PCCR_q[14]), .A2(n1298), .B1(n1366), .B2(n1293), .ZN(
        n1294) );
  OAI21_X1 U2166 ( .B1(n1295), .B2(n1368), .A(n1294), .ZN(PCCR_n[13]) );
  OAI21_X1 U2167 ( .B1(n1362), .B2(n1484), .A(csr_wdata_i[15]), .ZN(n1300) );
  HA_X1 U2168 ( .A(n1296), .B(PCCR_q[14]), .CO(n1301), .S(n1293) );
  AOI22_X1 U2169 ( .A1(PCCR_q[15]), .A2(n1298), .B1(n1366), .B2(n1297), .ZN(
        n1299) );
  OAI21_X1 U2170 ( .B1(n1300), .B2(n1368), .A(n1299), .ZN(PCCR_n[14]) );
  OAI21_X1 U2171 ( .B1(n1362), .B2(n1488), .A(csr_wdata_i[16]), .ZN(n1304) );
  HA_X1 U2172 ( .A(n1301), .B(PCCR_q[15]), .CO(n1305), .S(n1297) );
  AOI22_X1 U2173 ( .A1(PCCR_q[16]), .A2(n1315), .B1(n1366), .B2(n1302), .ZN(
        n1303) );
  OAI21_X1 U2174 ( .B1(n1304), .B2(n1368), .A(n1303), .ZN(PCCR_n[15]) );
  OAI21_X1 U2175 ( .B1(n1362), .B2(n1494), .A(csr_wdata_i[17]), .ZN(n1308) );
  HA_X1 U2176 ( .A(n1305), .B(PCCR_q[16]), .CO(n1309), .S(n1302) );
  AOI22_X1 U2177 ( .A1(PCCR_q[17]), .A2(n1315), .B1(n1366), .B2(n1306), .ZN(
        n1307) );
  OAI21_X1 U2178 ( .B1(n1308), .B2(n1368), .A(n1307), .ZN(PCCR_n[16]) );
  OAI21_X1 U2179 ( .B1(n1362), .B2(n1489), .A(csr_wdata_i[18]), .ZN(n1312) );
  HA_X1 U2180 ( .A(n1309), .B(PCCR_q[17]), .CO(n1313), .S(n1306) );
  AOI22_X1 U2181 ( .A1(PCCR_q[18]), .A2(n1315), .B1(n1366), .B2(n1310), .ZN(
        n1311) );
  OAI21_X1 U2182 ( .B1(n1312), .B2(n1368), .A(n1311), .ZN(PCCR_n[17]) );
  OAI21_X1 U2183 ( .B1(n1362), .B2(n1495), .A(csr_wdata_i[19]), .ZN(n1317) );
  HA_X1 U2184 ( .A(n1313), .B(PCCR_q[18]), .CO(n1318), .S(n1310) );
  AOI22_X1 U2185 ( .A1(PCCR_q[19]), .A2(n1315), .B1(n1366), .B2(n1314), .ZN(
        n1316) );
  OAI21_X1 U2186 ( .B1(n1317), .B2(n1368), .A(n1316), .ZN(PCCR_n[18]) );
  OAI21_X1 U2187 ( .B1(n1362), .B2(n1464), .A(csr_wdata_i[20]), .ZN(n1321) );
  HA_X1 U2188 ( .A(n1318), .B(PCCR_q[19]), .CO(n1322), .S(n1314) );
  AOI22_X1 U2189 ( .A1(PCCR_q[20]), .A2(n1298), .B1(n1366), .B2(n1319), .ZN(
        n1320) );
  OAI21_X1 U2190 ( .B1(n1321), .B2(n1368), .A(n1320), .ZN(PCCR_n[19]) );
  OAI21_X1 U2191 ( .B1(n1362), .B2(n1485), .A(csr_wdata_i[21]), .ZN(n1325) );
  HA_X1 U2192 ( .A(n1322), .B(PCCR_q[20]), .CO(n1326), .S(n1319) );
  AOI22_X1 U2193 ( .A1(PCCR_q[21]), .A2(n1315), .B1(n1366), .B2(n1323), .ZN(
        n1324) );
  OAI21_X1 U2194 ( .B1(n1325), .B2(n1368), .A(n1324), .ZN(PCCR_n[20]) );
  OAI21_X1 U2195 ( .B1(n1362), .B2(n1502), .A(csr_wdata_i[22]), .ZN(n1329) );
  HA_X1 U2196 ( .A(n1326), .B(PCCR_q[21]), .CO(n1330), .S(n1323) );
  AOI22_X1 U2197 ( .A1(PCCR_q[22]), .A2(n1298), .B1(n1366), .B2(n1327), .ZN(
        n1328) );
  OAI21_X1 U2198 ( .B1(n1368), .B2(n1329), .A(n1328), .ZN(PCCR_n[21]) );
  OAI21_X1 U2199 ( .B1(n1362), .B2(n1465), .A(csr_wdata_i[23]), .ZN(n1333) );
  HA_X1 U2200 ( .A(n1330), .B(PCCR_q[22]), .CO(n1334), .S(n1327) );
  AOI22_X1 U2201 ( .A1(PCCR_q[23]), .A2(n1315), .B1(n1366), .B2(n1331), .ZN(
        n1332) );
  OAI21_X1 U2202 ( .B1(n1333), .B2(n1368), .A(n1332), .ZN(PCCR_n[22]) );
  OAI21_X1 U2203 ( .B1(n1362), .B2(n1486), .A(csr_wdata_i[24]), .ZN(n1337) );
  HA_X1 U2204 ( .A(n1334), .B(PCCR_q[23]), .CO(n1338), .S(n1331) );
  AOI22_X1 U2205 ( .A1(PCCR_q[24]), .A2(n1298), .B1(n1366), .B2(n1335), .ZN(
        n1336) );
  OAI21_X1 U2206 ( .B1(n1337), .B2(n1368), .A(n1336), .ZN(PCCR_n[23]) );
  OAI21_X1 U2207 ( .B1(n1362), .B2(n1496), .A(csr_wdata_i[25]), .ZN(n1341) );
  HA_X1 U2208 ( .A(n1338), .B(PCCR_q[24]), .CO(n1342), .S(n1335) );
  AOI22_X1 U2209 ( .A1(PCCR_q[25]), .A2(n1298), .B1(n1366), .B2(n1339), .ZN(
        n1340) );
  OAI21_X1 U2210 ( .B1(n1368), .B2(n1341), .A(n1340), .ZN(PCCR_n[24]) );
  OAI21_X1 U2211 ( .B1(n1362), .B2(n1490), .A(csr_wdata_i[26]), .ZN(n1345) );
  HA_X1 U2212 ( .A(n1342), .B(PCCR_q[25]), .CO(n1346), .S(n1339) );
  AOI22_X1 U2213 ( .A1(PCCR_q[26]), .A2(n1315), .B1(n1366), .B2(n1343), .ZN(
        n1344) );
  OAI21_X1 U2214 ( .B1(n1345), .B2(n1368), .A(n1344), .ZN(PCCR_n[25]) );
  OAI21_X1 U2215 ( .B1(n1362), .B2(n1503), .A(csr_wdata_i[27]), .ZN(n1349) );
  HA_X1 U2216 ( .A(n1346), .B(PCCR_q[26]), .CO(n1350), .S(n1343) );
  AOI22_X1 U2217 ( .A1(PCCR_q[27]), .A2(n1298), .B1(n1366), .B2(n1347), .ZN(
        n1348) );
  OAI21_X1 U2218 ( .B1(n1349), .B2(n1368), .A(n1348), .ZN(PCCR_n[26]) );
  OAI21_X1 U2219 ( .B1(n1362), .B2(n1497), .A(csr_wdata_i[28]), .ZN(n1353) );
  HA_X1 U2220 ( .A(n1350), .B(PCCR_q[27]), .CO(n1354), .S(n1347) );
  AOI22_X1 U2221 ( .A1(PCCR_q[28]), .A2(n1315), .B1(n1366), .B2(n1351), .ZN(
        n1352) );
  OAI21_X1 U2222 ( .B1(n1353), .B2(n1368), .A(n1352), .ZN(PCCR_n[27]) );
  OAI21_X1 U2223 ( .B1(n1362), .B2(n1491), .A(csr_wdata_i[29]), .ZN(n1357) );
  HA_X1 U2224 ( .A(n1354), .B(PCCR_q[28]), .CO(n1358), .S(n1351) );
  AOI22_X1 U2225 ( .A1(PCCR_q[29]), .A2(n1298), .B1(n1366), .B2(n1355), .ZN(
        n1356) );
  OAI21_X1 U2226 ( .B1(n1357), .B2(n1368), .A(n1356), .ZN(PCCR_n[28]) );
  OAI21_X1 U2227 ( .B1(n1362), .B2(n1466), .A(csr_wdata_i[30]), .ZN(n1361) );
  HA_X1 U2228 ( .A(n1358), .B(PCCR_q[29]), .CO(n1363), .S(n1355) );
  AOI22_X1 U2229 ( .A1(PCCR_q[30]), .A2(n1315), .B1(n1271), .B2(n1359), .ZN(
        n1360) );
  OAI21_X1 U2230 ( .B1(n1361), .B2(n1368), .A(n1360), .ZN(PCCR_n[29]) );
  OAI21_X1 U2231 ( .B1(n1362), .B2(n1505), .A(csr_wdata_i[31]), .ZN(n1369) );
  HA_X1 U2232 ( .A(n1363), .B(PCCR_q[30]), .CO(n1364), .S(n1359) );
  XOR2_X1 U2233 ( .A(n1364), .B(PCCR_q[31]), .Z(n1365) );
  AOI22_X1 U2234 ( .A1(PCCR_q[31]), .A2(n1298), .B1(n1366), .B2(n1365), .ZN(
        n1367) );
  OAI21_X1 U2235 ( .B1(n1369), .B2(n1368), .A(n1367), .ZN(PCCR_n[30]) );
  NAND2_X1 U2237 ( .A1(n1706), .A2(n3700), .ZN(n1401) );
  NOR2_X1 U2238 ( .A1(n1380), .A2(n1401), .ZN(n1384) );
  NAND3_X1 U2239 ( .A1(n1371), .A2(n1373), .A3(n1372), .ZN(n1383) );
  AND2_X1 U2240 ( .A1(n1384), .A2(n1383), .ZN(n1428) );
  NAND3_X1 U2241 ( .A1(n1375), .A2(n1428), .A3(n1385), .ZN(n1377) );
  OR2_X1 U2242 ( .A1(n1374), .A2(n1377), .ZN(n1434) );
  NAND3_X1 U2243 ( .A1(csr_addr_i[1]), .A2(n1373), .A3(n1372), .ZN(n1396) );
  INV_X1 U2244 ( .A(n1398), .ZN(n1376) );
  NOR2_X1 U2245 ( .A1(n70), .A2(n1377), .ZN(n1419) );
  NOR2_X1 U2248 ( .A1(n1429), .A2(n1395), .ZN(n1379) );
  NAND3_X1 U2249 ( .A1(n1379), .A2(n1385), .A3(n1383), .ZN(n1400) );
  OR3_X1 U2250 ( .A1(n1380), .A2(csr_addr_i[11]), .A3(n1400), .ZN(n1382) );
  INV_X1 U2254 ( .A(n1383), .ZN(n1386) );
  NOR2_X1 U2277 ( .A1(n1395), .A2(n1394), .ZN(n1427) );
  NAND3_X1 U2278 ( .A1(n1396), .A2(n3700), .A3(n1427), .ZN(n1397) );
  NOR3_X1 U2279 ( .A1(n1398), .A2(n70), .A3(n1397), .ZN(n1399) );
  INV_X1 U2280 ( .A(n1399), .ZN(n1424) );
  NOR3_X1 U2286 ( .A1(n70), .A2(n1401), .A3(n1400), .ZN(n1403) );
  OAI22_X1 U2301 ( .A1(n1404), .A2(n1438), .B1(n1437), .B2(n1579), .ZN(n2764)
         );
  OAI22_X1 U2305 ( .A1(n1405), .A2(n1434), .B1(n1419), .B2(n1580), .ZN(n2761)
         );
  OAI22_X1 U2325 ( .A1(n1419), .A2(n1622), .B1(n1409), .B2(n1434), .ZN(n2741)
         );
  OAI22_X1 U2329 ( .A1(n1399), .A2(n1520), .B1(n1410), .B2(n1424), .ZN(n2737)
         );
  OAI22_X1 U2333 ( .A1(n1403), .A2(n1544), .B1(n1410), .B2(n1440), .ZN(n2733)
         );
  OAI22_X1 U2406 ( .A1(n1441), .A2(n1440), .B1(n1403), .B2(n1469), .ZN(n2663)
         );
  AOI22_X1 U2408 ( .A1(n1445), .A2(n1444), .B1(n1478), .B2(n1443), .ZN(n2136)
         );
  SDFFR_X1 dcsr_q_reg_xdebugver__30_ ( .D(1'b1), .SI(1'b0), .SE(1'b0), .CK(
        n3946), .RN(rst_n), .Q(dcsr_q_xdebugver__30_) );
  SDFFR_X1 PCER_q_reg_11_ ( .D(PCER_n[11]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .RN(rst_n), .Q(PCER_q[11]), .QN(n1479) );
  SDFFR_X1 PCER_q_reg_10_ ( .D(PCER_n[10]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .RN(rst_n), .Q(PCER_q[10]), .QN(n1480) );
  SDFFR_X1 PCER_q_reg_9_ ( .D(PCER_n[9]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .RN(rst_n), .Q(PCER_q[9]), .QN(n1477) );
  SDFFR_X1 PCER_q_reg_8_ ( .D(PCER_n[8]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .RN(rst_n), .Q(PCER_q[8]), .QN(n1476) );
  SDFFR_X1 PCER_q_reg_7_ ( .D(PCER_n[7]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .RN(rst_n), .Q(PCER_q[7]), .QN(n1474) );
  SDFFR_X1 PCER_q_reg_6_ ( .D(PCER_n[6]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .RN(rst_n), .Q(PCER_q[6]), .QN(n1472) );
  SDFFR_X1 PCER_q_reg_5_ ( .D(PCER_n[5]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .RN(rst_n), .Q(PCER_q[5]), .QN(n1471) );
  SDFFR_X1 PCER_q_reg_4_ ( .D(PCER_n[4]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .RN(rst_n), .Q(PCER_q[4]), .QN(n1457) );
  SDFFR_X1 PCER_q_reg_3_ ( .D(PCER_n[3]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .RN(rst_n), .Q(PCER_q[3]), .QN(n1475) );
  SDFFR_X1 PCER_q_reg_2_ ( .D(PCER_n[2]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .RN(rst_n), .Q(PCER_q[2]), .QN(n1473) );
  SDFFR_X1 PCER_q_reg_1_ ( .D(PCER_n[1]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .RN(rst_n), .Q(PCER_q[1]), .QN(n1458) );
  SDFFR_X1 PCER_q_reg_0_ ( .D(PCER_n[0]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .RN(rst_n), .Q(PCER_q[0]), .QN(n1468) );
  SDFFR_X1 PCCR_inc_q_reg_0_ ( .D(PCCR_inc_0_), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(rst_n), .Q(PCCR_inc_q_0_) );
  SDFFR_X1 PCCR_q_reg_0__1_ ( .D(PCCR_n[0]), .SI(1'b0), .SE(1'b0), .CK(n3914), 
        .RN(rst_n), .Q(PCCR_q[1]), .QN(n1498) );
  SDFFR_X1 PCCR_q_reg_0__2_ ( .D(PCCR_n[1]), .SI(1'b0), .SE(1'b0), .CK(n3914), 
        .RN(rst_n), .Q(PCCR_q[2]), .QN(n1452) );
  SDFFR_X1 PCCR_q_reg_0__3_ ( .D(PCCR_n[2]), .SI(1'b0), .SE(1'b0), .CK(n3914), 
        .RN(rst_n), .Q(PCCR_q[3]), .QN(n1460) );
  SDFFR_X1 PCCR_q_reg_0__4_ ( .D(PCCR_n[3]), .SI(1'b0), .SE(1'b0), .CK(n3914), 
        .RN(rst_n), .Q(PCCR_q[4]), .QN(n1492) );
  SDFFR_X1 PCCR_q_reg_0__5_ ( .D(PCCR_n[4]), .SI(1'b0), .SE(1'b0), .CK(n3914), 
        .RN(rst_n), .Q(PCCR_q[5]), .QN(n1482) );
  SDFFR_X1 PCCR_q_reg_0__6_ ( .D(PCCR_n[5]), .SI(1'b0), .SE(1'b0), .CK(n3914), 
        .RN(rst_n), .Q(PCCR_q[6]) );
  SDFFR_X1 PCCR_q_reg_0__7_ ( .D(PCCR_n[6]), .SI(1'b0), .SE(1'b0), .CK(n3914), 
        .RN(rst_n), .Q(PCCR_q[7]), .QN(n1499) );
  SDFFR_X1 PCCR_q_reg_0__8_ ( .D(PCCR_n[7]), .SI(1'b0), .SE(1'b0), .CK(n3914), 
        .RN(rst_n), .Q(PCCR_q[8]), .QN(n1463) );
  SDFFR_X1 PCCR_q_reg_0__9_ ( .D(PCCR_n[8]), .SI(1'b0), .SE(1'b0), .CK(n3914), 
        .RN(rst_n), .Q(PCCR_q[9]), .QN(n1500) );
  SDFFR_X1 PCCR_q_reg_0__10_ ( .D(PCCR_n[9]), .SI(1'b0), .SE(1'b0), .CK(n3914), 
        .RN(rst_n), .Q(PCCR_q[10]), .QN(n1493) );
  SDFFR_X1 PCCR_q_reg_0__11_ ( .D(PCCR_n[10]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[11]), .QN(n1501) );
  SDFFR_X1 PCCR_q_reg_0__12_ ( .D(PCCR_n[11]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[12]), .QN(n1462) );
  SDFFR_X1 mepc_q_reg_0_ ( .D(n4034), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(n3) );
  SDFFR_X1 mepc_q_reg_11_ ( .D(n4035), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[11]) );
  SDFFR_X1 depc_q_reg_0_ ( .D(n4002), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(n5) );
  SDFFR_X1 depc_q_reg_5_ ( .D(n4003), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[5]) );
  SDFFR_X1 uepc_q_reg_5_ ( .D(n3972), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[5]) );
  SDFFR_X1 mepc_q_reg_5_ ( .D(n4036), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[5]) );
  SDFFR_X1 dcsr_q_reg_zero0_ ( .D(n970), .SI(1'b0), .SE(1'b0), .CK(n3946), 
        .RN(rst_n), .Q(dcsr_q_zero0_) );
  SDFFR_X1 mscratch_q_reg_5_ ( .D(n4068), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[5]) );
  SDFFR_X1 dscratch0_q_reg_5_ ( .D(n4103), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[5]) );
  SDFFR_X1 dscratch1_q_reg_5_ ( .D(hwlp_data_o[5]), .SI(1'b0), .SE(1'b0), .CK(
        n4101), .RN(rst_n), .Q(dscratch1_q[5]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__5_ ( .D(n970), .SI(1'b0), .SE(1'b0), .CK(
        n4149), .RN(rst_n), .Q(pmp_addr_o[5]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__5_ ( .D(n970), .SI(1'b0), .SE(1'b0), .CK(
        n4163), .RN(rst_n), .Q(pmp_addr_o[37]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__5_ ( .D(n970), .SI(1'b0), .SE(1'b0), .CK(
        n4165), .RN(rst_n), .Q(pmp_addr_o[69]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__5_ ( .D(hwlp_data_o[5]), .SI(1'b0), .SE(
        1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[101]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__5_ ( .D(hwlp_data_o[5]), .SI(1'b0), .SE(
        1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[133]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__5_ ( .D(n970), .SI(1'b0), .SE(1'b0), .CK(
        n4171), .RN(rst_n), .Q(pmp_addr_o[165]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__5_ ( .D(n970), .SI(1'b0), .SE(1'b0), .CK(
        n4173), .RN(rst_n), .Q(pmp_addr_o[197]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__5_ ( .D(hwlp_data_o[5]), .SI(1'b0), .SE(
        1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[229]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__5_ ( .D(hwlp_data_o[5]), .SI(1'b0), .SE(
        1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[261]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__5_ ( .D(n970), .SI(1'b0), .SE(1'b0), .CK(
        n4180), .RN(rst_n), .Q(pmp_addr_o[293]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__5_ ( .D(n970), .SI(1'b0), .SE(1'b0), 
        .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[325]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__5_ ( .D(hwlp_data_o[5]), .SI(1'b0), .SE(
        1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[357]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__5_ ( .D(hwlp_data_o[5]), .SI(1'b0), .SE(
        1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[389]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__5_ ( .D(n970), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[421]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__5_ ( .D(n970), .SI(1'b0), .SE(1'b0), 
        .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[453]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__5_ ( .D(hwlp_data_o[5]), .SI(1'b0), .SE(
        1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[485]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__0__5_ ( .D(hwlp_data_o[5]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(n53) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__4__5_ ( .D(hwlp_data_o[5]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(n41) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__8__5_ ( .D(n970), .SI(1'b0), .SE(1'b0), .CK(
        n3964), .RN(rst_n), .Q(n29) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__12__5_ ( .D(n2051), .SI(1'b0), .SE(1'b0), 
        .CK(n3967), .RN(rst_n), .Q(n17) );
  SDFFR_X1 depc_q_reg_9_ ( .D(n4004), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[9]) );
  SDFFR_X1 uepc_q_reg_9_ ( .D(n3973), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[9]) );
  SDFFR_X1 mepc_q_reg_9_ ( .D(n4037), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[9]) );
  SDFFR_X1 mtvec_q_reg_1_ ( .D(n1681), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[1]), .QN(n1553) );
  SDFFR_X1 mscratch_q_reg_9_ ( .D(n4069), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[9]) );
  SDFFR_X1 dscratch0_q_reg_9_ ( .D(n4105), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[9]) );
  SDFFR_X1 dscratch1_q_reg_9_ ( .D(n1681), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[9]) );
  SDFFR_X1 utvec_q_reg_1_ ( .D(n1681), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[1]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[9]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[41]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[73]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[105]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[137]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[169]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[201]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[233]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[265]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[297]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[329]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[361]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[393]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[425]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[457]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__9_ ( .D(hwlp_data_o[9]), .SI(1'b0), .SE(
        1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[489]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__1__1_ ( .D(n2135), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(pmp_cfg_o[9]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__5__1_ ( .D(n2103), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(pmp_cfg_o[41]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__9__1_ ( .D(n2071), .SI(1'b0), .SE(1'b0), .CK(
        n3964), .RN(rst_n), .Q(pmp_cfg_o[73]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__13__1_ ( .D(n1681), .SI(1'b0), .SE(1'b0), 
        .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[105]) );
  SDFFR_X1 depc_q_reg_10_ ( .D(n4005), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[10]) );
  SDFFR_X1 uepc_q_reg_10_ ( .D(n3974), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[10]) );
  SDFFR_X1 mepc_q_reg_10_ ( .D(n4039), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[10]) );
  SDFFR_X1 mtvec_q_reg_2_ ( .D(n1682), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[2]) );
  SDFFR_X1 mscratch_q_reg_10_ ( .D(n4070), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[10]) );
  SDFFR_X1 dscratch0_q_reg_10_ ( .D(n4106), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[10]) );
  SDFFR_X1 dscratch1_q_reg_10_ ( .D(n1682), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[10]) );
  SDFFR_X1 utvec_q_reg_2_ ( .D(n1682), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[2]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[10]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[42]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[74]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[106]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[138]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[170]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[202]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[234]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[266]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[298]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[330]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[362]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[394]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[426]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[458]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__10_ ( .D(hwlp_data_o[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[490]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__1__2_ ( .D(n2136), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(pmp_cfg_o[10]), .QN(n1478) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__5__2_ ( .D(hwlp_data_o[10]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(pmp_cfg_o[42]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__9__2_ ( .D(hwlp_data_o[10]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[74]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__13__2_ ( .D(hwlp_data_o[10]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[106]) );
  SDFFR_X1 dcsr_q_reg_cause__6_ ( .D(n3917), .SI(1'b0), .SE(1'b0), .CK(n3922), 
        .RN(rst_n), .Q(dcsr_q_cause__6_) );
  SDFFR_X1 uepc_q_reg_6_ ( .D(n3975), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[6]) );
  SDFFR_X1 depc_q_reg_6_ ( .D(n4006), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[6]) );
  SDFFR_X1 mepc_q_reg_6_ ( .D(n4040), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[6]) );
  SDFFR_X1 mscratch_q_reg_6_ ( .D(n4071), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[6]) );
  SDFFR_X1 dscratch0_q_reg_6_ ( .D(n4107), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[6]) );
  SDFFR_X1 dscratch1_q_reg_6_ ( .D(hwlp_data_o[6]), .SI(1'b0), .SE(1'b0), .CK(
        n4101), .RN(rst_n), .Q(dscratch1_q[6]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__6_ ( .D(hwlp_data_o[6]), .SI(1'b0), .SE(
        1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[6]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__6_ ( .D(hwlp_data_o[6]), .SI(1'b0), .SE(
        1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[38]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__6_ ( .D(hwlp_data_o[6]), .SI(1'b0), .SE(
        1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[70]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__6_ ( .D(hwlp_data_o[6]), .SI(1'b0), .SE(
        1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[102]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__6_ ( .D(hwlp_data_o[6]), .SI(1'b0), .SE(
        1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[134]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__6_ ( .D(hwlp_data_o[6]), .SI(1'b0), .SE(
        1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[166]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__6_ ( .D(hwlp_data_o[6]), .SI(1'b0), .SE(
        1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[198]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__6_ ( .D(n483), .SI(1'b0), .SE(1'b0), .CK(
        n4176), .RN(rst_n), .Q(pmp_addr_o[230]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__6_ ( .D(n483), .SI(1'b0), .SE(1'b0), .CK(
        n4178), .RN(rst_n), .Q(pmp_addr_o[262]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__6_ ( .D(n483), .SI(1'b0), .SE(1'b0), .CK(
        n4180), .RN(rst_n), .Q(pmp_addr_o[294]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__6_ ( .D(n483), .SI(1'b0), .SE(1'b0), 
        .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[326]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__6_ ( .D(n483), .SI(1'b0), .SE(1'b0), 
        .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[358]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__6_ ( .D(n483), .SI(1'b0), .SE(1'b0), 
        .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[390]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__6_ ( .D(n483), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[422]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__6_ ( .D(n483), .SI(1'b0), .SE(1'b0), 
        .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[454]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__6_ ( .D(n483), .SI(1'b0), .SE(1'b0), 
        .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[486]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__0__6_ ( .D(n483), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(n52) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__4__6_ ( .D(n483), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(n40) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__8__6_ ( .D(n483), .SI(1'b0), .SE(1'b0), .CK(
        n3964), .RN(rst_n), .Q(n28) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__12__6_ ( .D(hwlp_data_o[6]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(n16) );
  SDFFR_X1 dcsr_q_reg_cause__8_ ( .D(n3918), .SI(1'b0), .SE(1'b0), .CK(n3922), 
        .RN(rst_n), .Q(dcsr_q_cause__8_) );
  SDFFR_X1 uepc_q_reg_8_ ( .D(n3976), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[8]) );
  SDFFR_X1 depc_q_reg_8_ ( .D(n4007), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[8]) );
  SDFFR_X1 mepc_q_reg_8_ ( .D(n4041), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[8]) );
  SDFFR_X1 mtvec_q_reg_0_ ( .D(hwlp_data_o[8]), .SI(1'b0), .SE(1'b0), .CK(
        n3962), .RN(rst_n), .Q(mtvec_o[0]) );
  SDFFR_X1 mscratch_q_reg_8_ ( .D(n4072), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[8]) );
  SDFFR_X1 dscratch0_q_reg_8_ ( .D(n4109), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[8]) );
  SDFFR_X1 dscratch1_q_reg_8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[8]) );
  SDFFR_X1 utvec_q_reg_0_ ( .D(n4175), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[0]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), 
        .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[8]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), 
        .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[40]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), 
        .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[72]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), 
        .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[104]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), 
        .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[136]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), 
        .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[168]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), 
        .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[200]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), 
        .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[232]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), 
        .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[264]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), 
        .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[296]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), 
        .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[328]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), 
        .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[360]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__8_ ( .D(hwlp_data_o[8]), .SI(1'b0), .SE(
        1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[392]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__8_ ( .D(hwlp_data_o[8]), .SI(1'b0), .SE(
        1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[424]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__8_ ( .D(hwlp_data_o[8]), .SI(1'b0), .SE(
        1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[456]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__8_ ( .D(n4175), .SI(1'b0), .SE(1'b0), 
        .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[488]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__1__0_ ( .D(hwlp_data_o[8]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(pmp_cfg_o[8]), .QN(n1607) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__5__0_ ( .D(hwlp_data_o[8]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(pmp_cfg_o[40]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__9__0_ ( .D(hwlp_data_o[8]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[72]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__13__0_ ( .D(hwlp_data_o[8]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[104]) );
  SDFFR_X1 mcause_q_reg_1_ ( .D(n3926), .SI(1'b0), .SE(1'b0), .CK(n3932), .RN(
        rst_n), .Q(mcause_q[1]) );
  SDFFR_X1 uepc_q_reg_1_ ( .D(n3977), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[1]) );
  SDFFR_X1 depc_q_reg_1_ ( .D(n4008), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[1]) );
  SDFFR_X1 mepc_q_reg_1_ ( .D(n4042), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[1]) );
  SDFFR_X1 ucause_q_reg_1_ ( .D(n3935), .SI(1'b0), .SE(1'b0), .CK(n3942), .RN(
        rst_n), .Q(ucause_q[1]) );
  SDFFR_X1 mscratch_q_reg_1_ ( .D(n4073), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[1]) );
  SDFFR_X1 dscratch0_q_reg_1_ ( .D(n4110), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[1]) );
  SDFFR_X1 dscratch1_q_reg_1_ ( .D(hwlp_data_o[1]), .SI(1'b0), .SE(1'b0), .CK(
        n4101), .RN(rst_n), .Q(dscratch1_q[1]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__1_ ( .D(n1031), .SI(1'b0), .SE(1'b0), 
        .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[1]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__1_ ( .D(n1031), .SI(1'b0), .SE(1'b0), 
        .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[33]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__1_ ( .D(n1031), .SI(1'b0), .SE(1'b0), 
        .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[65]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__1_ ( .D(n1031), .SI(1'b0), .SE(1'b0), 
        .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[97]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__1_ ( .D(hwlp_data_o[1]), .SI(1'b0), .SE(
        1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[129]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__1_ ( .D(hwlp_data_o[1]), .SI(1'b0), .SE(
        1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[161]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__1_ ( .D(n1031), .SI(1'b0), .SE(1'b0), 
        .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[193]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__1_ ( .D(n1031), .SI(1'b0), .SE(1'b0), 
        .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[225]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__1_ ( .D(hwlp_data_o[1]), .SI(1'b0), .SE(
        1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[257]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__1_ ( .D(hwlp_data_o[1]), .SI(1'b0), .SE(
        1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[289]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__1_ ( .D(n1031), .SI(1'b0), .SE(1'b0), 
        .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[321]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__1_ ( .D(n1031), .SI(1'b0), .SE(1'b0), 
        .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[353]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__1_ ( .D(n1031), .SI(1'b0), .SE(1'b0), 
        .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[385]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__1_ ( .D(hwlp_data_o[1]), .SI(1'b0), .SE(
        1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[449]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__0__1_ ( .D(n1031), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(pmp_cfg_o[1]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__4__1_ ( .D(hwlp_data_o[1]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(pmp_cfg_o[33]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__8__1_ ( .D(hwlp_data_o[1]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[65]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__12__1_ ( .D(hwlp_data_o[1]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[97]) );
  SDFFR_X1 mcause_q_reg_2_ ( .D(n3927), .SI(1'b0), .SE(1'b0), .CK(n3932), .RN(
        rst_n), .Q(mcause_q[2]) );
  SDFFR_X1 uepc_q_reg_2_ ( .D(n3978), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[2]) );
  SDFFR_X1 depc_q_reg_2_ ( .D(n4009), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[2]) );
  SDFFR_X1 mepc_q_reg_2_ ( .D(n4043), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[2]) );
  SDFFR_X1 ucause_q_reg_2_ ( .D(n3937), .SI(1'b0), .SE(1'b0), .CK(n3942), .RN(
        rst_n), .Q(ucause_q[2]) );
  SDFFR_X1 dcsr_q_reg_step_ ( .D(n4113), .SI(1'b0), .SE(1'b0), .CK(n3946), 
        .RN(rst_n), .Q(debug_single_step_o) );
  SDFFR_X1 mscratch_q_reg_2_ ( .D(n4074), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[2]) );
  SDFFR_X1 dscratch0_q_reg_2_ ( .D(n4112), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[2]) );
  SDFFR_X1 dscratch1_q_reg_2_ ( .D(n564), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[2]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__2_ ( .D(n4113), .SI(1'b0), .SE(1'b0), 
        .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[2]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__2_ ( .D(n4113), .SI(1'b0), .SE(1'b0), 
        .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[34]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__2_ ( .D(n4113), .SI(1'b0), .SE(1'b0), 
        .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[66]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__2_ ( .D(n4113), .SI(1'b0), .SE(1'b0), 
        .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[98]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__2_ ( .D(n4113), .SI(1'b0), .SE(1'b0), 
        .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[130]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__2_ ( .D(n4113), .SI(1'b0), .SE(1'b0), 
        .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[162]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__2_ ( .D(n4113), .SI(1'b0), .SE(1'b0), 
        .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[194]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__2_ ( .D(n4113), .SI(1'b0), .SE(1'b0), 
        .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[226]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__2_ ( .D(n4113), .SI(1'b0), .SE(1'b0), 
        .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[258]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__2_ ( .D(n4113), .SI(1'b0), .SE(1'b0), 
        .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[290]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__2_ ( .D(n4113), .SI(1'b0), .SE(1'b0), 
        .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[322]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__2_ ( .D(n4113), .SI(1'b0), .SE(1'b0), 
        .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[354]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__2_ ( .D(n4113), .SI(1'b0), .SE(1'b0), 
        .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[386]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__2_ ( .D(n564), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[418]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__2_ ( .D(n564), .SI(1'b0), .SE(1'b0), 
        .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[450]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__2_ ( .D(n564), .SI(1'b0), .SE(1'b0), 
        .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[482]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__0__2_ ( .D(n564), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(pmp_cfg_o[2]), .QN(n1470) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__8__2_ ( .D(n564), .SI(1'b0), .SE(1'b0), .CK(
        n3964), .RN(rst_n), .Q(pmp_cfg_o[66]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__12__2_ ( .D(n564), .SI(1'b0), .SE(1'b0), .CK(
        n3967), .RN(rst_n), .Q(pmp_cfg_o[98]) );
  SDFFR_X1 mcause_q_reg_4_ ( .D(n3928), .SI(1'b0), .SE(1'b0), .CK(n3932), .RN(
        rst_n), .Q(mcause_q[4]) );
  SDFFR_X1 uepc_q_reg_4_ ( .D(uepc_n[4]), .SI(1'b0), .SE(1'b0), .CK(n3999), 
        .RN(rst_n), .Q(uepc_o[4]) );
  SDFFR_X1 depc_q_reg_4_ ( .D(n4010), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[4]) );
  SDFFR_X1 mepc_q_reg_4_ ( .D(n4044), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[4]) );
  SDFFR_X1 ucause_q_reg_4_ ( .D(n3938), .SI(1'b0), .SE(1'b0), .CK(n3942), .RN(
        rst_n), .Q(ucause_q[4]) );
  SDFFR_X1 mstatus_q_reg_upie_ ( .D(n2807), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(rst_n), .Q(mstatus_q[4]) );
  SDFFR_X1 mstatus_q_reg_uie_ ( .D(mstatus_n[4]), .SI(1'b0), .SE(1'b0), .CK(
        clk), .RN(rst_n), .Q(mstatus_q[6]), .QN(n1455) );
  SDFFR_X1 mstatus_q_reg_mpie_ ( .D(mstatus_n[2]), .SI(1'b0), .SE(1'b0), .CK(
        clk), .RN(rst_n), .Q(mstatus_q[3]), .QN(n1461) );
  SDFFR_X1 mstatus_q_reg_mie_ ( .D(mstatus_n[3]), .SI(1'b0), .SE(1'b0), .CK(
        clk), .RN(rst_n), .Q(mstatus_q[5]), .QN(n1454) );
  SDFFR_X1 uepc_q_reg_3_ ( .D(n3979), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[3]) );
  SDFFR_X1 mcause_q_reg_3_ ( .D(n3929), .SI(1'b0), .SE(1'b0), .CK(n3932), .RN(
        rst_n), .Q(mcause_q[3]) );
  SDFFR_X1 depc_q_reg_3_ ( .D(n4011), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[3]) );
  SDFFR_X1 mepc_q_reg_3_ ( .D(n4045), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[3]) );
  SDFFR_X1 ucause_q_reg_3_ ( .D(n3939), .SI(1'b0), .SE(1'b0), .CK(n3942), .RN(
        rst_n), .Q(ucause_q[3]) );
  SDFFR_X1 mscratch_q_reg_3_ ( .D(n4075), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[3]) );
  SDFFR_X1 dscratch0_q_reg_3_ ( .D(n4114), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[3]) );
  SDFFR_X1 dscratch1_q_reg_3_ ( .D(hwlp_data_o[3]), .SI(1'b0), .SE(1'b0), .CK(
        n4101), .RN(rst_n), .Q(dscratch1_q[3]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__3_ ( .D(hwlp_data_o[3]), .SI(1'b0), .SE(
        1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[3]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__3_ ( .D(n4184), .SI(1'b0), .SE(1'b0), 
        .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[35]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__3_ ( .D(hwlp_data_o[3]), .SI(1'b0), .SE(
        1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[67]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__3_ ( .D(n4184), .SI(1'b0), .SE(1'b0), 
        .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[99]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__3_ ( .D(hwlp_data_o[3]), .SI(1'b0), .SE(
        1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[131]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__3_ ( .D(n4184), .SI(1'b0), .SE(1'b0), 
        .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[163]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__3_ ( .D(hwlp_data_o[3]), .SI(1'b0), .SE(
        1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[195]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__3_ ( .D(n4184), .SI(1'b0), .SE(1'b0), 
        .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[227]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__3_ ( .D(hwlp_data_o[3]), .SI(1'b0), .SE(
        1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[259]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__3_ ( .D(n4184), .SI(1'b0), .SE(1'b0), 
        .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[291]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__3_ ( .D(hwlp_data_o[3]), .SI(1'b0), .SE(
        1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[323]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__3_ ( .D(n4184), .SI(1'b0), .SE(1'b0), 
        .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[355]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__3_ ( .D(hwlp_data_o[3]), .SI(1'b0), .SE(
        1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[387]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__3_ ( .D(n4184), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[419]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__3_ ( .D(hwlp_data_o[3]), .SI(1'b0), .SE(
        1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[451]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__3_ ( .D(n4184), .SI(1'b0), .SE(1'b0), 
        .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[483]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__0__3_ ( .D(hwlp_data_o[3]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(pmp_cfg_o[3]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__4__3_ ( .D(n4184), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(pmp_cfg_o[35]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__8__3_ ( .D(hwlp_data_o[3]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[67]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__12__3_ ( .D(n4184), .SI(1'b0), .SE(1'b0), 
        .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[99]) );
  SDFFR_X1 uepc_q_reg_7_ ( .D(n3980), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[7]) );
  SDFFR_X1 depc_q_reg_7_ ( .D(n4012), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[7]) );
  SDFFR_X1 mepc_q_reg_7_ ( .D(n4046), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[7]) );
  SDFFR_X1 dcsr_q_reg_cause__7_ ( .D(n3919), .SI(1'b0), .SE(1'b0), .CK(n3922), 
        .RN(rst_n), .Q(dcsr_q_cause__7_) );
  SDFFR_X1 mscratch_q_reg_7_ ( .D(n4076), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[7]) );
  SDFFR_X1 dscratch0_q_reg_7_ ( .D(n4115), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[7]) );
  SDFFR_X1 dscratch1_q_reg_7_ ( .D(n520), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[7]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__7_ ( .D(n4116), .SI(1'b0), .SE(1'b0), 
        .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[7]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__7_ ( .D(n4116), .SI(1'b0), .SE(1'b0), 
        .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[39]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__7_ ( .D(n4116), .SI(1'b0), .SE(1'b0), 
        .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[71]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__7_ ( .D(n4116), .SI(1'b0), .SE(1'b0), 
        .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[103]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__7_ ( .D(n4116), .SI(1'b0), .SE(1'b0), 
        .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[135]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__7_ ( .D(n4116), .SI(1'b0), .SE(1'b0), 
        .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[167]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__7_ ( .D(n4116), .SI(1'b0), .SE(1'b0), 
        .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[199]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__7_ ( .D(n4116), .SI(1'b0), .SE(1'b0), 
        .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[231]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__7_ ( .D(n4116), .SI(1'b0), .SE(1'b0), 
        .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[263]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__7_ ( .D(n4116), .SI(1'b0), .SE(1'b0), 
        .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[295]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__7_ ( .D(n4116), .SI(1'b0), .SE(1'b0), 
        .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[327]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__7_ ( .D(n4116), .SI(1'b0), .SE(1'b0), 
        .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[359]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__7_ ( .D(n520), .SI(1'b0), .SE(1'b0), 
        .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[391]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__7_ ( .D(n520), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[423]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__7_ ( .D(n520), .SI(1'b0), .SE(1'b0), 
        .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[455]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__7_ ( .D(n520), .SI(1'b0), .SE(1'b0), 
        .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[487]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__0__7_ ( .D(n520), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(n51) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__4__7_ ( .D(n520), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(n39) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__8__7_ ( .D(n520), .SI(1'b0), .SE(1'b0), .CK(
        n3964), .RN(rst_n), .Q(n27) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__12__7_ ( .D(n520), .SI(1'b0), .SE(1'b0), .CK(
        n3967), .RN(rst_n), .Q(n15) );
  SDFFR_X1 uepc_q_reg_0_ ( .D(uepc_n[0]), .SI(1'b0), .SE(1'b0), .CK(n3999), 
        .RN(rst_n), .Q(n4) );
  SDFFR_X1 mcause_q_reg_0_ ( .D(n3930), .SI(1'b0), .SE(1'b0), .CK(n3932), .RN(
        rst_n), .Q(mcause_q[0]) );
  SDFFR_X1 ucause_q_reg_0_ ( .D(n3940), .SI(1'b0), .SE(1'b0), .CK(n3942), .RN(
        rst_n), .Q(ucause_q[0]) );
  SDFFR_X1 mscratch_q_reg_0_ ( .D(n4077), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[0]) );
  SDFFR_X1 dscratch0_q_reg_0_ ( .D(n4117), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[0]) );
  SDFFR_X1 dscratch1_q_reg_0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(1'b0), .CK(
        n4101), .RN(rst_n), .Q(dscratch1_q[0]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[0]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[32]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[64]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[96]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[160]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[192]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[224]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[256]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[288]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[320]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[352]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[384]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[448]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__0__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(pmp_cfg_o[0]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__4__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(pmp_cfg_o[32]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__8__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[64]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__12__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[96]) );
  SDFFR_X1 mscratch_q_reg_4_ ( .D(n4078), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[4]) );
  SDFFR_X1 dscratch0_q_reg_4_ ( .D(n4119), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[4]) );
  SDFFR_X1 dscratch1_q_reg_4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(1'b0), .CK(
        n4101), .RN(rst_n), .Q(dscratch1_q[4]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[4]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[36]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[68]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[100]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[132]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[164]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[196]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[228]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[260]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[292]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[324]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[356]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[388]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[420]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[452]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[484]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__0__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(pmp_cfg_o[4]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__4__4_ ( .D(n2114), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(pmp_cfg_o[36]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__8__4_ ( .D(n2082), .SI(1'b0), .SE(1'b0), .CK(
        n3964), .RN(rst_n), .Q(pmp_cfg_o[68]) );
  SDFFR_X1 uepc_q_reg_11_ ( .D(uepc_n[11]), .SI(1'b0), .SE(1'b0), .CK(n3999), 
        .RN(rst_n), .Q(uepc_o[11]) );
  SDFFR_X1 depc_q_reg_11_ ( .D(n4013), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[11]) );
  SDFFR_X1 dcsr_q_reg_stepie_ ( .D(hwlp_data_o[11]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(dcsr_q_stepie_) );
  SDFFR_X1 mtvec_q_reg_3_ ( .D(hwlp_data_o[11]), .SI(1'b0), .SE(1'b0), .CK(
        n3962), .RN(rst_n), .Q(mtvec_o[3]) );
  SDFFR_X1 mscratch_q_reg_11_ ( .D(n4079), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[11]) );
  SDFFR_X1 dscratch0_q_reg_11_ ( .D(n4120), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[11]) );
  SDFFR_X1 dscratch1_q_reg_11_ ( .D(n2764), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[11]), .QN(n1579) );
  SDFFR_X1 utvec_q_reg_3_ ( .D(hwlp_data_o[11]), .SI(1'b0), .SE(1'b0), .CK(
        n3958), .RN(rst_n), .Q(utvec_o[3]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[11]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[43]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[75]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[107]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[139]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[171]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[203]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[235]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[267]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[299]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[331]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[363]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[395]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[427]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[459]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__11_ ( .D(hwlp_data_o[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[491]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__1__3_ ( .D(hwlp_data_o[11]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(pmp_cfg_o[11]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__9__3_ ( .D(hwlp_data_o[11]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[75]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__13__3_ ( .D(n2041), .SI(1'b0), .SE(1'b0), 
        .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[107]) );
  SDFFR_X1 uepc_q_reg_12_ ( .D(uepc_n[12]), .SI(1'b0), .SE(1'b0), .CK(n3999), 
        .RN(rst_n), .Q(uepc_o[12]) );
  SDFFR_X1 depc_q_reg_12_ ( .D(n4014), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[12]) );
  SDFFR_X1 mepc_q_reg_12_ ( .D(n4048), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[12]) );
  SDFFR_X1 dcsr_q_reg_ebreaku_ ( .D(hwlp_data_o[12]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(debug_ebreaku_o) );
  SDFFR_X1 mtvec_q_reg_4_ ( .D(hwlp_data_o[12]), .SI(1'b0), .SE(1'b0), .CK(
        n3962), .RN(rst_n), .Q(mtvec_o[4]) );
  SDFFR_X1 mscratch_q_reg_12_ ( .D(n2761), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[12]), .QN(n1580) );
  SDFFR_X1 dscratch0_q_reg_12_ ( .D(n4121), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[12]) );
  SDFFR_X1 dscratch1_q_reg_12_ ( .D(hwlp_data_o[12]), .SI(1'b0), .SE(1'b0), 
        .CK(n4101), .RN(rst_n), .Q(dscratch1_q[12]) );
  SDFFR_X1 utvec_q_reg_4_ ( .D(hwlp_data_o[12]), .SI(1'b0), .SE(1'b0), .CK(
        n3958), .RN(rst_n), .Q(utvec_o[4]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[12]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[44]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[76]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[108]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[140]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[172]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[204]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[236]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[268]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[300]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[332]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[364]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[396]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[428]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[460]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__12_ ( .D(hwlp_data_o[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[492]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__1__4_ ( .D(n2138), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(pmp_cfg_o[12]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__5__4_ ( .D(hwlp_data_o[12]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(pmp_cfg_o[44]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__9__4_ ( .D(hwlp_data_o[12]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[76]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__13__4_ ( .D(hwlp_data_o[12]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[108]) );
  SDFFR_X1 PCCR_q_reg_0__13_ ( .D(PCCR_n[12]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[13]), .QN(n1487) );
  SDFFR_X1 uepc_q_reg_13_ ( .D(n3981), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[13]) );
  SDFFR_X1 depc_q_reg_13_ ( .D(n4015), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[13]) );
  SDFFR_X1 mepc_q_reg_13_ ( .D(n4049), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[13]) );
  SDFFR_X1 dcsr_q_reg_ebreaks_ ( .D(n3960), .SI(1'b0), .SE(1'b0), .CK(n3946), 
        .RN(rst_n), .Q(dcsr_q_ebreaks_) );
  SDFFR_X1 mtvec_q_reg_5_ ( .D(n3960), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[5]) );
  SDFFR_X1 mscratch_q_reg_13_ ( .D(n4080), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[13]) );
  SDFFR_X1 dscratch0_q_reg_13_ ( .D(n4122), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[13]) );
  SDFFR_X1 dscratch1_q_reg_13_ ( .D(n3960), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[13]) );
  SDFFR_X1 utvec_q_reg_5_ ( .D(n3960), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[5]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__13_ ( .D(n3960), .SI(1'b0), .SE(1'b0), 
        .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[13]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__13_ ( .D(n501), .SI(1'b0), .SE(1'b0), 
        .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[45]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__13_ ( .D(n501), .SI(1'b0), .SE(1'b0), 
        .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[77]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__13_ ( .D(n501), .SI(1'b0), .SE(1'b0), 
        .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[109]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__13_ ( .D(n501), .SI(1'b0), .SE(1'b0), 
        .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[141]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__13_ ( .D(n501), .SI(1'b0), .SE(1'b0), 
        .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[173]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__13_ ( .D(n501), .SI(1'b0), .SE(1'b0), 
        .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[205]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__13_ ( .D(n501), .SI(1'b0), .SE(1'b0), 
        .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[237]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__13_ ( .D(n501), .SI(1'b0), .SE(1'b0), 
        .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[269]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__13_ ( .D(n501), .SI(1'b0), .SE(1'b0), 
        .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[301]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__13_ ( .D(n3960), .SI(1'b0), .SE(1'b0), 
        .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[333]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__13_ ( .D(n3960), .SI(1'b0), .SE(1'b0), 
        .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[365]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__13_ ( .D(n3960), .SI(1'b0), .SE(1'b0), 
        .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[397]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__13_ ( .D(n3960), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[429]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__13_ ( .D(n3960), .SI(1'b0), .SE(1'b0), 
        .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[461]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__13_ ( .D(n3960), .SI(1'b0), .SE(1'b0), 
        .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[493]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__1__5_ ( .D(n3960), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(n50) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__5__5_ ( .D(n3960), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(n38) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__9__5_ ( .D(n3960), .SI(1'b0), .SE(1'b0), .CK(
        n3964), .RN(rst_n), .Q(n26) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__13__5_ ( .D(n3960), .SI(1'b0), .SE(1'b0), 
        .CK(n3967), .RN(rst_n), .Q(n14) );
  SDFFR_X1 PCCR_q_reg_0__14_ ( .D(PCCR_n[13]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[14]), .QN(n1483) );
  SDFFR_X1 uepc_q_reg_14_ ( .D(n3982), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[14]) );
  SDFFR_X1 depc_q_reg_14_ ( .D(n4016), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[14]) );
  SDFFR_X1 mepc_q_reg_14_ ( .D(n4050), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[14]) );
  SDFFR_X1 dcsr_q_reg_zero1_ ( .D(hwlp_data_o[14]), .SI(1'b0), .SE(1'b0), .CK(
        n3946), .RN(rst_n), .Q(dcsr_q_zero1_) );
  SDFFR_X1 mtvec_q_reg_6_ ( .D(hwlp_data_o[14]), .SI(1'b0), .SE(1'b0), .CK(
        n3962), .RN(rst_n), .Q(mtvec_o[6]) );
  SDFFR_X1 mscratch_q_reg_14_ ( .D(n4081), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[14]) );
  SDFFR_X1 dscratch0_q_reg_14_ ( .D(n4123), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[14]) );
  SDFFR_X1 dscratch1_q_reg_14_ ( .D(hwlp_data_o[14]), .SI(1'b0), .SE(1'b0), 
        .CK(n4101), .RN(rst_n), .Q(dscratch1_q[14]) );
  SDFFR_X1 utvec_q_reg_6_ ( .D(hwlp_data_o[14]), .SI(1'b0), .SE(1'b0), .CK(
        n3958), .RN(rst_n), .Q(utvec_o[6]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__14_ ( .D(hwlp_data_o[14]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[14]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__14_ ( .D(hwlp_data_o[14]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[46]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__14_ ( .D(hwlp_data_o[14]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[78]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__14_ ( .D(hwlp_data_o[14]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[110]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__14_ ( .D(hwlp_data_o[14]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[142]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__14_ ( .D(hwlp_data_o[14]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[174]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__14_ ( .D(n443), .SI(1'b0), .SE(1'b0), 
        .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[206]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__14_ ( .D(n443), .SI(1'b0), .SE(1'b0), 
        .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[238]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__14_ ( .D(n443), .SI(1'b0), .SE(1'b0), 
        .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[270]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__14_ ( .D(n443), .SI(1'b0), .SE(1'b0), 
        .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[302]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__14_ ( .D(n443), .SI(1'b0), .SE(1'b0), 
        .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[334]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__14_ ( .D(n443), .SI(1'b0), .SE(1'b0), 
        .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[366]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__14_ ( .D(n443), .SI(1'b0), .SE(1'b0), 
        .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[398]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__14_ ( .D(n443), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[430]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__14_ ( .D(n443), .SI(1'b0), .SE(1'b0), 
        .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[462]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__14_ ( .D(n443), .SI(1'b0), .SE(1'b0), 
        .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[494]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__1__6_ ( .D(n443), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(n49) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__5__6_ ( .D(n443), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(n37) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__9__6_ ( .D(hwlp_data_o[14]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(n25) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__13__6_ ( .D(hwlp_data_o[14]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(n13) );
  SDFFR_X1 PCCR_q_reg_0__15_ ( .D(PCCR_n[14]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[15]), .QN(n1484) );
  SDFFR_X1 uepc_q_reg_15_ ( .D(n3983), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[15]) );
  SDFFR_X1 depc_q_reg_15_ ( .D(n4017), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[15]) );
  SDFFR_X1 mepc_q_reg_15_ ( .D(n4051), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[15]) );
  SDFFR_X1 dcsr_q_reg_ebreakm_ ( .D(hwlp_data_o[15]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(debug_ebreakm_o) );
  SDFFR_X1 mtvec_q_reg_7_ ( .D(hwlp_data_o[15]), .SI(1'b0), .SE(1'b0), .CK(
        n3962), .RN(rst_n), .Q(mtvec_o[7]) );
  SDFFR_X1 mscratch_q_reg_15_ ( .D(n4082), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[15]) );
  SDFFR_X1 dscratch0_q_reg_15_ ( .D(n4125), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[15]) );
  SDFFR_X1 dscratch1_q_reg_15_ ( .D(hwlp_data_o[15]), .SI(1'b0), .SE(1'b0), 
        .CK(n4101), .RN(rst_n), .Q(dscratch1_q[15]) );
  SDFFR_X1 utvec_q_reg_7_ ( .D(hwlp_data_o[15]), .SI(1'b0), .SE(1'b0), .CK(
        n3958), .RN(rst_n), .Q(utvec_o[7]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__15_ ( .D(hwlp_data_o[15]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[15]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__15_ ( .D(hwlp_data_o[15]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[47]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__15_ ( .D(hwlp_data_o[15]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[79]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__15_ ( .D(hwlp_data_o[15]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[111]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__15_ ( .D(n543), .SI(1'b0), .SE(1'b0), 
        .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[143]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__15_ ( .D(n543), .SI(1'b0), .SE(1'b0), 
        .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[175]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__15_ ( .D(n543), .SI(1'b0), .SE(1'b0), 
        .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[207]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__15_ ( .D(n543), .SI(1'b0), .SE(1'b0), 
        .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[239]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__15_ ( .D(n543), .SI(1'b0), .SE(1'b0), 
        .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[271]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__15_ ( .D(n543), .SI(1'b0), .SE(1'b0), 
        .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[303]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__15_ ( .D(n543), .SI(1'b0), .SE(1'b0), 
        .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[335]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__15_ ( .D(n543), .SI(1'b0), .SE(1'b0), 
        .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[367]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__15_ ( .D(n543), .SI(1'b0), .SE(1'b0), 
        .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[399]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__15_ ( .D(n543), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[431]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__15_ ( .D(n543), .SI(1'b0), .SE(1'b0), 
        .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[463]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__15_ ( .D(n543), .SI(1'b0), .SE(1'b0), 
        .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[495]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__1__7_ ( .D(hwlp_data_o[15]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(n48) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__5__7_ ( .D(hwlp_data_o[15]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(n36) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__9__7_ ( .D(hwlp_data_o[15]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(n24) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__13__7_ ( .D(hwlp_data_o[15]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(n12) );
  SDFFR_X1 PCCR_q_reg_0__16_ ( .D(PCCR_n[15]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[16]), .QN(n1488) );
  SDFFR_X1 uepc_q_reg_16_ ( .D(uepc_n[16]), .SI(1'b0), .SE(1'b0), .CK(n3999), 
        .RN(rst_n), .Q(uepc_o[16]) );
  SDFFR_X1 depc_q_reg_16_ ( .D(depc_n[16]), .SI(1'b0), .SE(1'b0), .CK(n4031), 
        .RN(rst_n), .Q(depc_o[16]) );
  SDFFR_X1 mepc_q_reg_16_ ( .D(mepc_n[16]), .SI(1'b0), .SE(1'b0), .CK(n4065), 
        .RN(rst_n), .Q(mepc_o[16]) );
  SDFFR_X1 dcsr_q_reg_zero2__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(dcsr_q_zero2__16_) );
  SDFFR_X1 mtvec_q_reg_8_ ( .D(hwlp_data_o[16]), .SI(1'b0), .SE(1'b0), .CK(
        n3962), .RN(rst_n), .Q(mtvec_o[8]) );
  SDFFR_X1 mscratch_q_reg_16_ ( .D(n2741), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[16]), .QN(n1622) );
  SDFFR_X1 dscratch0_q_reg_16_ ( .D(n4127), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[16]) );
  SDFFR_X1 dscratch1_q_reg_16_ ( .D(hwlp_data_o[16]), .SI(1'b0), .SE(1'b0), 
        .CK(n4101), .RN(rst_n), .Q(dscratch1_q[16]) );
  SDFFR_X1 utvec_q_reg_8_ ( .D(hwlp_data_o[16]), .SI(1'b0), .SE(1'b0), .CK(
        n3958), .RN(rst_n), .Q(utvec_o[8]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[16]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[48]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[80]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[112]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[144]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[176]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[208]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[240]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[272]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[304]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[336]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[368]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[400]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[432]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[464]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__16_ ( .D(hwlp_data_o[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[496]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__2__0_ ( .D(hwlp_data_o[16]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(pmp_cfg_o[16]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__6__0_ ( .D(hwlp_data_o[16]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(pmp_cfg_o[48]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__10__0_ ( .D(hwlp_data_o[16]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[80]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__14__0_ ( .D(hwlp_data_o[16]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[112]) );
  SDFFR_X1 PCCR_q_reg_0__17_ ( .D(PCCR_n[16]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[17]), .QN(n1494) );
  SDFFR_X1 uepc_q_reg_17_ ( .D(n3984), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[17]) );
  SDFFR_X1 depc_q_reg_17_ ( .D(depc_n[17]), .SI(1'b0), .SE(1'b0), .CK(n4031), 
        .RN(rst_n), .Q(depc_o[17]) );
  SDFFR_X1 mepc_q_reg_17_ ( .D(mepc_n[17]), .SI(1'b0), .SE(1'b0), .CK(n4065), 
        .RN(rst_n), .Q(mepc_o[17]) );
  SDFFR_X1 dcsr_q_reg_zero2__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(dcsr_q_zero2__17_) );
  SDFFR_X1 mstatus_q_reg_mprv_ ( .D(N2756), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .RN(rst_n), .Q(mstatus_q[0]) );
  SDFFR_X1 mtvec_q_reg_9_ ( .D(n2737), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[9]), .QN(n1520) );
  SDFFR_X1 mscratch_q_reg_17_ ( .D(n4083), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[17]) );
  SDFFR_X1 dscratch0_q_reg_17_ ( .D(n4128), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[17]) );
  SDFFR_X1 dscratch1_q_reg_17_ ( .D(hwlp_data_o[17]), .SI(1'b0), .SE(1'b0), 
        .CK(n4101), .RN(rst_n), .Q(dscratch1_q[17]) );
  SDFFR_X1 utvec_q_reg_9_ ( .D(n2733), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[9]), .QN(n1544) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[17]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[49]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[81]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[113]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[145]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[177]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[209]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[241]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[273]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[305]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[337]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[369]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[401]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[433]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[465]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__17_ ( .D(hwlp_data_o[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[497]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__2__1_ ( .D(hwlp_data_o[17]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(pmp_cfg_o[17]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__6__1_ ( .D(hwlp_data_o[17]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(pmp_cfg_o[49]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__10__1_ ( .D(hwlp_data_o[17]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[81]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__14__1_ ( .D(hwlp_data_o[17]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[113]) );
  SDFFR_X1 PCCR_q_reg_0__18_ ( .D(PCCR_n[17]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[18]), .QN(n1489) );
  SDFFR_X1 uepc_q_reg_18_ ( .D(n3985), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[18]) );
  SDFFR_X1 depc_q_reg_18_ ( .D(n4018), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[18]) );
  SDFFR_X1 mepc_q_reg_18_ ( .D(n4052), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[18]) );
  SDFFR_X1 dcsr_q_reg_zero2__18_ ( .D(hwlp_data_o[18]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(dcsr_q_zero2__18_) );
  SDFFR_X1 mtvec_q_reg_10_ ( .D(hwlp_data_o[18]), .SI(1'b0), .SE(1'b0), .CK(
        n3962), .RN(rst_n), .Q(mtvec_o[10]) );
  SDFFR_X1 mscratch_q_reg_18_ ( .D(n4084), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[18]) );
  SDFFR_X1 dscratch0_q_reg_18_ ( .D(n4130), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[18]) );
  SDFFR_X1 dscratch1_q_reg_18_ ( .D(hwlp_data_o[18]), .SI(1'b0), .SE(1'b0), 
        .CK(n4101), .RN(rst_n), .Q(dscratch1_q[18]) );
  SDFFR_X1 utvec_q_reg_10_ ( .D(hwlp_data_o[18]), .SI(1'b0), .SE(1'b0), .CK(
        n3958), .RN(rst_n), .Q(utvec_o[10]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__18_ ( .D(hwlp_data_o[18]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[18]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__18_ ( .D(hwlp_data_o[18]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[50]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__18_ ( .D(hwlp_data_o[18]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[82]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__18_ ( .D(hwlp_data_o[18]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[114]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__18_ ( .D(hwlp_data_o[18]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[146]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__18_ ( .D(hwlp_data_o[18]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[178]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__18_ ( .D(n1675), .SI(1'b0), .SE(1'b0), 
        .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[210]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__18_ ( .D(n1675), .SI(1'b0), .SE(1'b0), 
        .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[242]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__18_ ( .D(n1675), .SI(1'b0), .SE(1'b0), 
        .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[274]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__18_ ( .D(n1675), .SI(1'b0), .SE(1'b0), 
        .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[306]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__18_ ( .D(n1675), .SI(1'b0), .SE(1'b0), 
        .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[338]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__18_ ( .D(n1675), .SI(1'b0), .SE(1'b0), 
        .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[370]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__18_ ( .D(n1675), .SI(1'b0), .SE(1'b0), 
        .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[402]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__18_ ( .D(n1675), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[434]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__18_ ( .D(n1675), .SI(1'b0), .SE(1'b0), 
        .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[466]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__18_ ( .D(n1675), .SI(1'b0), .SE(1'b0), 
        .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[498]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__2__2_ ( .D(n1675), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(pmp_cfg_o[18]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__6__2_ ( .D(n1675), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(pmp_cfg_o[50]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__10__2_ ( .D(hwlp_data_o[18]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[82]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__14__2_ ( .D(hwlp_data_o[18]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[114]) );
  SDFFR_X1 PCCR_q_reg_0__19_ ( .D(PCCR_n[18]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[19]), .QN(n1495) );
  SDFFR_X1 uepc_q_reg_19_ ( .D(n3986), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[19]) );
  SDFFR_X1 depc_q_reg_19_ ( .D(n4019), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[19]) );
  SDFFR_X1 mepc_q_reg_19_ ( .D(n4053), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[19]) );
  SDFFR_X1 dcsr_q_reg_zero2__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(dcsr_q_zero2__19_) );
  SDFFR_X1 mtvec_q_reg_11_ ( .D(n3951), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[11]) );
  SDFFR_X1 mscratch_q_reg_19_ ( .D(n4085), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[19]) );
  SDFFR_X1 dscratch0_q_reg_19_ ( .D(n4132), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[19]) );
  SDFFR_X1 dscratch1_q_reg_19_ ( .D(n3951), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[19]) );
  SDFFR_X1 utvec_q_reg_11_ ( .D(n3951), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[11]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[19]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[51]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[83]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[115]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[147]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[179]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[211]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[243]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[275]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[307]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[339]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[371]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[403]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[435]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[467]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__19_ ( .D(hwlp_data_o[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[499]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__2__3_ ( .D(n2129), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(pmp_cfg_o[19]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__6__3_ ( .D(n2097), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(pmp_cfg_o[51]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__10__3_ ( .D(n2065), .SI(1'b0), .SE(1'b0), 
        .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[83]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__14__3_ ( .D(n2033), .SI(1'b0), .SE(1'b0), 
        .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[115]) );
  SDFFR_X1 PCCR_q_reg_0__20_ ( .D(PCCR_n[19]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[20]), .QN(n1464) );
  SDFFR_X1 uepc_q_reg_20_ ( .D(n3987), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[20]) );
  SDFFR_X1 depc_q_reg_20_ ( .D(n4020), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[20]) );
  SDFFR_X1 mepc_q_reg_20_ ( .D(n4054), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[20]) );
  SDFFR_X1 dcsr_q_reg_zero2__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(dcsr_q_zero2__20_) );
  SDFFR_X1 mtvec_q_reg_12_ ( .D(n1678), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[12]) );
  SDFFR_X1 mscratch_q_reg_20_ ( .D(n4086), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[20]) );
  SDFFR_X1 dscratch0_q_reg_20_ ( .D(n4133), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[20]) );
  SDFFR_X1 dscratch1_q_reg_20_ ( .D(n1678), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[20]) );
  SDFFR_X1 utvec_q_reg_12_ ( .D(n1678), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[12]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[20]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[52]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[84]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[116]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[148]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[180]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[212]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[244]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[276]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[308]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[340]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[372]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[404]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[436]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[468]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__20_ ( .D(hwlp_data_o[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[500]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__2__4_ ( .D(hwlp_data_o[20]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(pmp_cfg_o[20]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__6__4_ ( .D(n2098), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(pmp_cfg_o[52]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__14__4_ ( .D(n2034), .SI(1'b0), .SE(1'b0), 
        .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[116]) );
  SDFFR_X1 PCCR_q_reg_0__21_ ( .D(PCCR_n[20]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[21]), .QN(n1485) );
  SDFFR_X1 uepc_q_reg_21_ ( .D(n3988), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[21]) );
  SDFFR_X1 depc_q_reg_21_ ( .D(n4021), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[21]) );
  SDFFR_X1 mepc_q_reg_21_ ( .D(n4055), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[21]) );
  SDFFR_X1 dcsr_q_reg_zero2__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(dcsr_q_zero2__21_) );
  SDFFR_X1 mtvec_q_reg_13_ ( .D(n4183), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[13]) );
  SDFFR_X1 mscratch_q_reg_21_ ( .D(n4087), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[21]) );
  SDFFR_X1 dscratch0_q_reg_21_ ( .D(n4134), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[21]) );
  SDFFR_X1 dscratch1_q_reg_21_ ( .D(n4183), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[21]) );
  SDFFR_X1 utvec_q_reg_13_ ( .D(hwlp_data_o[21]), .SI(1'b0), .SE(1'b0), .CK(
        n3958), .RN(rst_n), .Q(utvec_o[13]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[21]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[53]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[85]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[117]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[149]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[181]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[245]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[277]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[309]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[341]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[373]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[405]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[437]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[469]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[501]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__2__5_ ( .D(hwlp_data_o[21]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(n47) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__6__5_ ( .D(n2099), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(n35) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__10__5_ ( .D(hwlp_data_o[21]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(n23) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__14__5_ ( .D(n2035), .SI(1'b0), .SE(1'b0), 
        .CK(n3967), .RN(rst_n), .Q(n11) );
  SDFFR_X1 PCCR_q_reg_0__22_ ( .D(PCCR_n[21]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[22]), .QN(n1502) );
  SDFFR_X1 uepc_q_reg_22_ ( .D(n3989), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[22]) );
  SDFFR_X1 depc_q_reg_22_ ( .D(n4022), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[22]) );
  SDFFR_X1 mepc_q_reg_22_ ( .D(n4056), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[22]) );
  SDFFR_X1 dcsr_q_reg_zero2__22_ ( .D(hwlp_data_o[22]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(dcsr_q_zero2__22_) );
  SDFFR_X1 mtvec_q_reg_14_ ( .D(hwlp_data_o[22]), .SI(1'b0), .SE(1'b0), .CK(
        n3962), .RN(rst_n), .Q(mtvec_o[14]) );
  SDFFR_X1 mscratch_q_reg_22_ ( .D(n4088), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[22]) );
  SDFFR_X1 dscratch0_q_reg_22_ ( .D(n4135), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[22]) );
  SDFFR_X1 dscratch1_q_reg_22_ ( .D(hwlp_data_o[22]), .SI(1'b0), .SE(1'b0), 
        .CK(n4101), .RN(rst_n), .Q(dscratch1_q[22]) );
  SDFFR_X1 utvec_q_reg_14_ ( .D(hwlp_data_o[22]), .SI(1'b0), .SE(1'b0), .CK(
        n3958), .RN(rst_n), .Q(utvec_o[14]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__22_ ( .D(hwlp_data_o[22]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[22]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__22_ ( .D(n1007), .SI(1'b0), .SE(1'b0), 
        .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[54]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__22_ ( .D(n1007), .SI(1'b0), .SE(1'b0), 
        .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[86]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__22_ ( .D(hwlp_data_o[22]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[118]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__22_ ( .D(hwlp_data_o[22]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[150]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__22_ ( .D(n1007), .SI(1'b0), .SE(1'b0), 
        .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[182]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__22_ ( .D(n1007), .SI(1'b0), .SE(1'b0), 
        .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[214]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__22_ ( .D(hwlp_data_o[22]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[246]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__22_ ( .D(hwlp_data_o[22]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[278]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__22_ ( .D(n1007), .SI(1'b0), .SE(1'b0), 
        .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[310]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__22_ ( .D(n1007), .SI(1'b0), .SE(1'b0), 
        .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[342]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__22_ ( .D(hwlp_data_o[22]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[374]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__22_ ( .D(hwlp_data_o[22]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[406]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__22_ ( .D(n1007), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[438]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__22_ ( .D(n1007), .SI(1'b0), .SE(1'b0), 
        .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[470]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__22_ ( .D(hwlp_data_o[22]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[502]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__2__6_ ( .D(hwlp_data_o[22]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(n46) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__6__6_ ( .D(hwlp_data_o[22]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(n34) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__10__6_ ( .D(n2068), .SI(1'b0), .SE(1'b0), 
        .CK(n3964), .RN(rst_n), .Q(n22) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__14__6_ ( .D(n1007), .SI(1'b0), .SE(1'b0), 
        .CK(n3967), .RN(rst_n), .Q(n10) );
  SDFFR_X1 PCCR_q_reg_0__23_ ( .D(PCCR_n[22]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[23]), .QN(n1465) );
  SDFFR_X1 uepc_q_reg_23_ ( .D(n3990), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[23]) );
  SDFFR_X1 depc_q_reg_23_ ( .D(n4023), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[23]) );
  SDFFR_X1 mepc_q_reg_23_ ( .D(n4057), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[23]) );
  SDFFR_X1 dcsr_q_reg_zero2__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(dcsr_q_zero2__23_) );
  SDFFR_X1 mtvec_q_reg_15_ ( .D(n3952), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[15]) );
  SDFFR_X1 mscratch_q_reg_23_ ( .D(n4089), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[23]) );
  SDFFR_X1 dscratch0_q_reg_23_ ( .D(n4136), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[23]) );
  SDFFR_X1 dscratch1_q_reg_23_ ( .D(n3952), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[23]) );
  SDFFR_X1 utvec_q_reg_15_ ( .D(n3952), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[15]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[23]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[55]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[87]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[119]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[151]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[183]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[215]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[247]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[279]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[311]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[343]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[375]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[407]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[439]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[471]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__23_ ( .D(hwlp_data_o[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[503]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__2__7_ ( .D(hwlp_data_o[23]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(n45) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__6__7_ ( .D(hwlp_data_o[23]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(n33) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__10__7_ ( .D(hwlp_data_o[23]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(n21) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__14__7_ ( .D(hwlp_data_o[23]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(n9) );
  SDFFR_X1 PCCR_q_reg_0__24_ ( .D(PCCR_n[23]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[24]), .QN(n1486) );
  SDFFR_X1 uepc_q_reg_24_ ( .D(n3991), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[24]) );
  SDFFR_X1 depc_q_reg_24_ ( .D(n4024), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[24]) );
  SDFFR_X1 mepc_q_reg_24_ ( .D(mepc_n[24]), .SI(1'b0), .SE(1'b0), .CK(n4065), 
        .RN(rst_n), .Q(mepc_o[24]) );
  SDFFR_X1 dcsr_q_reg_zero2__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(dcsr_q_zero2__24_) );
  SDFFR_X1 mtvec_q_reg_16_ ( .D(n3953), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[16]) );
  SDFFR_X1 mscratch_q_reg_24_ ( .D(n4090), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[24]) );
  SDFFR_X1 dscratch0_q_reg_24_ ( .D(n4137), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[24]) );
  SDFFR_X1 dscratch1_q_reg_24_ ( .D(n3953), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[24]) );
  SDFFR_X1 utvec_q_reg_16_ ( .D(n3953), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[16]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[24]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[56]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[88]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[120]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[152]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[184]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[216]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[248]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[280]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[312]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[344]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[376]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[408]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[440]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[472]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__24_ ( .D(hwlp_data_o[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[504]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__3__0_ ( .D(n2126), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(pmp_cfg_o[24]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__7__0_ ( .D(n2094), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(pmp_cfg_o[56]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__11__0_ ( .D(n2062), .SI(1'b0), .SE(1'b0), 
        .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[88]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__15__0_ ( .D(hwlp_data_o[24]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[120]) );
  SDFFR_X1 PCCR_q_reg_0__25_ ( .D(PCCR_n[24]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[25]), .QN(n1496) );
  SDFFR_X1 uepc_q_reg_25_ ( .D(n3992), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[25]) );
  SDFFR_X1 depc_q_reg_25_ ( .D(n4025), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[25]) );
  SDFFR_X1 mepc_q_reg_25_ ( .D(n4058), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[25]) );
  SDFFR_X1 dcsr_q_reg_zero2__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(dcsr_q_zero2__25_) );
  SDFFR_X1 mtvec_q_reg_17_ ( .D(n3954), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[17]) );
  SDFFR_X1 mscratch_q_reg_25_ ( .D(n4091), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[25]) );
  SDFFR_X1 dscratch0_q_reg_25_ ( .D(n4138), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[25]) );
  SDFFR_X1 dscratch1_q_reg_25_ ( .D(n3954), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[25]) );
  SDFFR_X1 utvec_q_reg_17_ ( .D(n3954), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[17]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[25]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[57]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[89]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[121]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[153]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[185]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[217]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[249]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[281]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[313]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[345]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[377]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[409]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[441]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[473]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__25_ ( .D(hwlp_data_o[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[505]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__3__1_ ( .D(hwlp_data_o[25]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(pmp_cfg_o[25]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__7__1_ ( .D(hwlp_data_o[25]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(pmp_cfg_o[57]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__11__1_ ( .D(hwlp_data_o[25]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[89]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__15__1_ ( .D(hwlp_data_o[25]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[121]) );
  SDFFR_X1 PCCR_q_reg_0__26_ ( .D(PCCR_n[25]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[26]), .QN(n1490) );
  SDFFR_X1 uepc_q_reg_26_ ( .D(n3993), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[26]) );
  SDFFR_X1 depc_q_reg_26_ ( .D(n4026), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[26]) );
  SDFFR_X1 mepc_q_reg_26_ ( .D(n4059), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[26]) );
  SDFFR_X1 dcsr_q_reg_zero2__26_ ( .D(n3955), .SI(1'b0), .SE(1'b0), .CK(n3946), 
        .RN(rst_n), .Q(dcsr_q_zero2__26_) );
  SDFFR_X1 mtvec_q_reg_18_ ( .D(n3955), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[18]) );
  SDFFR_X1 mscratch_q_reg_26_ ( .D(n4092), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[26]) );
  SDFFR_X1 dscratch0_q_reg_26_ ( .D(n4139), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[26]) );
  SDFFR_X1 dscratch1_q_reg_26_ ( .D(n3955), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[26]) );
  SDFFR_X1 utvec_q_reg_18_ ( .D(n3955), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[18]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__26_ ( .D(n3955), .SI(1'b0), .SE(1'b0), 
        .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[26]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__26_ ( .D(n3955), .SI(1'b0), .SE(1'b0), 
        .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[58]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__26_ ( .D(n3955), .SI(1'b0), .SE(1'b0), 
        .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[90]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__26_ ( .D(hwlp_data_o[26]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[122]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__26_ ( .D(hwlp_data_o[26]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[154]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__26_ ( .D(hwlp_data_o[26]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[186]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__26_ ( .D(hwlp_data_o[26]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[218]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__26_ ( .D(hwlp_data_o[26]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[250]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__26_ ( .D(hwlp_data_o[26]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[282]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__26_ ( .D(hwlp_data_o[26]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[314]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__26_ ( .D(hwlp_data_o[26]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[346]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__26_ ( .D(hwlp_data_o[26]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[378]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__26_ ( .D(n3955), .SI(1'b0), .SE(1'b0), 
        .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[410]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__26_ ( .D(n3955), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[442]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__26_ ( .D(n3955), .SI(1'b0), .SE(1'b0), 
        .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[474]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__26_ ( .D(n3955), .SI(1'b0), .SE(1'b0), 
        .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[506]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__3__2_ ( .D(n2120), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(pmp_cfg_o[26]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__7__2_ ( .D(n2088), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(pmp_cfg_o[58]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__11__2_ ( .D(n2056), .SI(1'b0), .SE(1'b0), 
        .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[90]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__15__2_ ( .D(n2024), .SI(1'b0), .SE(1'b0), 
        .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[122]) );
  SDFFR_X1 PCCR_q_reg_0__27_ ( .D(PCCR_n[26]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[27]), .QN(n1503) );
  SDFFR_X1 uepc_q_reg_27_ ( .D(n3994), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[27]) );
  SDFFR_X1 depc_q_reg_27_ ( .D(n4027), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[27]) );
  SDFFR_X1 mepc_q_reg_27_ ( .D(n4060), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[27]) );
  SDFFR_X1 dcsr_q_reg_zero2__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), .SE(1'b0), 
        .CK(n3946), .RN(rst_n), .Q(dcsr_q_zero2__27_) );
  SDFFR_X1 mtvec_q_reg_19_ ( .D(n3956), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[19]) );
  SDFFR_X1 mscratch_q_reg_27_ ( .D(n4093), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[27]) );
  SDFFR_X1 dscratch0_q_reg_27_ ( .D(n4140), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[27]) );
  SDFFR_X1 dscratch1_q_reg_27_ ( .D(n3956), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[27]) );
  SDFFR_X1 utvec_q_reg_19_ ( .D(n3956), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[19]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[27]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[59]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[91]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[123]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[155]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[187]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[219]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[251]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[283]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[315]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[347]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[379]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[411]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[443]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[475]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__27_ ( .D(hwlp_data_o[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[507]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__3__3_ ( .D(n2121), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(pmp_cfg_o[27]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__7__3_ ( .D(n2089), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(pmp_cfg_o[59]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__11__3_ ( .D(n2057), .SI(1'b0), .SE(1'b0), 
        .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[91]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__15__3_ ( .D(n2025), .SI(1'b0), .SE(1'b0), 
        .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[123]) );
  SDFFR_X1 uepc_q_reg_28_ ( .D(n3995), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[28]) );
  SDFFR_X1 depc_q_reg_28_ ( .D(n4028), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[28]) );
  SDFFR_X1 mepc_q_reg_28_ ( .D(n4061), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[28]) );
  SDFFR_X1 mtvec_q_reg_20_ ( .D(n3957), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[20]) );
  SDFFR_X1 mscratch_q_reg_28_ ( .D(n4094), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[28]) );
  SDFFR_X1 dscratch0_q_reg_28_ ( .D(n4141), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[28]) );
  SDFFR_X1 dscratch1_q_reg_28_ ( .D(n3957), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[28]) );
  SDFFR_X1 utvec_q_reg_20_ ( .D(n3957), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[20]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[28]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[60]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[92]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[124]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[156]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[188]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[220]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[252]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[284]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[316]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[348]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[380]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[412]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[444]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[476]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__28_ ( .D(hwlp_data_o[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[508]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__3__4_ ( .D(n2122), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(pmp_cfg_o[28]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__7__4_ ( .D(n2090), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(pmp_cfg_o[60]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__11__4_ ( .D(n2058), .SI(1'b0), .SE(1'b0), 
        .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[92]) );
  SDFFR_X1 uepc_q_reg_29_ ( .D(n3996), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[29]) );
  SDFFR_X1 depc_q_reg_29_ ( .D(n4029), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[29]) );
  SDFFR_X1 mepc_q_reg_29_ ( .D(n4062), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[29]) );
  SDFFR_X1 mtvec_q_reg_21_ ( .D(n4143), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[21]) );
  SDFFR_X1 mscratch_q_reg_29_ ( .D(n4095), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[29]) );
  SDFFR_X1 dscratch0_q_reg_29_ ( .D(n4142), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[29]) );
  SDFFR_X1 dscratch1_q_reg_29_ ( .D(n4143), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[29]) );
  SDFFR_X1 utvec_q_reg_21_ ( .D(n4143), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[21]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__29_ ( .D(n4143), .SI(1'b0), .SE(1'b0), 
        .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[29]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__29_ ( .D(n929), .SI(1'b0), .SE(1'b0), 
        .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[61]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__29_ ( .D(n929), .SI(1'b0), .SE(1'b0), 
        .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[93]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__29_ ( .D(n4143), .SI(1'b0), .SE(1'b0), 
        .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[125]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__29_ ( .D(n4143), .SI(1'b0), .SE(1'b0), 
        .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[157]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__29_ ( .D(n4143), .SI(1'b0), .SE(1'b0), 
        .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[189]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__29_ ( .D(n4143), .SI(1'b0), .SE(1'b0), 
        .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[221]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__29_ ( .D(n4143), .SI(1'b0), .SE(1'b0), 
        .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[253]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__29_ ( .D(n4143), .SI(1'b0), .SE(1'b0), 
        .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[285]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__29_ ( .D(n4143), .SI(1'b0), .SE(1'b0), 
        .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[317]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__29_ ( .D(n4143), .SI(1'b0), .SE(1'b0), 
        .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[349]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__29_ ( .D(n4143), .SI(1'b0), .SE(1'b0), 
        .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[381]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__29_ ( .D(n929), .SI(1'b0), .SE(1'b0), 
        .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[413]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__29_ ( .D(n929), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[445]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__29_ ( .D(n929), .SI(1'b0), .SE(1'b0), 
        .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[477]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__29_ ( .D(n929), .SI(1'b0), .SE(1'b0), 
        .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[509]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__3__5_ ( .D(n4143), .SI(1'b0), .SE(1'b0), .CK(
        n3970), .RN(rst_n), .Q(n44) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__7__5_ ( .D(n929), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(n32) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__11__5_ ( .D(n929), .SI(1'b0), .SE(1'b0), .CK(
        n3964), .RN(rst_n), .Q(n20) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__15__5_ ( .D(n929), .SI(1'b0), .SE(1'b0), .CK(
        n3967), .RN(rst_n), .Q(n8) );
  SDFFR_X1 uepc_q_reg_30_ ( .D(n3997), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[30]) );
  SDFFR_X1 depc_q_reg_30_ ( .D(depc_n[30]), .SI(1'b0), .SE(1'b0), .CK(n4031), 
        .RN(rst_n), .Q(depc_o[30]) );
  SDFFR_X1 mepc_q_reg_30_ ( .D(n4063), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[30]) );
  SDFFR_X1 mtvec_q_reg_22_ ( .D(n931), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[22]) );
  SDFFR_X1 mscratch_q_reg_30_ ( .D(n4096), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[30]) );
  SDFFR_X1 dscratch0_q_reg_30_ ( .D(n4144), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[30]) );
  SDFFR_X1 dscratch1_q_reg_30_ ( .D(n931), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[30]) );
  SDFFR_X1 utvec_q_reg_22_ ( .D(n931), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[22]), .QN(n1467) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__30_ ( .D(hwlp_data_o[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[30]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__30_ ( .D(n931), .SI(1'b0), .SE(1'b0), 
        .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[62]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__30_ ( .D(n931), .SI(1'b0), .SE(1'b0), 
        .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[94]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__30_ ( .D(hwlp_data_o[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[126]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__30_ ( .D(hwlp_data_o[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[158]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__30_ ( .D(hwlp_data_o[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[190]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__30_ ( .D(hwlp_data_o[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[222]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__30_ ( .D(hwlp_data_o[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[254]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__9__30_ ( .D(hwlp_data_o[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n4180), .RN(rst_n), .Q(pmp_addr_o[318]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__30_ ( .D(hwlp_data_o[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[350]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__30_ ( .D(hwlp_data_o[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[382]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__30_ ( .D(n931), .SI(1'b0), .SE(1'b0), 
        .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[414]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__30_ ( .D(n931), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[446]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__30_ ( .D(hwlp_data_o[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[478]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__30_ ( .D(hwlp_data_o[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[510]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__3__6_ ( .D(hwlp_data_o[30]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(n43) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__7__6_ ( .D(hwlp_data_o[30]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(n31) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__11__6_ ( .D(hwlp_data_o[30]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(n19) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__15__6_ ( .D(hwlp_data_o[30]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(n7) );
  SDFFR_X1 uepc_q_reg_31_ ( .D(n3998), .SI(1'b0), .SE(1'b0), .CK(n3999), .RN(
        rst_n), .Q(uepc_o[31]) );
  SDFFR_X1 mcause_q_reg_5_ ( .D(n3931), .SI(1'b0), .SE(1'b0), .CK(n3932), .RN(
        rst_n), .Q(mcause_q[5]) );
  SDFFR_X1 depc_q_reg_31_ ( .D(n4030), .SI(1'b0), .SE(1'b0), .CK(n4031), .RN(
        rst_n), .Q(depc_o[31]) );
  SDFFR_X1 mepc_q_reg_31_ ( .D(n4064), .SI(1'b0), .SE(1'b0), .CK(n4065), .RN(
        rst_n), .Q(mepc_o[31]) );
  SDFFR_X1 ucause_q_reg_5_ ( .D(n3941), .SI(1'b0), .SE(1'b0), .CK(n3942), .RN(
        rst_n), .Q(ucause_q[5]) );
  SDFFR_X1 mtvec_q_reg_23_ ( .D(n3961), .SI(1'b0), .SE(1'b0), .CK(n3962), .RN(
        rst_n), .Q(mtvec_o[23]) );
  SDFFR_X1 mscratch_q_reg_31_ ( .D(n4100), .SI(1'b0), .SE(1'b0), .CK(n4097), 
        .RN(rst_n), .Q(mscratch_q[31]) );
  SDFFR_X1 dscratch0_q_reg_31_ ( .D(n4148), .SI(1'b0), .SE(1'b0), .CK(n4145), 
        .RN(rst_n), .Q(dscratch0_q[31]) );
  SDFFR_X1 dscratch1_q_reg_31_ ( .D(n935), .SI(1'b0), .SE(1'b0), .CK(n4101), 
        .RN(rst_n), .Q(dscratch1_q[31]) );
  SDFFR_X1 utvec_q_reg_23_ ( .D(n2663), .SI(1'b0), .SE(1'b0), .CK(n3958), .RN(
        rst_n), .Q(utvec_o[23]), .QN(n1469) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__0__31_ ( .D(hwlp_data_o[31]), .SI(1'b0), 
        .SE(1'b0), .CK(n4149), .RN(rst_n), .Q(pmp_addr_o[31]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__1__31_ ( .D(n935), .SI(1'b0), .SE(1'b0), 
        .CK(n4163), .RN(rst_n), .Q(pmp_addr_o[63]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__2__31_ ( .D(n935), .SI(1'b0), .SE(1'b0), 
        .CK(n4165), .RN(rst_n), .Q(pmp_addr_o[95]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__3__31_ ( .D(n935), .SI(1'b0), .SE(1'b0), 
        .CK(n4167), .RN(rst_n), .Q(pmp_addr_o[127]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__4__31_ ( .D(n935), .SI(1'b0), .SE(1'b0), 
        .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[159]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__5__31_ ( .D(hwlp_data_o[31]), .SI(1'b0), 
        .SE(1'b0), .CK(n4171), .RN(rst_n), .Q(pmp_addr_o[191]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__31_ ( .D(n935), .SI(1'b0), .SE(1'b0), 
        .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[223]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__7__31_ ( .D(hwlp_data_o[31]), .SI(1'b0), 
        .SE(1'b0), .CK(n4176), .RN(rst_n), .Q(pmp_addr_o[255]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__31_ ( .D(hwlp_data_o[31]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[287]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__10__31_ ( .D(hwlp_data_o[31]), .SI(1'b0), 
        .SE(1'b0), .CK(n4151), .RN(rst_n), .Q(pmp_addr_o[351]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__11__31_ ( .D(hwlp_data_o[31]), .SI(1'b0), 
        .SE(1'b0), .CK(n4153), .RN(rst_n), .Q(pmp_addr_o[383]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__12__31_ ( .D(n935), .SI(1'b0), .SE(1'b0), 
        .CK(n4155), .RN(rst_n), .Q(pmp_addr_o[415]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__13__31_ ( .D(n935), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[447]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__14__31_ ( .D(n935), .SI(1'b0), .SE(1'b0), 
        .CK(n4159), .RN(rst_n), .Q(pmp_addr_o[479]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__15__31_ ( .D(hwlp_data_o[31]), .SI(1'b0), 
        .SE(1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[511]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__3__7_ ( .D(hwlp_data_o[31]), .SI(1'b0), .SE(
        1'b0), .CK(n3970), .RN(rst_n), .Q(n42) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__7__7_ ( .D(hwlp_data_o[31]), .SI(1'b0), .SE(
        1'b0), .CK(n3948), .RN(rst_n), .Q(n30) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__11__7_ ( .D(hwlp_data_o[31]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(n18) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__15__7_ ( .D(hwlp_data_o[31]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(n6) );
  SDFFS_X1 PCMR_q_reg_1_ ( .D(PCMR_n[1]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .SN(rst_n), .Q(PCMR_q[1]), .QN(n1584) );
  SDFFS_X1 PCMR_q_reg_0_ ( .D(PCMR_n[0]), .SI(1'b0), .SE(1'b0), .CK(n3911), 
        .SN(rst_n), .Q(PCMR_q[0]), .QN(n1456) );
  SDFFS_X1 mstatus_q_reg_mpp__1_ ( .D(mstatus_n[1]), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(rst_n), .Q(mstatus_q[2]) );
  SDFFS_X1 mstatus_q_reg_mpp__0_ ( .D(mstatus_n[0]), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(rst_n), .Q(mstatus_q[1]) );
  SDFFS_X1 dcsr_q_reg_prv__0_ ( .D(n3920), .SI(1'b0), .SE(1'b0), .CK(n3922), 
        .SN(rst_n), .Q(dcsr_q_prv__0_) );
  SDFFS_X1 dcsr_q_reg_prv__1_ ( .D(n3921), .SI(1'b0), .SE(1'b0), .CK(n3922), 
        .SN(rst_n), .Q(dcsr_q_prv__1_) );
  SDFFR_X1 id_valid_q_reg ( .D(id_valid_i), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(rst_n), .Q(id_valid_q) );
  SDFFS_X1 pmp_reg_q_reg_pmpaddr__9__31_ ( .D(n1441), .SI(1'b0), .SE(1'b0), 
        .CK(n4180), .SN(rst_n), .QN(pmp_addr_o[319]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__5__3_ ( .D(n2105), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(pmp_cfg_o[43]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__15__4_ ( .D(n2026), .SI(1'b0), .SE(1'b0), 
        .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[124]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__4__2_ ( .D(n564), .SI(1'b0), .SE(1'b0), .CK(
        n3948), .RN(rst_n), .Q(pmp_cfg_o[34]) );
  SDFFS_X1 priv_lvl_q_reg_1_ ( .D(n2022), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        rst_n), .Q(priv_lvl_o[1]), .QN(n1459) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__12__4_ ( .D(hwlp_data_o[4]), .SI(1'b0), .SE(
        1'b0), .CK(n3967), .RN(rst_n), .Q(pmp_cfg_o[100]) );
  SDFFR_X1 pmp_reg_q_reg_pmpcfg__10__4_ ( .D(hwlp_data_o[20]), .SI(1'b0), .SE(
        1'b0), .CK(n3964), .RN(rst_n), .Q(pmp_cfg_o[84]) );
  SDFFS_X1 PCCR_q_reg_0__0_ ( .D(n1450), .SI(1'b0), .SE(1'b0), .CK(n3914), 
        .SN(rst_n), .QN(PCCR_q[0]) );
  INV_X1 U80 ( .A(hwlp_data_o[8]), .ZN(n1402) );
  SDFFR_X2 pmp_reg_q_reg_pmpaddr__15__1_ ( .D(hwlp_data_o[1]), .SI(1'b0), .SE(
        1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[481]) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_0 clk_gate_pmp_reg_q_reg_pmpaddr__9__31_ ( 
        .CLK(clk), .EN(n1688), .ENCLK(n4180), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_1 clk_gate_pmp_reg_q_reg_pmpaddr__8__31_ ( 
        .CLK(clk), .EN(n1692), .ENCLK(n4178), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_2 clk_gate_pmp_reg_q_reg_pmpaddr__7__31_ ( 
        .CLK(clk), .EN(n1695), .ENCLK(n4176), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_3 clk_gate_pmp_reg_q_reg_pmpaddr__6__31_ ( 
        .CLK(clk), .EN(n1684), .ENCLK(n4173), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_4 clk_gate_pmp_reg_q_reg_pmpaddr__5__31_ ( 
        .CLK(clk), .EN(n1687), .ENCLK(n4171), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_5 clk_gate_pmp_reg_q_reg_pmpaddr__4__31_ ( 
        .CLK(clk), .EN(n1686), .ENCLK(n4169), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_6 clk_gate_pmp_reg_q_reg_pmpaddr__3__31_ ( 
        .CLK(clk), .EN(n1685), .ENCLK(n4167), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_7 clk_gate_pmp_reg_q_reg_pmpaddr__2__31_ ( 
        .CLK(clk), .EN(n1698), .ENCLK(n4165), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_8 clk_gate_pmp_reg_q_reg_pmpaddr__1__31_ ( 
        .CLK(clk), .EN(n1693), .ENCLK(n4163), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_9 clk_gate_pmp_reg_q_reg_pmpaddr__15__31_ ( 
        .CLK(clk), .EN(n1690), .ENCLK(n4161), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_10 clk_gate_pmp_reg_q_reg_pmpaddr__14__31_ ( 
        .CLK(clk), .EN(n932), .ENCLK(n4159), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_11 clk_gate_pmp_reg_q_reg_pmpaddr__13__31_ ( 
        .CLK(clk), .EN(n928), .ENCLK(n4157), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_12 clk_gate_pmp_reg_q_reg_pmpaddr__12__31_ ( 
        .CLK(clk), .EN(n926), .ENCLK(n4155), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_13 clk_gate_pmp_reg_q_reg_pmpaddr__11__31_ ( 
        .CLK(clk), .EN(n1691), .ENCLK(n4153), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_14 clk_gate_pmp_reg_q_reg_pmpaddr__10__31_ ( 
        .CLK(clk), .EN(n1696), .ENCLK(n4151), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_15 clk_gate_pmp_reg_q_reg_pmpaddr__0__31_ ( 
        .CLK(clk), .EN(n1694), .ENCLK(n4149), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_16 clk_gate_dscratch0_q_reg_31_ ( 
        .CLK(clk), .EN(n4147), .ENCLK(n4145), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_17 clk_gate_dscratch1_q_reg_31_ ( 
        .CLK(clk), .EN(n1437), .ENCLK(n4101), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_18 clk_gate_mscratch_q_reg_31_ ( 
        .CLK(clk), .EN(n4099), .ENCLK(n4097), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_19 clk_gate_mepc_q_reg_31_ ( 
        .CLK(clk), .EN(n4067), .ENCLK(n4065), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_20 clk_gate_depc_q_reg_31_ ( 
        .CLK(clk), .EN(n4033), .ENCLK(n4031), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_21 clk_gate_uepc_q_reg_31_ ( 
        .CLK(clk), .EN(n4001), .ENCLK(n3999), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_22 clk_gate_pmp_reg_q_reg_pmpcfg__3__7_ ( 
        .CLK(clk), .EN(n1445), .ENCLK(n3970), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_23 clk_gate_pmp_reg_q_reg_pmpcfg__12__4_ ( 
        .CLK(clk), .EN(n3969), .ENCLK(n3967), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_24 clk_gate_pmp_reg_q_reg_pmpcfg__10__4_ ( 
        .CLK(clk), .EN(n3966), .ENCLK(n3964), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_25 clk_gate_mtvec_q_reg_23_ ( 
        .CLK(clk), .EN(n1399), .ENCLK(n3962), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_26 clk_gate_utvec_q_reg_22_ ( 
        .CLK(clk), .EN(n1403), .ENCLK(n3958), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_27 clk_gate_pmp_reg_q_reg_pmpcfg__4__2_ ( 
        .CLK(clk), .EN(n241), .ENCLK(n3948), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_28 clk_gate_dcsr_q_reg_zero2__27_ ( 
        .CLK(clk), .EN(n198), .ENCLK(n3946), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_29 clk_gate_ucause_q_reg_5_ ( 
        .CLK(clk), .EN(n3944), .ENCLK(n3942), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_30 clk_gate_mcause_q_reg_5_ ( 
        .CLK(clk), .EN(n3934), .ENCLK(n3932), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_31 clk_gate_dcsr_q_reg_prv__1_ ( 
        .CLK(clk), .EN(n3924), .ENCLK(n3922), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_32 clk_gate_PCCR_q_reg_0__9_ ( 
        .CLK(clk), .EN(n3916), .ENCLK(n3914), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16_33 clk_gate_mstatus_q_reg_mprv_ ( 
        .CLK(clk), .EN(n3913), .ENCLK(n3911), .TE(1'b0) );
  SDFFR_X2 pmp_reg_q_reg_pmpaddr__4__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4169), .RN(rst_n), .Q(pmp_addr_o[128]) );
  SDFFR_X2 pmp_reg_q_reg_pmpaddr__13__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[416]) );
  SDFFR_X2 pmp_reg_q_reg_pmpaddr__15__0_ ( .D(hwlp_data_o[0]), .SI(1'b0), .SE(
        1'b0), .CK(n4161), .RN(rst_n), .Q(pmp_addr_o[480]) );
  SDFFR_X2 pmp_reg_q_reg_pmpaddr__13__1_ ( .D(n1031), .SI(1'b0), .SE(1'b0), 
        .CK(n4157), .RN(rst_n), .Q(pmp_addr_o[417]) );
  SDFFR_X1 PCCR_q_reg_0__28_ ( .D(PCCR_n[27]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[28]), .QN(n1497) );
  SDFFR_X1 PCCR_q_reg_0__29_ ( .D(PCCR_n[28]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[29]), .QN(n1491) );
  SDFFR_X1 PCCR_q_reg_0__30_ ( .D(PCCR_n[29]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[30]), .QN(n1466) );
  SDFFR_X1 PCCR_q_reg_0__31_ ( .D(PCCR_n[30]), .SI(1'b0), .SE(1'b0), .CK(n3914), .RN(rst_n), .Q(PCCR_q[31]), .QN(n1505) );
  SDFFR_X2 priv_lvl_q_reg_0_ ( .D(n1449), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(
        rst_n), .Q(n1481), .QN(\priv_lvl_o[0] ) );
  INV_X1 U1972 ( .A(n1129), .ZN(n1125) );
  NOR2_X2 U1975 ( .A1(csr_save_ex_i_BAR), .A2(n1125), .ZN(n1141) );
  BUF_X1 U10 ( .A(n1012), .Z(n62) );
  BUF_X1 U8 ( .A(n1142), .Z(n58) );
  CLKBUF_X2 U12 ( .A(n1070), .Z(n55) );
  CLKBUF_X2 U3 ( .A(n1079), .Z(n57) );
  CLKBUF_X2 U6 ( .A(n1155), .Z(n60) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__6__21_ ( .D(hwlp_data_o[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n4173), .RN(rst_n), .Q(pmp_addr_o[213]) );
  SDFFR_X1 pmp_reg_q_reg_pmpaddr__8__30_ ( .D(hwlp_data_o[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n4178), .RN(rst_n), .Q(pmp_addr_o[286]) );
  CLKBUF_X1 U4 ( .A(n3884), .Z(n1705) );
  CLKBUF_X2 U5 ( .A(n971), .Z(n63) );
  INV_X2 U7 ( .A(n1050), .ZN(n1677) );
  NOR2_X1 U9 ( .A1(debug_csr_save_i), .A2(n1122), .ZN(n1129) );
  NAND2_X2 U13 ( .A1(n1209), .A2(n951), .ZN(n958) );
  INV_X1 U15 ( .A(n1412), .ZN(n1678) );
  INV_X2 U17 ( .A(n1404), .ZN(hwlp_data_o[11]) );
  INV_X2 U19 ( .A(n1405), .ZN(hwlp_data_o[12]) );
  INV_X1 U27 ( .A(n1447), .ZN(n1681) );
  INV_X1 U28 ( .A(n1444), .ZN(n1682) );
  INV_X2 U29 ( .A(n1390), .ZN(hwlp_data_o[4]) );
  INV_X1 U32 ( .A(n714), .ZN(n734) );
  CLKBUF_X1 U33 ( .A(n153), .Z(n691) );
  NOR2_X1 U34 ( .A1(n940), .A2(n1038), .ZN(n942) );
  CLKBUF_X2 U35 ( .A(n1057), .Z(n56) );
  NOR3_X1 U36 ( .A1(n133), .A2(n195), .A3(n1198), .ZN(n911) );
  OR2_X1 U37 ( .A1(n831), .A2(n1038), .ZN(n1212) );
  AND2_X1 U38 ( .A1(n911), .A2(n906), .ZN(n1684) );
  AND2_X1 U41 ( .A1(n911), .A2(n894), .ZN(n1685) );
  AND2_X1 U44 ( .A1(n911), .A2(n898), .ZN(n1686) );
  AND2_X1 U47 ( .A1(n911), .A2(n902), .ZN(n1687) );
  AND2_X1 U75 ( .A1(n923), .A2(n1046), .ZN(n1688) );
  AND3_X1 U76 ( .A1(n1370), .A2(n1373), .A3(n1372), .ZN(n1689) );
  AND2_X1 U77 ( .A1(n1371), .A2(n937), .ZN(n1690) );
  AND2_X1 U78 ( .A1(n923), .A2(n922), .ZN(n1691) );
  AND2_X1 U79 ( .A1(n923), .A2(n914), .ZN(n1692) );
  AND2_X1 U96 ( .A1(n911), .A2(n886), .ZN(n1693) );
  AND2_X1 U137 ( .A1(n911), .A2(n882), .ZN(n1694) );
  AND2_X1 U190 ( .A1(n911), .A2(n910), .ZN(n1695) );
  AND2_X1 U191 ( .A1(n923), .A2(n919), .ZN(n1696) );
  OR2_X1 U193 ( .A1(n1199), .A2(n1198), .ZN(n1697) );
  AND2_X1 U234 ( .A1(n911), .A2(n890), .ZN(n1698) );
  AND4_X1 U240 ( .A1(n145), .A2(n144), .A3(n143), .A4(n142), .ZN(n1699) );
  INV_X1 U241 ( .A(n4183), .ZN(n1700) );
  INV_X1 U243 ( .A(n1700), .ZN(hwlp_data_o[21]) );
  OAI21_X1 U245 ( .B1(n424), .B2(csr_wdata_i[21]), .A(n423), .ZN(n4183) );
  INV_X1 U246 ( .A(n4184), .ZN(n1702) );
  INV_X1 U255 ( .A(n1702), .ZN(hwlp_data_o[3]) );
  INV_X1 U277 ( .A(hwlp_data_o[26]), .ZN(n1704) );
  OAI21_X1 U278 ( .B1(n403), .B2(csr_wdata_i[26]), .A(n402), .ZN(
        hwlp_data_o[26]) );
  NAND2_X2 U283 ( .A1(n1046), .A2(n1373), .ZN(n1054) );
  INV_X1 U284 ( .A(n1415), .ZN(n3952) );
  INV_X1 U285 ( .A(n1411), .ZN(n3951) );
  INV_X1 U286 ( .A(n1704), .ZN(n3955) );
  INV_X1 U287 ( .A(n1418), .ZN(n3954) );
  INV_X1 U288 ( .A(n1421), .ZN(n3956) );
  INV_X1 U289 ( .A(n1422), .ZN(n3957) );
  INV_X1 U306 ( .A(n1416), .ZN(n3953) );
  INV_X1 U307 ( .A(n1426), .ZN(hwlp_data_o[30]) );
  INV_X2 U311 ( .A(n1689), .ZN(n1706) );
  INV_X1 U312 ( .A(n1402), .ZN(n4175) );
  NAND4_X1 U341 ( .A1(n1699), .A2(n163), .A3(n1714), .A4(n164), .ZN(
        csr_rdata_o[8]) );
  AND2_X1 U343 ( .A1(n162), .A2(n165), .ZN(n1714) );
  INV_X1 U344 ( .A(n1374), .ZN(n1395) );
  OR2_X2 U345 ( .A1(n118), .A2(n881), .ZN(n1374) );
  INV_X1 U346 ( .A(csr_access_i), .ZN(n1715) );
  INV_X1 U348 ( .A(n1441), .ZN(hwlp_data_o[31]) );
  INV_X1 U349 ( .A(n935), .ZN(n1441) );
  NOR2_X1 U350 ( .A1(n1054), .A2(n1677), .ZN(n3833) );
  AOI21_X1 U351 ( .B1(csr_save_cause_i), .B2(n1048), .A(n3925), .ZN(n1050) );
  INV_X1 U370 ( .A(n1129), .ZN(n3890) );
  NOR4_X1 U3225 ( .A1(csr_addr_i[1]), .A2(csr_addr_i[2]), .A3(n1394), .A4(
        n3692), .ZN(n3913) );
  OAI221_X1 U3226 ( .B1(csr_addr_i[7]), .B2(n3693), .C1(csr_addr_i[7]), .C2(
        n3694), .A(n3695), .ZN(n3692) );
  AOI211_X1 U3227 ( .C1(csr_addr_i[7]), .C2(n3696), .A(csr_addr_i[4]), .B(
        csr_addr_i[3]), .ZN(n3695) );
  NAND3_X1 U3228 ( .A1(csr_addr_i[6]), .A2(csr_addr_i[10]), .A3(n3697), .ZN(
        n3696) );
  AOI21_X1 U3229 ( .B1(csr_addr_i[5]), .B2(n3698), .A(n3699), .ZN(n3697) );
  AOI21_X1 U3230 ( .B1(csr_addr_i[11]), .B2(n155), .A(csr_addr_i[5]), .ZN(
        n3699) );
  NOR4_X1 U3231 ( .A1(csr_addr_i[6]), .A2(csr_addr_i[5]), .A3(csr_addr_i[10]), 
        .A4(csr_addr_i[0]), .ZN(n3694) );
  INV_X1 U3232 ( .A(n3698), .ZN(n3693) );
  NAND3_X1 U3233 ( .A1(csr_addr_i[8]), .A2(csr_addr_i[9]), .A3(n3700), .ZN(
        n3698) );
  INV_X1 U3234 ( .A(csr_addr_i[11]), .ZN(n3700) );
  INV_X1 U3235 ( .A(n3701), .ZN(n3916) );
  AOI221_X1 U3236 ( .B1(n814), .B2(n790), .C1(csr_op_i[0]), .C2(n790), .A(
        PCCR_inc_q_0_), .ZN(n3701) );
  OAI21_X1 U3237 ( .B1(debug_cause_i[2]), .B2(n1221), .A(n3702), .ZN(n3917) );
  NAND2_X1 U3238 ( .A1(n1221), .A2(hwlp_data_o[6]), .ZN(n3702) );
  MUX2_X1 U3239 ( .A(debug_cause_i[2]), .B(hwlp_data_o[8]), .S(n1221), .Z(
        n3918) );
  MUX2_X1 U3240 ( .A(n4116), .B(debug_cause_i[1]), .S(n3925), .Z(n3919) );
  OR2_X1 U3241 ( .A1(n3925), .A2(\priv_lvl_o[0] ), .ZN(n3920) );
  OR2_X1 U3242 ( .A1(n3925), .A2(priv_lvl_o[1]), .ZN(n3921) );
  OR2_X1 U3243 ( .A1(n198), .A2(n3925), .ZN(n3924) );
  INV_X1 U3244 ( .A(n1221), .ZN(n3925) );
  MUX2_X1 U3245 ( .A(n1031), .B(n3936), .S(n1037), .Z(n3926) );
  MUX2_X1 U3246 ( .A(n564), .B(csr_cause_i_2_), .S(n1037), .Z(n3927) );
  MUX2_X1 U3247 ( .A(hwlp_data_o[4]), .B(csr_cause_i_4_), .S(n1037), .Z(n3928)
         );
  MUX2_X1 U3248 ( .A(hwlp_data_o[3]), .B(csr_cause_i_3_), .S(n1037), .Z(n3929)
         );
  MUX2_X1 U3249 ( .A(hwlp_data_o[0]), .B(csr_cause_i_0_), .S(n1037), .Z(n3930)
         );
  AOI22_X1 U3250 ( .A1(n3703), .A2(n1441), .B1(n1045), .B2(csr_cause_i_5__BAR), 
        .ZN(n3931) );
  OAI21_X1 U3251 ( .B1(csr_irq_sec_i), .B2(n1042), .A(n1045), .ZN(n3703) );
  OR2_X1 U3252 ( .A1(n1041), .A2(n1037), .ZN(n3934) );
  MUX2_X1 U3253 ( .A(n3936), .B(hwlp_data_o[1]), .S(n1212), .Z(n3935) );
  INV_X1 U3254 ( .A(csr_cause_i_1__BAR), .ZN(n3936) );
  MUX2_X1 U3255 ( .A(csr_cause_i_2_), .B(n4113), .S(n1212), .Z(n3937) );
  MUX2_X1 U3256 ( .A(csr_cause_i_4_), .B(hwlp_data_o[4]), .S(n1212), .Z(n3938)
         );
  MUX2_X1 U3257 ( .A(csr_cause_i_3_), .B(n4184), .S(n1212), .Z(n3939) );
  MUX2_X1 U3258 ( .A(csr_cause_i_0_), .B(hwlp_data_o[0]), .S(n1212), .Z(n3940)
         );
  NAND2_X1 U3259 ( .A1(n1212), .A2(n1441), .ZN(n3941) );
  NAND2_X1 U3260 ( .A1(n1212), .A2(n1697), .ZN(n3944) );
  AND2_X1 U3261 ( .A1(hwlp_data_o[31]), .A2(n1429), .ZN(n3961) );
  OAI21_X1 U3262 ( .B1(n958), .B2(n3704), .A(n3705), .ZN(n3972) );
  AOI22_X1 U3263 ( .A1(pc_id_i[5]), .A2(n3750), .B1(n958), .B2(hwlp_data_o[5]), 
        .ZN(n3705) );
  AOI22_X1 U3264 ( .A1(pc_if_i[5]), .A2(n3907), .B1(pc_ex_i[5]), .B2(n3723), 
        .ZN(n3704) );
  OAI211_X1 U3265 ( .C1(n958), .C2(n3706), .A(n3707), .B(n3708), .ZN(n3973) );
  NAND2_X1 U3266 ( .A1(n958), .A2(n1681), .ZN(n3708) );
  NAND2_X1 U3267 ( .A1(n62), .A2(pc_id_i[9]), .ZN(n3707) );
  AOI21_X1 U3268 ( .B1(pc_ex_i[9]), .B2(n3723), .A(n4038), .ZN(n3706) );
  NAND2_X1 U3269 ( .A1(n983), .A2(n3709), .ZN(n3974) );
  AOI22_X1 U3270 ( .A1(pc_if_i[10]), .A2(n3732), .B1(n958), .B2(n1682), .ZN(
        n3709) );
  NAND2_X1 U3271 ( .A1(n975), .A2(n3710), .ZN(n3975) );
  AOI22_X1 U3272 ( .A1(pc_if_i[6]), .A2(n3732), .B1(n958), .B2(hwlp_data_o[6]), 
        .ZN(n3710) );
  NAND2_X1 U3273 ( .A1(n979), .A2(n3711), .ZN(n3976) );
  AOI22_X1 U3274 ( .A1(pc_ex_i[8]), .A2(n63), .B1(n958), .B2(n4175), .ZN(n3711) );
  OAI211_X1 U3275 ( .C1(n958), .C2(n3712), .A(n3713), .B(n3714), .ZN(n3977) );
  NAND2_X1 U3276 ( .A1(n958), .A2(hwlp_data_o[1]), .ZN(n3714) );
  NAND2_X1 U3277 ( .A1(n62), .A2(pc_id_i[1]), .ZN(n3713) );
  AOI22_X1 U3278 ( .A1(pc_if_i[1]), .A2(n3907), .B1(pc_ex_i[1]), .B2(n3723), 
        .ZN(n3712) );
  NAND2_X1 U3279 ( .A1(n964), .A2(n3715), .ZN(n3978) );
  AOI22_X1 U3280 ( .A1(pc_if_i[2]), .A2(n3732), .B1(n958), .B2(n4113), .ZN(
        n3715) );
  NAND2_X1 U3281 ( .A1(n966), .A2(n3716), .ZN(n3979) );
  AOI22_X1 U3282 ( .A1(pc_if_i[3]), .A2(n3732), .B1(n958), .B2(hwlp_data_o[3]), 
        .ZN(n3716) );
  OAI21_X1 U3283 ( .B1(n958), .B2(n3717), .A(n3718), .ZN(n3980) );
  AOI22_X1 U3284 ( .A1(pc_id_i[7]), .A2(n3750), .B1(n958), .B2(n4116), .ZN(
        n3718) );
  AOI21_X1 U3285 ( .B1(pc_ex_i[7]), .B2(n3723), .A(n4047), .ZN(n3717) );
  NAND2_X1 U3286 ( .A1(n989), .A2(n3719), .ZN(n3981) );
  AOI22_X1 U3287 ( .A1(pc_if_i[13]), .A2(n3732), .B1(n958), .B2(n3960), .ZN(
        n3719) );
  OAI211_X1 U3288 ( .C1(n1126), .C2(n3720), .A(n3721), .B(n3722), .ZN(n3982)
         );
  NAND3_X1 U3289 ( .A1(pc_ex_i[14]), .A2(n3723), .A3(n3748), .ZN(n3722) );
  INV_X1 U3290 ( .A(csr_save_ex_i_BAR), .ZN(n3723) );
  AOI22_X1 U3291 ( .A1(n64), .A2(pc_if_i[14]), .B1(hwlp_data_o[14]), .B2(n958), 
        .ZN(n3721) );
  NAND2_X1 U3292 ( .A1(pc_id_i[14]), .A2(n3748), .ZN(n3720) );
  OAI211_X1 U3293 ( .C1(n958), .C2(n3724), .A(n3725), .B(n3726), .ZN(n3983) );
  NAND2_X1 U3294 ( .A1(n958), .A2(hwlp_data_o[15]), .ZN(n3726) );
  NAND2_X1 U3295 ( .A1(n62), .A2(pc_id_i[15]), .ZN(n3725) );
  AOI22_X1 U3296 ( .A1(pc_if_i[15]), .A2(n3907), .B1(pc_ex_i[15]), .B2(n3723), 
        .ZN(n3724) );
  NAND2_X1 U3297 ( .A1(n998), .A2(n3727), .ZN(n3984) );
  AOI22_X1 U3298 ( .A1(pc_if_i[17]), .A2(n3732), .B1(n958), .B2(
        hwlp_data_o[17]), .ZN(n3727) );
  NAND2_X1 U3299 ( .A1(n1000), .A2(n3728), .ZN(n3985) );
  AOI22_X1 U3300 ( .A1(pc_ex_i[18]), .A2(n971), .B1(n958), .B2(hwlp_data_o[18]), .ZN(n3728) );
  NAND2_X1 U3301 ( .A1(n1002), .A2(n3729), .ZN(n3986) );
  AOI22_X1 U3302 ( .A1(pc_id_i[19]), .A2(n3750), .B1(n958), .B2(
        hwlp_data_o[19]), .ZN(n3729) );
  NAND2_X1 U3303 ( .A1(n1004), .A2(n3730), .ZN(n3987) );
  AOI22_X1 U3304 ( .A1(pc_ex_i[20]), .A2(n971), .B1(n958), .B2(n1678), .ZN(
        n3730) );
  NAND2_X1 U3305 ( .A1(n1006), .A2(n3731), .ZN(n3988) );
  AOI22_X1 U3306 ( .A1(pc_if_i[21]), .A2(n3732), .B1(n958), .B2(n4183), .ZN(
        n3731) );
  NOR2_X1 U3307 ( .A1(n1124), .A2(n958), .ZN(n3732) );
  NAND2_X1 U3308 ( .A1(n1009), .A2(n3733), .ZN(n3989) );
  AOI22_X1 U3309 ( .A1(pc_if_i[22]), .A2(n3732), .B1(n958), .B2(
        hwlp_data_o[22]), .ZN(n3733) );
  NAND2_X1 U3310 ( .A1(n1011), .A2(n3734), .ZN(n3990) );
  AOI22_X1 U3311 ( .A1(pc_ex_i[23]), .A2(n971), .B1(n958), .B2(n3952), .ZN(
        n3734) );
  OAI211_X1 U3312 ( .C1(n958), .C2(n3735), .A(n3736), .B(n3737), .ZN(n3991) );
  NAND2_X1 U3313 ( .A1(n958), .A2(hwlp_data_o[24]), .ZN(n3737) );
  NAND2_X1 U3314 ( .A1(n64), .A2(pc_if_i[24]), .ZN(n3736) );
  AOI22_X1 U3315 ( .A1(pc_id_i[24]), .A2(n3838), .B1(pc_ex_i[24]), .B2(n3723), 
        .ZN(n3735) );
  OAI211_X1 U3316 ( .C1(n1124), .C2(n3738), .A(n3739), .B(n3740), .ZN(n3992)
         );
  NAND3_X1 U3317 ( .A1(pc_id_i[25]), .A2(n3838), .A3(n3748), .ZN(n3740) );
  AOI22_X1 U3318 ( .A1(n63), .A2(pc_ex_i[25]), .B1(n3954), .B2(n958), .ZN(
        n3739) );
  NAND2_X1 U3319 ( .A1(pc_if_i[25]), .A2(n3748), .ZN(n3738) );
  NAND2_X1 U3320 ( .A1(n1018), .A2(n3741), .ZN(n3993) );
  AOI22_X1 U3321 ( .A1(pc_id_i[26]), .A2(n3750), .B1(n958), .B2(n3955), .ZN(
        n3741) );
  NAND2_X1 U3322 ( .A1(n1020), .A2(n3742), .ZN(n3994) );
  AOI22_X1 U3323 ( .A1(pc_ex_i[27]), .A2(n971), .B1(n958), .B2(n3956), .ZN(
        n3742) );
  NAND2_X1 U3324 ( .A1(n1022), .A2(n3743), .ZN(n3995) );
  AOI22_X1 U3325 ( .A1(pc_ex_i[28]), .A2(n63), .B1(n958), .B2(hwlp_data_o[28]), 
        .ZN(n3743) );
  NAND2_X1 U3326 ( .A1(n1024), .A2(n3744), .ZN(n3996) );
  AOI22_X1 U3327 ( .A1(pc_id_i[29]), .A2(n3750), .B1(n958), .B2(n4143), .ZN(
        n3744) );
  OAI211_X1 U3328 ( .C1(n1124), .C2(n3745), .A(n3746), .B(n3747), .ZN(n3997)
         );
  NAND3_X1 U3329 ( .A1(pc_id_i[30]), .A2(n3838), .A3(n3748), .ZN(n3747) );
  AOI22_X1 U3330 ( .A1(n63), .A2(pc_ex_i[30]), .B1(hwlp_data_o[30]), .B2(n958), 
        .ZN(n3746) );
  NAND2_X1 U3331 ( .A1(pc_if_i[30]), .A2(n3748), .ZN(n3745) );
  INV_X1 U3332 ( .A(n958), .ZN(n3748) );
  NAND2_X1 U3333 ( .A1(n1028), .A2(n3749), .ZN(n3998) );
  AOI22_X1 U3334 ( .A1(pc_id_i[31]), .A2(n3750), .B1(n958), .B2(
        hwlp_data_o[31]), .ZN(n3749) );
  NOR2_X1 U3335 ( .A1(n1126), .A2(n958), .ZN(n3750) );
  NAND2_X1 U3336 ( .A1(n958), .A2(n956), .ZN(n4001) );
  NAND2_X1 U3337 ( .A1(n1051), .A2(n3751), .ZN(n4002) );
  NAND2_X1 U3338 ( .A1(pc_if_i[0]), .A2(n56), .ZN(n3751) );
  NAND2_X1 U3339 ( .A1(n1065), .A2(n3752), .ZN(n4003) );
  AOI21_X1 U3340 ( .B1(pc_ex_i[5]), .B2(n55), .A(n3753), .ZN(n3752) );
  NOR3_X1 U3341 ( .A1(n1677), .A2(n1054), .A3(n3754), .ZN(n3753) );
  NAND2_X1 U3342 ( .A1(n1385), .A2(hwlp_data_o[5]), .ZN(n3754) );
  NAND2_X1 U3343 ( .A1(n1074), .A2(n3755), .ZN(n4004) );
  AOI21_X1 U3344 ( .B1(n55), .B2(pc_ex_i[9]), .A(n3756), .ZN(n3755) );
  NOR3_X1 U3345 ( .A1(n1677), .A2(n1054), .A3(n3757), .ZN(n3756) );
  NAND2_X1 U3346 ( .A1(n1385), .A2(n1681), .ZN(n3757) );
  NAND2_X1 U3347 ( .A1(n1076), .A2(n3758), .ZN(n4005) );
  AOI21_X1 U3348 ( .B1(n55), .B2(pc_ex_i[10]), .A(n3759), .ZN(n3758) );
  NOR3_X1 U3349 ( .A1(n1677), .A2(n1054), .A3(n3760), .ZN(n3759) );
  NAND2_X1 U3350 ( .A1(n1385), .A2(n1682), .ZN(n3760) );
  NAND2_X1 U3351 ( .A1(n1067), .A2(n3761), .ZN(n4006) );
  AOI21_X1 U3352 ( .B1(n57), .B2(pc_id_i[6]), .A(n3762), .ZN(n3761) );
  NOR3_X1 U3353 ( .A1(n1677), .A2(n1054), .A3(n3763), .ZN(n3762) );
  NAND2_X1 U3354 ( .A1(n1385), .A2(hwlp_data_o[6]), .ZN(n3763) );
  NAND2_X1 U3355 ( .A1(n1072), .A2(n3764), .ZN(n4007) );
  AOI21_X1 U3356 ( .B1(n55), .B2(pc_ex_i[8]), .A(n3765), .ZN(n3764) );
  NOR3_X1 U3357 ( .A1(n1677), .A2(n1054), .A3(n3766), .ZN(n3765) );
  NAND2_X1 U3358 ( .A1(n1385), .A2(n4175), .ZN(n3766) );
  NAND2_X1 U3359 ( .A1(n1056), .A2(n3767), .ZN(n4008) );
  AOI21_X1 U3360 ( .B1(pc_ex_i[1]), .B2(n55), .A(n3768), .ZN(n3767) );
  NOR3_X1 U3361 ( .A1(n1677), .A2(n1054), .A3(n3769), .ZN(n3768) );
  NAND2_X1 U3362 ( .A1(n1385), .A2(hwlp_data_o[1]), .ZN(n3769) );
  NAND2_X1 U3363 ( .A1(n1059), .A2(n3770), .ZN(n4009) );
  AOI21_X1 U3364 ( .B1(n57), .B2(pc_id_i[2]), .A(n3771), .ZN(n3770) );
  NOR3_X1 U3365 ( .A1(n1677), .A2(n1054), .A3(n3772), .ZN(n3771) );
  NAND2_X1 U3366 ( .A1(n1385), .A2(n4113), .ZN(n3772) );
  OAI211_X1 U3367 ( .C1(n1124), .C2(n3773), .A(n3774), .B(n3775), .ZN(n4010)
         );
  NAND3_X1 U3368 ( .A1(hwlp_data_o[4]), .A2(n1385), .A3(n3833), .ZN(n3775) );
  AOI22_X1 U3369 ( .A1(n55), .A2(pc_ex_i[4]), .B1(pc_id_i[4]), .B2(n1079), 
        .ZN(n3774) );
  NAND2_X1 U3370 ( .A1(pc_if_i[4]), .A2(n1677), .ZN(n3773) );
  NAND2_X1 U3371 ( .A1(n1061), .A2(n3776), .ZN(n4011) );
  AOI21_X1 U3372 ( .B1(n57), .B2(pc_id_i[3]), .A(n3777), .ZN(n3776) );
  NOR3_X1 U3373 ( .A1(n1677), .A2(n1054), .A3(n3778), .ZN(n3777) );
  NAND2_X1 U3374 ( .A1(n1385), .A2(n4184), .ZN(n3778) );
  NAND2_X1 U3375 ( .A1(n1069), .A2(n3779), .ZN(n4012) );
  AOI21_X1 U3376 ( .B1(n56), .B2(pc_if_i[7]), .A(n3780), .ZN(n3779) );
  NOR3_X1 U3377 ( .A1(n1677), .A2(n1054), .A3(n3781), .ZN(n3780) );
  NAND2_X1 U3378 ( .A1(n1385), .A2(n4116), .ZN(n3781) );
  NAND2_X1 U3379 ( .A1(n1078), .A2(n3782), .ZN(n4013) );
  AOI21_X1 U3380 ( .B1(n56), .B2(pc_if_i[11]), .A(n3783), .ZN(n3782) );
  NOR3_X1 U3381 ( .A1(n1677), .A2(n1054), .A3(n3784), .ZN(n3783) );
  NAND2_X1 U3382 ( .A1(n1385), .A2(hwlp_data_o[11]), .ZN(n3784) );
  NAND2_X1 U3383 ( .A1(n1081), .A2(n3785), .ZN(n4014) );
  AOI21_X1 U3384 ( .B1(n56), .B2(pc_if_i[12]), .A(n3786), .ZN(n3785) );
  NOR3_X1 U3385 ( .A1(n1677), .A2(n1054), .A3(n3787), .ZN(n3786) );
  NAND2_X1 U3386 ( .A1(n1385), .A2(hwlp_data_o[12]), .ZN(n3787) );
  OAI211_X1 U3387 ( .C1(n1126), .C2(n3788), .A(n3789), .B(n3790), .ZN(n4015)
         );
  NAND3_X1 U3388 ( .A1(n3960), .A2(n1385), .A3(n3833), .ZN(n3790) );
  AOI22_X1 U3389 ( .A1(n55), .A2(pc_ex_i[13]), .B1(pc_if_i[13]), .B2(n56), 
        .ZN(n3789) );
  NAND2_X1 U3390 ( .A1(pc_id_i[13]), .A2(n1677), .ZN(n3788) );
  NAND2_X1 U3391 ( .A1(n1085), .A2(n3791), .ZN(n4016) );
  AOI21_X1 U3392 ( .B1(n56), .B2(pc_if_i[14]), .A(n3792), .ZN(n3791) );
  NOR3_X1 U3393 ( .A1(n1677), .A2(n1054), .A3(n3793), .ZN(n3792) );
  NAND2_X1 U3394 ( .A1(n1385), .A2(hwlp_data_o[14]), .ZN(n3793) );
  NAND2_X1 U3395 ( .A1(n1087), .A2(n3794), .ZN(n4017) );
  AOI21_X1 U3396 ( .B1(n56), .B2(pc_if_i[15]), .A(n3795), .ZN(n3794) );
  NOR3_X1 U3397 ( .A1(n1677), .A2(n1054), .A3(n3796), .ZN(n3795) );
  NAND2_X1 U3398 ( .A1(n1385), .A2(hwlp_data_o[15]), .ZN(n3796) );
  NAND2_X1 U3399 ( .A1(n1094), .A2(n3797), .ZN(n4018) );
  AOI21_X1 U3400 ( .B1(n55), .B2(pc_ex_i[18]), .A(n3798), .ZN(n3797) );
  NOR3_X1 U3401 ( .A1(n1677), .A2(n1054), .A3(n3799), .ZN(n3798) );
  NAND2_X1 U3402 ( .A1(n1385), .A2(hwlp_data_o[18]), .ZN(n3799) );
  NAND2_X1 U3403 ( .A1(n1096), .A2(n3800), .ZN(n4019) );
  AOI21_X1 U3404 ( .B1(n55), .B2(pc_ex_i[19]), .A(n3801), .ZN(n3800) );
  NOR3_X1 U3405 ( .A1(n1677), .A2(n1054), .A3(n3802), .ZN(n3801) );
  NAND2_X1 U3406 ( .A1(n1385), .A2(hwlp_data_o[19]), .ZN(n3802) );
  NAND2_X1 U3407 ( .A1(n1098), .A2(n3803), .ZN(n4020) );
  AOI21_X1 U3408 ( .B1(n55), .B2(pc_ex_i[20]), .A(n3804), .ZN(n3803) );
  NOR3_X1 U3409 ( .A1(n1677), .A2(n1054), .A3(n3805), .ZN(n3804) );
  NAND2_X1 U3410 ( .A1(n1385), .A2(n1678), .ZN(n3805) );
  NAND2_X1 U3411 ( .A1(n1100), .A2(n3806), .ZN(n4021) );
  AOI21_X1 U3412 ( .B1(n1079), .B2(pc_id_i[21]), .A(n3807), .ZN(n3806) );
  NOR3_X1 U3413 ( .A1(n1677), .A2(n1054), .A3(n3808), .ZN(n3807) );
  NAND2_X1 U3414 ( .A1(n1385), .A2(hwlp_data_o[21]), .ZN(n3808) );
  NAND2_X1 U3415 ( .A1(n1102), .A2(n3809), .ZN(n4022) );
  AOI21_X1 U3416 ( .B1(pc_ex_i[22]), .B2(n55), .A(n3810), .ZN(n3809) );
  NOR3_X1 U3417 ( .A1(n1677), .A2(n1054), .A3(n3811), .ZN(n3810) );
  NAND2_X1 U3418 ( .A1(n1385), .A2(n1007), .ZN(n3811) );
  OAI211_X1 U3419 ( .C1(n1126), .C2(n3812), .A(n3813), .B(n3814), .ZN(n4023)
         );
  NAND3_X1 U3420 ( .A1(n3952), .A2(n1385), .A3(n3833), .ZN(n3814) );
  AOI22_X1 U3421 ( .A1(n55), .A2(pc_ex_i[23]), .B1(pc_if_i[23]), .B2(n56), 
        .ZN(n3813) );
  NAND2_X1 U3422 ( .A1(pc_id_i[23]), .A2(n1677), .ZN(n3812) );
  NAND2_X1 U3423 ( .A1(n1106), .A2(n3815), .ZN(n4024) );
  AOI21_X1 U3424 ( .B1(n55), .B2(pc_ex_i[24]), .A(n3816), .ZN(n3815) );
  NOR3_X1 U3425 ( .A1(n1677), .A2(n1054), .A3(n3817), .ZN(n3816) );
  NAND2_X1 U3426 ( .A1(n1385), .A2(hwlp_data_o[24]), .ZN(n3817) );
  NAND2_X1 U3427 ( .A1(n1109), .A2(n3818), .ZN(n4025) );
  AOI21_X1 U3428 ( .B1(pc_if_i[25]), .B2(n56), .A(n3819), .ZN(n3818) );
  NOR3_X1 U3429 ( .A1(n1677), .A2(n1054), .A3(n3820), .ZN(n3819) );
  NAND2_X1 U3430 ( .A1(n1385), .A2(n3954), .ZN(n3820) );
  OAI211_X1 U3431 ( .C1(n1124), .C2(n3821), .A(n3822), .B(n3823), .ZN(n4026)
         );
  NAND3_X1 U3432 ( .A1(n3955), .A2(n1385), .A3(n3833), .ZN(n3823) );
  AOI22_X1 U3433 ( .A1(n55), .A2(pc_ex_i[26]), .B1(pc_id_i[26]), .B2(n1079), 
        .ZN(n3822) );
  NAND2_X1 U3434 ( .A1(pc_if_i[26]), .A2(n1677), .ZN(n3821) );
  NAND2_X1 U3435 ( .A1(n1113), .A2(n3824), .ZN(n4027) );
  AOI21_X1 U3436 ( .B1(n55), .B2(pc_ex_i[27]), .A(n3825), .ZN(n3824) );
  NOR3_X1 U3437 ( .A1(n1677), .A2(n1054), .A3(n3826), .ZN(n3825) );
  NAND2_X1 U3438 ( .A1(n1385), .A2(hwlp_data_o[27]), .ZN(n3826) );
  NAND2_X1 U3439 ( .A1(n1115), .A2(n3827), .ZN(n4028) );
  AOI21_X1 U3440 ( .B1(n1057), .B2(pc_if_i[28]), .A(n3828), .ZN(n3827) );
  NOR3_X1 U3441 ( .A1(n1677), .A2(n1054), .A3(n3829), .ZN(n3828) );
  NAND2_X1 U3442 ( .A1(n1385), .A2(hwlp_data_o[28]), .ZN(n3829) );
  OAI211_X1 U3443 ( .C1(n1124), .C2(n3830), .A(n3831), .B(n3832), .ZN(n4029)
         );
  NAND3_X1 U3444 ( .A1(n4143), .A2(n1385), .A3(n3833), .ZN(n3832) );
  AOI22_X1 U3445 ( .A1(n55), .A2(pc_ex_i[29]), .B1(pc_id_i[29]), .B2(n1079), 
        .ZN(n3831) );
  NAND2_X1 U3446 ( .A1(pc_if_i[29]), .A2(n1677), .ZN(n3830) );
  OAI21_X1 U3447 ( .B1(n1050), .B2(n3834), .A(n3835), .ZN(n4030) );
  AOI21_X1 U3448 ( .B1(pc_if_i[31]), .B2(n56), .A(n3836), .ZN(n3835) );
  NOR3_X1 U3449 ( .A1(n1054), .A2(n1677), .A3(n3837), .ZN(n3836) );
  NAND2_X1 U3450 ( .A1(n1385), .A2(hwlp_data_o[31]), .ZN(n3837) );
  AOI22_X1 U3451 ( .A1(pc_id_i[31]), .A2(n3838), .B1(pc_ex_i[31]), .B2(n3723), 
        .ZN(n3834) );
  INV_X1 U3452 ( .A(n1126), .ZN(n3838) );
  NAND3_X1 U3453 ( .A1(n3839), .A2(n1090), .A3(n1051), .ZN(n4033) );
  NAND2_X1 U3454 ( .A1(n56), .A2(pc_if_i[0]), .ZN(n3839) );
  NAND2_X1 U3455 ( .A1(n1127), .A2(n3840), .ZN(n4034) );
  NAND2_X1 U3456 ( .A1(pc_if_i[0]), .A2(n58), .ZN(n3840) );
  NAND2_X1 U3457 ( .A1(n1154), .A2(n3841), .ZN(n4035) );
  AOI22_X1 U3458 ( .A1(hwlp_data_o[11]), .A2(n3884), .B1(n1141), .B2(
        pc_ex_i[11]), .ZN(n3841) );
  NAND2_X1 U3459 ( .A1(n1140), .A2(n3842), .ZN(n4036) );
  AOI22_X1 U3460 ( .A1(hwlp_data_o[5]), .A2(n3884), .B1(pc_id_i[5]), .B2(n60), 
        .ZN(n3842) );
  OAI21_X1 U3461 ( .B1(n1125), .B2(n3843), .A(n3844), .ZN(n4037) );
  AOI22_X1 U3462 ( .A1(n1681), .A2(n3884), .B1(n60), .B2(pc_id_i[9]), .ZN(
        n3844) );
  AOI21_X1 U3463 ( .B1(pc_ex_i[9]), .B2(n3723), .A(n3845), .ZN(n3843) );
  AOI21_X1 U3464 ( .B1(n3890), .B2(n1124), .A(n3846), .ZN(n3845) );
  OAI21_X1 U3465 ( .B1(n3907), .B2(n3890), .A(pc_if_i[9]), .ZN(n3846) );
  AND2_X1 U3466 ( .A1(pc_if_i[9]), .A2(n3907), .ZN(n4038) );
  OAI21_X1 U3467 ( .B1(n1125), .B2(n3847), .A(n3848), .ZN(n4039) );
  AOI22_X1 U3468 ( .A1(n1682), .A2(n3894), .B1(n60), .B2(pc_id_i[10]), .ZN(
        n3848) );
  AOI21_X1 U3469 ( .B1(pc_if_i[10]), .B2(n3907), .A(n3849), .ZN(n3847) );
  AOI21_X1 U3470 ( .B1(n3890), .B2(csr_save_ex_i_BAR), .A(n3850), .ZN(n3849)
         );
  OAI21_X1 U3471 ( .B1(n3723), .B2(n3890), .A(pc_ex_i[10]), .ZN(n3850) );
  NAND2_X1 U3472 ( .A1(n1144), .A2(n3851), .ZN(n4040) );
  AOI22_X1 U3473 ( .A1(hwlp_data_o[6]), .A2(n1705), .B1(n58), .B2(pc_if_i[6]), 
        .ZN(n3851) );
  NAND2_X1 U3474 ( .A1(n1148), .A2(n3852), .ZN(n4041) );
  AOI22_X1 U3475 ( .A1(n4175), .A2(n1705), .B1(n58), .B2(pc_if_i[8]), .ZN(
        n3852) );
  NAND2_X1 U3476 ( .A1(n1132), .A2(n3853), .ZN(n4042) );
  AOI22_X1 U3477 ( .A1(hwlp_data_o[1]), .A2(n3894), .B1(pc_ex_i[1]), .B2(n1141), .ZN(n3853) );
  NAND2_X1 U3478 ( .A1(n1134), .A2(n3854), .ZN(n4043) );
  AOI22_X1 U3479 ( .A1(n4113), .A2(n1705), .B1(n1141), .B2(pc_ex_i[2]), .ZN(
        n3854) );
  OAI21_X1 U3480 ( .B1(n1125), .B2(n3855), .A(n3856), .ZN(n4044) );
  AOI22_X1 U3481 ( .A1(hwlp_data_o[4]), .A2(n1705), .B1(n60), .B2(pc_id_i[4]), 
        .ZN(n3856) );
  AOI21_X1 U3482 ( .B1(pc_ex_i[4]), .B2(n3723), .A(n3857), .ZN(n3855) );
  AOI21_X1 U3483 ( .B1(n3890), .B2(n1124), .A(n3858), .ZN(n3857) );
  OAI21_X1 U3484 ( .B1(n3907), .B2(n3890), .A(pc_if_i[4]), .ZN(n3858) );
  NAND2_X1 U3485 ( .A1(n1136), .A2(n3859), .ZN(n4045) );
  AOI22_X1 U3486 ( .A1(hwlp_data_o[3]), .A2(n1705), .B1(n1141), .B2(pc_ex_i[3]), .ZN(n3859) );
  OAI21_X1 U3487 ( .B1(n1125), .B2(n3860), .A(n3861), .ZN(n4046) );
  AOI22_X1 U3488 ( .A1(n4116), .A2(n1705), .B1(n60), .B2(pc_id_i[7]), .ZN(
        n3861) );
  AOI21_X1 U3489 ( .B1(pc_ex_i[7]), .B2(n3723), .A(n3862), .ZN(n3860) );
  AOI21_X1 U3490 ( .B1(n3890), .B2(n1124), .A(n3863), .ZN(n3862) );
  OAI21_X1 U3491 ( .B1(n3907), .B2(n3890), .A(pc_if_i[7]), .ZN(n3863) );
  AND2_X1 U3492 ( .A1(pc_if_i[7]), .A2(n3907), .ZN(n4047) );
  NAND2_X1 U3493 ( .A1(n1157), .A2(n3864), .ZN(n4048) );
  AOI22_X1 U3494 ( .A1(hwlp_data_o[12]), .A2(n3894), .B1(n1141), .B2(
        pc_ex_i[12]), .ZN(n3864) );
  NAND2_X1 U3495 ( .A1(n1159), .A2(n3865), .ZN(n4049) );
  AOI22_X1 U3496 ( .A1(n3960), .A2(n1705), .B1(n1141), .B2(pc_ex_i[13]), .ZN(
        n3865) );
  OAI211_X1 U3497 ( .C1(n1126), .C2(n3866), .A(n1161), .B(n3867), .ZN(n4050)
         );
  NAND2_X1 U3498 ( .A1(hwlp_data_o[14]), .A2(n3873), .ZN(n3867) );
  NAND2_X1 U3499 ( .A1(n1129), .A2(pc_id_i[14]), .ZN(n3866) );
  NAND2_X1 U3500 ( .A1(n1163), .A2(n3868), .ZN(n4051) );
  AOI22_X1 U3501 ( .A1(hwlp_data_o[15]), .A2(n1705), .B1(n58), .B2(pc_if_i[15]), .ZN(n3868) );
  NAND2_X1 U3502 ( .A1(n1170), .A2(n3869), .ZN(n4052) );
  AOI22_X1 U3503 ( .A1(n58), .A2(pc_if_i[18]), .B1(hwlp_data_o[18]), .B2(n3890), .ZN(n3869) );
  NAND2_X1 U3504 ( .A1(n1172), .A2(n3870), .ZN(n4053) );
  AOI22_X1 U3505 ( .A1(n1141), .A2(pc_ex_i[19]), .B1(hwlp_data_o[19]), .B2(
        n3890), .ZN(n3870) );
  OAI211_X1 U3506 ( .C1(n1126), .C2(n3871), .A(n1174), .B(n3872), .ZN(n4054)
         );
  NAND2_X1 U3507 ( .A1(n1678), .A2(n3873), .ZN(n3872) );
  NOR3_X1 U3508 ( .A1(n1198), .A2(n1129), .A3(n1130), .ZN(n3873) );
  NAND2_X1 U3509 ( .A1(n1129), .A2(pc_id_i[20]), .ZN(n3871) );
  OAI21_X1 U3510 ( .B1(n1125), .B2(n3874), .A(n3875), .ZN(n4055) );
  AOI22_X1 U3511 ( .A1(pc_id_i[21]), .A2(n60), .B1(n4183), .B2(n3890), .ZN(
        n3875) );
  AOI21_X1 U3512 ( .B1(pc_ex_i[21]), .B2(n3723), .A(n3876), .ZN(n3874) );
  AOI21_X1 U3513 ( .B1(n3890), .B2(n1124), .A(n3877), .ZN(n3876) );
  OAI21_X1 U3514 ( .B1(n3907), .B2(n3890), .A(pc_if_i[21]), .ZN(n3877) );
  NAND2_X1 U3515 ( .A1(n1178), .A2(n3878), .ZN(n4056) );
  AOI22_X1 U3516 ( .A1(hwlp_data_o[22]), .A2(n3894), .B1(pc_if_i[22]), .B2(n58), .ZN(n3878) );
  OAI21_X1 U3517 ( .B1(n1125), .B2(n3879), .A(n3880), .ZN(n4057) );
  AOI22_X1 U3518 ( .A1(n1141), .A2(pc_ex_i[23]), .B1(n3952), .B2(n3890), .ZN(
        n3880) );
  AOI22_X1 U3519 ( .A1(pc_id_i[23]), .A2(n3838), .B1(pc_if_i[23]), .B2(n3907), 
        .ZN(n3879) );
  NAND2_X1 U3520 ( .A1(n1185), .A2(n3881), .ZN(n4058) );
  AOI22_X1 U3521 ( .A1(n3954), .A2(n3884), .B1(pc_if_i[25]), .B2(n58), .ZN(
        n3881) );
  OAI21_X1 U3522 ( .B1(n1125), .B2(n3882), .A(n3883), .ZN(n4059) );
  AOI22_X1 U3523 ( .A1(n3955), .A2(n3884), .B1(n58), .B2(pc_if_i[26]), .ZN(
        n3883) );
  NOR3_X1 U3524 ( .A1(n1129), .A2(n1130), .A3(n1198), .ZN(n3884) );
  AOI21_X1 U3525 ( .B1(pc_id_i[26]), .B2(n3838), .A(n3885), .ZN(n3882) );
  AOI21_X1 U3526 ( .B1(n3890), .B2(csr_save_ex_i_BAR), .A(n3886), .ZN(n3885)
         );
  OAI21_X1 U3527 ( .B1(n3723), .B2(n3890), .A(pc_ex_i[26]), .ZN(n3886) );
  OAI21_X1 U3528 ( .B1(n1125), .B2(n3887), .A(n3888), .ZN(n4060) );
  AOI22_X1 U3529 ( .A1(n3956), .A2(n3894), .B1(n60), .B2(pc_id_i[27]), .ZN(
        n3888) );
  AOI21_X1 U3530 ( .B1(pc_if_i[27]), .B2(n3907), .A(n3889), .ZN(n3887) );
  AOI21_X1 U3531 ( .B1(n3890), .B2(csr_save_ex_i_BAR), .A(n3891), .ZN(n3889)
         );
  OAI21_X1 U3532 ( .B1(n3723), .B2(n3890), .A(pc_ex_i[27]), .ZN(n3891) );
  OAI21_X1 U3533 ( .B1(n1125), .B2(n3892), .A(n3893), .ZN(n4061) );
  AOI22_X1 U3534 ( .A1(hwlp_data_o[28]), .A2(n1705), .B1(n60), .B2(pc_id_i[28]), .ZN(n3893) );
  NOR3_X1 U3535 ( .A1(n1129), .A2(n1130), .A3(n1198), .ZN(n3894) );
  AOI21_X1 U3536 ( .B1(pc_if_i[28]), .B2(n3907), .A(n3895), .ZN(n3892) );
  AOI21_X1 U3537 ( .B1(n3890), .B2(csr_save_ex_i_BAR), .A(n3896), .ZN(n3895)
         );
  OAI21_X1 U3538 ( .B1(n3723), .B2(n3890), .A(pc_ex_i[28]), .ZN(n3896) );
  OAI21_X1 U3539 ( .B1(n1125), .B2(n3897), .A(n3898), .ZN(n4062) );
  AOI22_X1 U3540 ( .A1(n4143), .A2(n3899), .B1(n60), .B2(pc_id_i[29]), .ZN(
        n3898) );
  NOR3_X1 U3541 ( .A1(n1130), .A2(n1198), .A3(n1129), .ZN(n3899) );
  AOI22_X1 U3542 ( .A1(pc_if_i[29]), .A2(n3907), .B1(pc_ex_i[29]), .B2(n3723), 
        .ZN(n3897) );
  OAI21_X1 U3543 ( .B1(n1125), .B2(n3900), .A(n3901), .ZN(n4063) );
  AOI22_X1 U3544 ( .A1(n931), .A2(n1705), .B1(n60), .B2(pc_id_i[30]), .ZN(
        n3901) );
  AOI21_X1 U3545 ( .B1(pc_if_i[30]), .B2(n3907), .A(n3902), .ZN(n3900) );
  AOI21_X1 U3546 ( .B1(n3890), .B2(csr_save_ex_i_BAR), .A(n3903), .ZN(n3902)
         );
  OAI21_X1 U3547 ( .B1(n3723), .B2(n3890), .A(pc_ex_i[30]), .ZN(n3903) );
  OAI21_X1 U3548 ( .B1(n1125), .B2(n3904), .A(n3905), .ZN(n4064) );
  NAND2_X1 U3549 ( .A1(hwlp_data_o[31]), .A2(n3906), .ZN(n3905) );
  NOR3_X1 U3550 ( .A1(n1130), .A2(n1129), .A3(n1198), .ZN(n3906) );
  AOI222_X1 U3551 ( .A1(n3907), .A2(pc_if_i[31]), .B1(n3723), .B2(pc_ex_i[31]), 
        .C1(n3838), .C2(pc_id_i[31]), .ZN(n3904) );
  INV_X1 U3552 ( .A(n1124), .ZN(n3907) );
  NAND3_X1 U3553 ( .A1(n3908), .A2(n1166), .A3(n1127), .ZN(n4067) );
  NAND2_X1 U3554 ( .A1(n58), .A2(pc_if_i[0]), .ZN(n3908) );
  NOR2_X1 U3555 ( .A1(n1374), .A2(n1391), .ZN(n4068) );
  NOR2_X1 U3556 ( .A1(n1374), .A2(n1447), .ZN(n4069) );
  NOR2_X1 U3557 ( .A1(n1374), .A2(n1444), .ZN(n4070) );
  NOR2_X1 U3558 ( .A1(n1374), .A2(n1392), .ZN(n4071) );
  NOR2_X1 U3559 ( .A1(n1374), .A2(n1402), .ZN(n4072) );
  NOR2_X1 U3560 ( .A1(n1374), .A2(n1388), .ZN(n4073) );
  NOR2_X1 U3561 ( .A1(n1374), .A2(n1442), .ZN(n4074) );
  NOR2_X1 U3562 ( .A1(n1374), .A2(n1702), .ZN(n4075) );
  NOR2_X1 U3563 ( .A1(n1374), .A2(n1393), .ZN(n4076) );
  NOR2_X1 U3564 ( .A1(n1374), .A2(n1387), .ZN(n4077) );
  NOR2_X1 U3565 ( .A1(n1374), .A2(n1390), .ZN(n4078) );
  NOR2_X1 U3566 ( .A1(n1374), .A2(n1404), .ZN(n4079) );
  NOR2_X1 U3567 ( .A1(n1374), .A2(n1406), .ZN(n4080) );
  NOR2_X1 U3568 ( .A1(n1374), .A2(n1407), .ZN(n4081) );
  NOR2_X1 U3569 ( .A1(n1374), .A2(n1408), .ZN(n4082) );
  NOR2_X1 U3570 ( .A1(n1374), .A2(n1410), .ZN(n4083) );
  NOR2_X1 U3571 ( .A1(n1374), .A2(n68), .ZN(n4084) );
  NOR2_X1 U3572 ( .A1(n1374), .A2(n1411), .ZN(n4085) );
  NOR2_X1 U3573 ( .A1(n1374), .A2(n1412), .ZN(n4086) );
  NOR2_X1 U3574 ( .A1(n1374), .A2(n1700), .ZN(n4087) );
  NOR2_X1 U3575 ( .A1(n1374), .A2(n1414), .ZN(n4088) );
  NOR2_X1 U3576 ( .A1(n1374), .A2(n1415), .ZN(n4089) );
  NOR2_X1 U3577 ( .A1(n1374), .A2(n1416), .ZN(n4090) );
  NOR2_X1 U3578 ( .A1(n1374), .A2(n1418), .ZN(n4091) );
  NOR2_X1 U3579 ( .A1(n1374), .A2(n1704), .ZN(n4092) );
  NOR2_X1 U3580 ( .A1(n1374), .A2(n1421), .ZN(n4093) );
  NOR2_X1 U3581 ( .A1(n1374), .A2(n1422), .ZN(n4094) );
  NOR2_X1 U3582 ( .A1(n1374), .A2(n1423), .ZN(n4095) );
  NOR2_X1 U3583 ( .A1(n1374), .A2(n1426), .ZN(n4096) );
  AOI21_X1 U3584 ( .B1(n70), .B2(n3909), .A(n1377), .ZN(n4099) );
  INV_X1 U3585 ( .A(n4100), .ZN(n3909) );
  NOR2_X1 U3586 ( .A1(n1374), .A2(n1441), .ZN(n4100) );
  NOR2_X1 U3587 ( .A1(n1706), .A2(n1391), .ZN(n4103) );
  INV_X1 U3588 ( .A(n1391), .ZN(hwlp_data_o[5]) );
  NOR2_X1 U3589 ( .A1(n1706), .A2(n1447), .ZN(n4105) );
  NOR2_X1 U3590 ( .A1(n1706), .A2(n1444), .ZN(n4106) );
  NOR2_X1 U3591 ( .A1(n1706), .A2(n1392), .ZN(n4107) );
  INV_X1 U3592 ( .A(n1392), .ZN(hwlp_data_o[6]) );
  NOR2_X1 U3593 ( .A1(n1706), .A2(n1402), .ZN(n4109) );
  NOR2_X1 U3594 ( .A1(n1706), .A2(n1388), .ZN(n4110) );
  INV_X1 U3595 ( .A(n1388), .ZN(hwlp_data_o[1]) );
  NOR2_X1 U3596 ( .A1(n1706), .A2(n1442), .ZN(n4112) );
  INV_X1 U3597 ( .A(n1442), .ZN(n4113) );
  NOR2_X1 U3598 ( .A1(n1706), .A2(n1702), .ZN(n4114) );
  NOR2_X1 U3599 ( .A1(n1706), .A2(n1393), .ZN(n4115) );
  INV_X1 U3600 ( .A(n1393), .ZN(n4116) );
  NOR2_X1 U3601 ( .A1(n1706), .A2(n1387), .ZN(n4117) );
  INV_X1 U3602 ( .A(n1387), .ZN(hwlp_data_o[0]) );
  NOR2_X1 U3603 ( .A1(n1706), .A2(n1390), .ZN(n4119) );
  NOR2_X1 U3604 ( .A1(n1706), .A2(n1404), .ZN(n4120) );
  NOR2_X1 U3605 ( .A1(n1706), .A2(n1405), .ZN(n4121) );
  NOR2_X1 U3606 ( .A1(n1706), .A2(n1406), .ZN(n4122) );
  NOR2_X1 U3607 ( .A1(n1706), .A2(n1407), .ZN(n4123) );
  INV_X1 U3608 ( .A(n1407), .ZN(hwlp_data_o[14]) );
  NOR2_X1 U3609 ( .A1(n1706), .A2(n1408), .ZN(n4125) );
  INV_X1 U3610 ( .A(n1408), .ZN(hwlp_data_o[15]) );
  NOR2_X1 U3611 ( .A1(n1706), .A2(n1409), .ZN(n4127) );
  NOR2_X1 U3612 ( .A1(n1706), .A2(n1410), .ZN(n4128) );
  INV_X1 U3613 ( .A(n1410), .ZN(hwlp_data_o[17]) );
  NOR2_X1 U3614 ( .A1(n1706), .A2(n68), .ZN(n4130) );
  INV_X1 U3615 ( .A(n68), .ZN(hwlp_data_o[18]) );
  NOR2_X1 U3616 ( .A1(n1706), .A2(n1411), .ZN(n4132) );
  NOR2_X1 U3617 ( .A1(n1706), .A2(n1412), .ZN(n4133) );
  NOR2_X1 U3618 ( .A1(n1706), .A2(n1700), .ZN(n4134) );
  NOR2_X1 U3619 ( .A1(n1706), .A2(n1414), .ZN(n4135) );
  NOR2_X1 U3620 ( .A1(n1706), .A2(n1415), .ZN(n4136) );
  NOR2_X1 U3621 ( .A1(n1706), .A2(n1416), .ZN(n4137) );
  NOR2_X1 U3622 ( .A1(n1706), .A2(n1418), .ZN(n4138) );
  NOR2_X1 U3623 ( .A1(n1706), .A2(n1704), .ZN(n4139) );
  NOR2_X1 U3624 ( .A1(n1706), .A2(n1421), .ZN(n4140) );
  NOR2_X1 U3625 ( .A1(n1706), .A2(n1422), .ZN(n4141) );
  NOR2_X1 U3626 ( .A1(n1706), .A2(n1423), .ZN(n4142) );
  INV_X1 U3627 ( .A(n1423), .ZN(n4143) );
  NOR2_X1 U3628 ( .A1(n1706), .A2(n1426), .ZN(n4144) );
  AOI21_X1 U3629 ( .B1(n70), .B2(n3910), .A(n1382), .ZN(n4147) );
  INV_X1 U3630 ( .A(n4148), .ZN(n3910) );
  NOR2_X1 U3631 ( .A1(n1706), .A2(n1441), .ZN(n4148) );
  INV_X1 U3640 ( .A(n1409), .ZN(hwlp_data_o[16]) );
  INV_X1 U3642 ( .A(n1406), .ZN(n3960) );
  INV_X1 U3645 ( .A(n865), .ZN(n3966) );
  INV_X1 U3647 ( .A(n1446), .ZN(n3969) );
endmodule


module riscv_load_store_unit ( clk, rst_n, data_req_o, data_gnt_i, 
        data_rvalid_i, data_addr_o, data_we_o, data_be_o, data_wdata_o, 
        data_rdata_i, data_we_ex_i, data_type_ex_i, data_wdata_ex_i, 
        data_reg_offset_ex_i, data_sign_ext_ex_i, data_rdata_ex_o, 
        data_req_ex_i, operand_a_ex_i, operand_b_ex_i, data_misaligned_o, 
        lsu_ready_ex_o, lsu_ready_wb_o, ex_valid_i, busy_o, data_err_i_BAR, 
        data_misaligned_ex_i_BAR, addr_useincr_ex_i );
  output [31:0] data_addr_o;
  output [3:0] data_be_o;
  output [31:0] data_wdata_o;
  input [31:0] data_rdata_i;
  input [1:0] data_type_ex_i;
  input [31:0] data_wdata_ex_i;
  input [1:0] data_reg_offset_ex_i;
  input [1:0] data_sign_ext_ex_i;
  output [31:0] data_rdata_ex_o;
  input [31:0] operand_a_ex_i;
  input [31:0] operand_b_ex_i;
  input clk, rst_n, data_gnt_i, data_rvalid_i, data_we_ex_i, data_req_ex_i,
         ex_valid_i, data_err_i_BAR, data_misaligned_ex_i_BAR,
         addr_useincr_ex_i;
  output data_req_o, data_we_o, data_misaligned_o, lsu_ready_ex_o,
         lsu_ready_wb_o, busy_o;
  wire   data_we_ex_i, data_misaligned_ex_i, data_sign_ext_q_0_, n429, n430,
         n2, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n423, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n586, n587, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n633, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n713, n715, n717, n719, n721, n723, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908;
  wire   [1:0] data_type_q;
  wire   [1:0] rdata_offset_q;
  wire   [31:0] rdata_q;
  wire   [1:0] CS;
  assign data_we_o = data_we_ex_i;
  assign data_misaligned_ex_i = data_misaligned_ex_i_BAR;

  AND2_X4 U4 ( .A1(n8), .A2(n7), .ZN(n263) );
  XNOR2_X1 U7 ( .A(n146), .B(operand_a_ex_i[1]), .ZN(n2) );
  CLKBUF_X1 U11 ( .A(data_gnt_i), .Z(n584) );
  MUX2_X2 U12 ( .A(rdata_q[22]), .B(n537), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[22]) );
  MUX2_X2 U13 ( .A(rdata_q[23]), .B(n476), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[23]) );
  MUX2_X2 U14 ( .A(rdata_q[20]), .B(n473), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[20]) );
  MUX2_X2 U15 ( .A(rdata_q[14]), .B(n534), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[14]) );
  MUX2_X2 U16 ( .A(rdata_q[12]), .B(n481), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[12]) );
  MUX2_X2 U17 ( .A(rdata_q[11]), .B(n451), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[11]) );
  MUX2_X2 U18 ( .A(rdata_q[13]), .B(n489), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[13]) );
  MUX2_X2 U19 ( .A(rdata_q[9]), .B(n465), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[9]) );
  MUX2_X2 U20 ( .A(rdata_q[10]), .B(n500), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[10]) );
  MUX2_X2 U21 ( .A(rdata_q[8]), .B(n470), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[8]) );
  AOI21_X2 U22 ( .B1(n573), .B2(n572), .A(n571), .ZN(data_misaligned_o) );
  OR2_X1 U23 ( .A1(n11), .A2(n12), .ZN(n9) );
  OAI21_X1 U24 ( .B1(n45), .B2(n34), .A(n33), .ZN(n86) );
  INV_X1 U25 ( .A(data_type_ex_i[0]), .ZN(n569) );
  NOR2_X1 U26 ( .A1(n774), .A2(data_type_ex_i[1]), .ZN(n570) );
  OR2_X1 U27 ( .A1(data_gnt_i), .A2(n9), .ZN(lsu_ready_ex_o) );
  INV_X1 U28 ( .A(n84), .ZN(n8) );
  NAND2_X1 U29 ( .A1(n570), .A2(data_req_ex_i), .ZN(n571) );
  NAND2_X1 U30 ( .A1(data_addr_o[0]), .A2(n569), .ZN(n572) );
  INV_X2 U32 ( .A(n444), .ZN(data_rdata_ex_o[2]) );
  INV_X2 U33 ( .A(n431), .ZN(data_rdata_ex_o[4]) );
  INV_X2 U34 ( .A(n357), .ZN(data_rdata_ex_o[3]) );
  INV_X2 U35 ( .A(n436), .ZN(data_rdata_ex_o[5]) );
  INV_X2 U36 ( .A(n367), .ZN(data_rdata_ex_o[0]) );
  INV_X2 U37 ( .A(n362), .ZN(data_rdata_ex_o[6]) );
  INV_X2 U38 ( .A(n460), .ZN(data_rdata_ex_o[1]) );
  NAND2_X2 U39 ( .A1(n5), .A2(n6), .ZN(data_rdata_ex_o[19]) );
  NAND2_X1 U40 ( .A1(data_rvalid_i), .A2(n492), .ZN(n5) );
  NAND2_X1 U41 ( .A1(rdata_q[19]), .A2(n459), .ZN(n6) );
  NAND2_X1 U42 ( .A1(n85), .A2(n86), .ZN(n7) );
  NOR2_X1 U43 ( .A1(data_type_q[1]), .A2(data_type_q[0]), .ZN(n509) );
  NOR2_X1 U45 ( .A1(n770), .A2(n16), .ZN(n152) );
  OR2_X1 U46 ( .A1(data_addr_o[0]), .A2(n569), .ZN(n568) );
  XNOR2_X1 U47 ( .A(n152), .B(operand_a_ex_i[0]), .ZN(n153) );
  XOR2_X1 U48 ( .A(n147), .B(n2), .Z(data_addr_o[1]) );
  NOR2_X1 U49 ( .A1(CS[1]), .A2(CS[0]), .ZN(n637) );
  AND2_X1 U50 ( .A1(n637), .A2(data_req_ex_i), .ZN(n10) );
  OR2_X1 U51 ( .A1(n576), .A2(n10), .ZN(data_req_o) );
  INV_X1 U52 ( .A(data_err_i_BAR), .ZN(n12) );
  INV_X1 U53 ( .A(data_req_o), .ZN(n11) );
  INV_X1 U54 ( .A(operand_b_ex_i[2]), .ZN(n13) );
  NOR2_X1 U55 ( .A1(n770), .A2(n13), .ZN(n19) );
  NOR2_X1 U56 ( .A1(n19), .A2(operand_a_ex_i[2]), .ZN(n62) );
  INV_X1 U57 ( .A(operand_b_ex_i[3]), .ZN(n14) );
  NOR2_X1 U58 ( .A1(n769), .A2(n14), .ZN(n20) );
  NOR2_X1 U60 ( .A1(n62), .A2(n57), .ZN(n22) );
  INV_X1 U61 ( .A(operand_b_ex_i[1]), .ZN(n15) );
  NOR2_X1 U62 ( .A1(n770), .A2(n15), .ZN(n146) );
  NOR2_X1 U63 ( .A1(n146), .A2(operand_a_ex_i[1]), .ZN(n18) );
  INV_X1 U64 ( .A(operand_b_ex_i[0]), .ZN(n16) );
  NAND2_X1 U65 ( .A1(n152), .A2(operand_a_ex_i[0]), .ZN(n147) );
  NAND2_X1 U66 ( .A1(n146), .A2(operand_a_ex_i[1]), .ZN(n17) );
  OAI21_X1 U67 ( .B1(n18), .B2(n147), .A(n17), .ZN(n56) );
  NAND2_X1 U68 ( .A1(n19), .A2(operand_a_ex_i[2]), .ZN(n63) );
  NAND2_X1 U69 ( .A1(n20), .A2(operand_a_ex_i[3]), .ZN(n58) );
  OAI21_X1 U70 ( .B1(n57), .B2(n63), .A(n58), .ZN(n21) );
  AOI21_X1 U71 ( .B1(n22), .B2(n56), .A(n21), .ZN(n45) );
  INV_X1 U72 ( .A(operand_b_ex_i[4]), .ZN(n23) );
  NOR2_X1 U73 ( .A1(n770), .A2(n23), .ZN(n27) );
  NOR2_X1 U74 ( .A1(n27), .A2(operand_a_ex_i[4]), .ZN(n46) );
  INV_X1 U75 ( .A(operand_b_ex_i[5]), .ZN(n24) );
  NOR2_X1 U76 ( .A1(n768), .A2(n24), .ZN(n28) );
  NOR2_X1 U78 ( .A1(n46), .A2(n48), .ZN(n235) );
  INV_X1 U79 ( .A(operand_b_ex_i[6]), .ZN(n25) );
  NOR2_X1 U80 ( .A1(n770), .A2(n25), .ZN(n29) );
  INV_X1 U82 ( .A(operand_b_ex_i[7]), .ZN(n26) );
  NOR2_X1 U83 ( .A1(n770), .A2(n26), .ZN(n30) );
  NOR2_X1 U84 ( .A1(n30), .A2(operand_a_ex_i[7]), .ZN(n229) );
  NOR2_X1 U85 ( .A1(n237), .A2(n229), .ZN(n32) );
  NAND2_X1 U86 ( .A1(n235), .A2(n32), .ZN(n34) );
  NAND2_X1 U87 ( .A1(n27), .A2(operand_a_ex_i[4]), .ZN(n53) );
  NAND2_X1 U88 ( .A1(n28), .A2(operand_a_ex_i[5]), .ZN(n49) );
  OAI21_X1 U89 ( .B1(n48), .B2(n53), .A(n49), .ZN(n234) );
  NAND2_X1 U90 ( .A1(n29), .A2(operand_a_ex_i[6]), .ZN(n238) );
  NAND2_X1 U91 ( .A1(n30), .A2(operand_a_ex_i[7]), .ZN(n230) );
  OAI21_X1 U92 ( .B1(n229), .B2(n238), .A(n230), .ZN(n31) );
  AOI21_X1 U93 ( .B1(n32), .B2(n234), .A(n31), .ZN(n33) );
  INV_X1 U94 ( .A(n86), .ZN(n299) );
  INV_X1 U95 ( .A(operand_b_ex_i[8]), .ZN(n35) );
  NOR2_X1 U96 ( .A1(n770), .A2(n35), .ZN(n37) );
  NOR2_X1 U97 ( .A1(n37), .A2(operand_a_ex_i[8]), .ZN(n255) );
  INV_X1 U98 ( .A(operand_b_ex_i[9]), .ZN(n36) );
  NOR2_X1 U99 ( .A1(n769), .A2(n36), .ZN(n38) );
  NOR2_X1 U100 ( .A1(n255), .A2(n256), .ZN(n242) );
  INV_X1 U101 ( .A(n242), .ZN(n40) );
  NAND2_X1 U102 ( .A1(n37), .A2(operand_a_ex_i[8]), .ZN(n254) );
  NAND2_X1 U103 ( .A1(n38), .A2(operand_a_ex_i[9]), .ZN(n257) );
  OAI21_X1 U104 ( .B1(n256), .B2(n254), .A(n257), .ZN(n246) );
  INV_X1 U105 ( .A(n246), .ZN(n39) );
  OAI21_X1 U106 ( .B1(n299), .B2(n40), .A(n39), .ZN(n44) );
  INV_X1 U107 ( .A(operand_b_ex_i[10]), .ZN(n41) );
  NOR2_X1 U108 ( .A1(n769), .A2(n41), .ZN(n42) );
  NOR2_X1 U109 ( .A1(n42), .A2(operand_a_ex_i[10]), .ZN(n68) );
  INV_X1 U110 ( .A(n68), .ZN(n245) );
  NAND2_X1 U111 ( .A1(n42), .A2(operand_a_ex_i[10]), .ZN(n243) );
  NAND2_X1 U112 ( .A1(n245), .A2(n243), .ZN(n43) );
  XNOR2_X1 U113 ( .A(n44), .B(n43), .ZN(data_addr_o[10]) );
  INV_X1 U114 ( .A(n45), .ZN(n236) );
  INV_X1 U115 ( .A(n46), .ZN(n54) );
  INV_X1 U116 ( .A(n53), .ZN(n47) );
  AOI21_X1 U117 ( .B1(n236), .B2(n54), .A(n47), .ZN(n52) );
  INV_X1 U118 ( .A(n48), .ZN(n50) );
  NAND2_X1 U119 ( .A1(n50), .A2(n49), .ZN(n51) );
  XOR2_X1 U120 ( .A(n52), .B(n51), .Z(data_addr_o[5]) );
  NAND2_X1 U121 ( .A1(n54), .A2(n53), .ZN(n55) );
  XNOR2_X1 U122 ( .A(n236), .B(n55), .ZN(data_addr_o[4]) );
  INV_X1 U123 ( .A(n56), .ZN(n66) );
  OAI21_X1 U124 ( .B1(n66), .B2(n62), .A(n63), .ZN(n61) );
  INV_X1 U125 ( .A(n57), .ZN(n59) );
  NAND2_X1 U126 ( .A1(n59), .A2(n58), .ZN(n60) );
  XNOR2_X1 U127 ( .A(n61), .B(n60), .ZN(data_addr_o[3]) );
  INV_X1 U128 ( .A(n62), .ZN(n64) );
  NAND2_X1 U129 ( .A1(n64), .A2(n63), .ZN(n65) );
  XOR2_X1 U130 ( .A(n66), .B(n65), .Z(data_addr_o[2]) );
  INV_X1 U131 ( .A(operand_b_ex_i[11]), .ZN(n67) );
  NOR2_X1 U132 ( .A1(n769), .A2(n67), .ZN(n73) );
  NOR2_X1 U134 ( .A1(n68), .A2(n249), .ZN(n75) );
  NAND2_X1 U135 ( .A1(n242), .A2(n75), .ZN(n271) );
  INV_X1 U136 ( .A(operand_b_ex_i[12]), .ZN(n69) );
  NOR2_X1 U137 ( .A1(n770), .A2(n69), .ZN(n76) );
  NOR2_X1 U138 ( .A1(n76), .A2(operand_a_ex_i[12]), .ZN(n268) );
  INV_X1 U139 ( .A(operand_b_ex_i[13]), .ZN(n70) );
  NOR2_X1 U140 ( .A1(n768), .A2(n70), .ZN(n77) );
  NOR2_X1 U141 ( .A1(n77), .A2(operand_a_ex_i[13]), .ZN(n277) );
  INV_X1 U143 ( .A(operand_b_ex_i[14]), .ZN(n71) );
  NOR2_X1 U144 ( .A1(n770), .A2(n71), .ZN(n78) );
  NOR2_X1 U145 ( .A1(n78), .A2(operand_a_ex_i[14]), .ZN(n292) );
  INV_X1 U146 ( .A(operand_b_ex_i[15]), .ZN(n72) );
  NOR2_X1 U147 ( .A1(n770), .A2(n72), .ZN(n79) );
  NOR2_X1 U148 ( .A1(n79), .A2(operand_a_ex_i[15]), .ZN(n300) );
  NOR2_X1 U149 ( .A1(n292), .A2(n300), .ZN(n81) );
  NAND2_X1 U150 ( .A1(n287), .A2(n81), .ZN(n83) );
  NOR2_X1 U151 ( .A1(n271), .A2(n83), .ZN(n85) );
  NAND2_X1 U152 ( .A1(n73), .A2(operand_a_ex_i[11]), .ZN(n250) );
  OAI21_X1 U153 ( .B1(n249), .B2(n243), .A(n250), .ZN(n74) );
  AOI21_X1 U154 ( .B1(n75), .B2(n246), .A(n74), .ZN(n267) );
  NAND2_X1 U155 ( .A1(n76), .A2(operand_a_ex_i[12]), .ZN(n272) );
  NAND2_X1 U156 ( .A1(n77), .A2(operand_a_ex_i[13]), .ZN(n278) );
  OAI21_X1 U157 ( .B1(n277), .B2(n272), .A(n278), .ZN(n290) );
  NAND2_X1 U158 ( .A1(n78), .A2(operand_a_ex_i[14]), .ZN(n291) );
  NAND2_X1 U159 ( .A1(n79), .A2(operand_a_ex_i[15]), .ZN(n301) );
  OAI21_X1 U160 ( .B1(n300), .B2(n291), .A(n301), .ZN(n80) );
  AOI21_X1 U161 ( .B1(n81), .B2(n290), .A(n80), .ZN(n82) );
  OAI21_X1 U162 ( .B1(n267), .B2(n83), .A(n82), .ZN(n84) );
  INV_X1 U163 ( .A(operand_b_ex_i[16]), .ZN(n87) );
  NOR2_X1 U164 ( .A1(n768), .A2(n87), .ZN(n88) );
  NOR2_X1 U165 ( .A1(n88), .A2(operand_a_ex_i[16]), .ZN(n148) );
  NAND2_X1 U166 ( .A1(n88), .A2(operand_a_ex_i[16]), .ZN(n149) );
  OAI21_X1 U167 ( .B1(n263), .B2(n148), .A(n149), .ZN(n93) );
  INV_X1 U168 ( .A(operand_b_ex_i[17]), .ZN(n89) );
  NOR2_X1 U169 ( .A1(n768), .A2(n89), .ZN(n90) );
  NOR2_X1 U170 ( .A1(n90), .A2(operand_a_ex_i[17]), .ZN(n109) );
  INV_X1 U171 ( .A(n109), .ZN(n91) );
  NAND2_X1 U172 ( .A1(n90), .A2(operand_a_ex_i[17]), .ZN(n108) );
  NAND2_X1 U173 ( .A1(n91), .A2(n108), .ZN(n92) );
  XNOR2_X1 U174 ( .A(n93), .B(n92), .ZN(data_addr_o[17]) );
  NOR2_X1 U175 ( .A1(n148), .A2(n109), .ZN(n202) );
  INV_X1 U176 ( .A(operand_b_ex_i[18]), .ZN(n94) );
  NOR2_X1 U177 ( .A1(n770), .A2(n94), .ZN(n110) );
  NOR2_X1 U178 ( .A1(n110), .A2(operand_a_ex_i[18]), .ZN(n183) );
  INV_X1 U179 ( .A(operand_b_ex_i[19]), .ZN(n95) );
  NOR2_X1 U180 ( .A1(n770), .A2(n95), .ZN(n111) );
  NOR2_X1 U181 ( .A1(n111), .A2(operand_a_ex_i[19]), .ZN(n187) );
  NOR2_X1 U182 ( .A1(n183), .A2(n187), .ZN(n113) );
  NAND2_X1 U183 ( .A1(n202), .A2(n113), .ZN(n262) );
  INV_X1 U184 ( .A(operand_b_ex_i[20]), .ZN(n96) );
  NOR2_X1 U185 ( .A1(n768), .A2(n96), .ZN(n114) );
  NOR2_X1 U186 ( .A1(n114), .A2(operand_a_ex_i[20]), .ZN(n264) );
  INV_X1 U187 ( .A(operand_b_ex_i[21]), .ZN(n97) );
  NOR2_X1 U188 ( .A1(n768), .A2(n97), .ZN(n115) );
  NOR2_X1 U189 ( .A1(n115), .A2(operand_a_ex_i[21]), .ZN(n312) );
  NOR2_X1 U190 ( .A1(n264), .A2(n312), .ZN(n210) );
  INV_X1 U191 ( .A(operand_b_ex_i[22]), .ZN(n98) );
  NOR2_X1 U192 ( .A1(n770), .A2(n98), .ZN(n116) );
  NOR2_X1 U193 ( .A1(n116), .A2(operand_a_ex_i[22]), .ZN(n214) );
  INV_X1 U194 ( .A(operand_b_ex_i[23]), .ZN(n99) );
  NOR2_X1 U195 ( .A1(n770), .A2(n99), .ZN(n117) );
  NOR2_X1 U196 ( .A1(n117), .A2(operand_a_ex_i[23]), .ZN(n220) );
  NOR2_X1 U197 ( .A1(n214), .A2(n220), .ZN(n119) );
  NAND2_X1 U198 ( .A1(n210), .A2(n119), .ZN(n121) );
  INV_X1 U200 ( .A(operand_b_ex_i[24]), .ZN(n101) );
  NOR2_X1 U201 ( .A1(n769), .A2(n101), .ZN(n122) );
  NOR2_X1 U202 ( .A1(n122), .A2(operand_a_ex_i[24]), .ZN(n180) );
  INV_X1 U203 ( .A(operand_b_ex_i[25]), .ZN(n102) );
  NOR2_X1 U204 ( .A1(n770), .A2(n102), .ZN(n123) );
  NOR2_X1 U205 ( .A1(n123), .A2(operand_a_ex_i[25]), .ZN(n197) );
  NOR2_X1 U206 ( .A1(n180), .A2(n197), .ZN(n322) );
  INV_X1 U207 ( .A(operand_b_ex_i[26]), .ZN(n103) );
  NOR2_X1 U208 ( .A1(n769), .A2(n103), .ZN(n124) );
  NOR2_X1 U209 ( .A1(n124), .A2(operand_a_ex_i[26]), .ZN(n326) );
  INV_X1 U210 ( .A(operand_b_ex_i[27]), .ZN(n104) );
  NOR2_X1 U211 ( .A1(n770), .A2(n104), .ZN(n125) );
  NOR2_X1 U212 ( .A1(n125), .A2(operand_a_ex_i[27]), .ZN(n332) );
  NOR2_X1 U213 ( .A1(n326), .A2(n332), .ZN(n127) );
  NAND2_X1 U214 ( .A1(n322), .A2(n127), .ZN(n337) );
  INV_X1 U215 ( .A(operand_b_ex_i[28]), .ZN(n105) );
  NOR2_X1 U216 ( .A1(n770), .A2(n105), .ZN(n128) );
  NOR2_X1 U217 ( .A1(n128), .A2(operand_a_ex_i[28]), .ZN(n340) );
  INV_X1 U218 ( .A(operand_b_ex_i[29]), .ZN(n106) );
  NOR2_X1 U219 ( .A1(n769), .A2(n106), .ZN(n129) );
  NOR2_X1 U220 ( .A1(n129), .A2(operand_a_ex_i[29]), .ZN(n347) );
  NOR2_X1 U221 ( .A1(n340), .A2(n347), .ZN(n161) );
  INV_X1 U222 ( .A(operand_b_ex_i[30]), .ZN(n107) );
  NOR2_X1 U223 ( .A1(n770), .A2(n107), .ZN(n130) );
  OR2_X1 U224 ( .A1(n130), .A2(operand_a_ex_i[30]), .ZN(n170) );
  NAND2_X1 U225 ( .A1(n161), .A2(n170), .ZN(n133) );
  NOR2_X1 U226 ( .A1(n337), .A2(n133), .ZN(n135) );
  NAND2_X1 U227 ( .A1(n338), .A2(n135), .ZN(n137) );
  OAI21_X1 U228 ( .B1(n109), .B2(n149), .A(n108), .ZN(n203) );
  NAND2_X1 U229 ( .A1(n110), .A2(operand_a_ex_i[18]), .ZN(n206) );
  NAND2_X1 U230 ( .A1(n111), .A2(operand_a_ex_i[19]), .ZN(n188) );
  OAI21_X1 U231 ( .B1(n187), .B2(n206), .A(n188), .ZN(n112) );
  AOI21_X1 U232 ( .B1(n113), .B2(n203), .A(n112), .ZN(n261) );
  NAND2_X1 U233 ( .A1(n114), .A2(operand_a_ex_i[20]), .ZN(n306) );
  NAND2_X1 U234 ( .A1(n115), .A2(operand_a_ex_i[21]), .ZN(n313) );
  OAI21_X1 U235 ( .B1(n312), .B2(n306), .A(n313), .ZN(n212) );
  NAND2_X1 U236 ( .A1(n116), .A2(operand_a_ex_i[22]), .ZN(n213) );
  NAND2_X1 U237 ( .A1(n117), .A2(operand_a_ex_i[23]), .ZN(n221) );
  OAI21_X1 U238 ( .B1(n220), .B2(n213), .A(n221), .ZN(n118) );
  AOI21_X1 U239 ( .B1(n119), .B2(n212), .A(n118), .ZN(n120) );
  NAND2_X1 U241 ( .A1(n122), .A2(operand_a_ex_i[24]), .ZN(n192) );
  NAND2_X1 U242 ( .A1(n123), .A2(operand_a_ex_i[25]), .ZN(n198) );
  OAI21_X1 U243 ( .B1(n197), .B2(n192), .A(n198), .ZN(n324) );
  NAND2_X1 U244 ( .A1(n124), .A2(operand_a_ex_i[26]), .ZN(n325) );
  NAND2_X1 U245 ( .A1(n125), .A2(operand_a_ex_i[27]), .ZN(n333) );
  OAI21_X1 U246 ( .B1(n332), .B2(n325), .A(n333), .ZN(n126) );
  AOI21_X1 U247 ( .B1(n127), .B2(n324), .A(n126), .ZN(n341) );
  NAND2_X1 U248 ( .A1(n128), .A2(operand_a_ex_i[28]), .ZN(n339) );
  NAND2_X1 U249 ( .A1(n129), .A2(operand_a_ex_i[29]), .ZN(n348) );
  OAI21_X1 U250 ( .B1(n347), .B2(n339), .A(n348), .ZN(n162) );
  NAND2_X1 U251 ( .A1(n130), .A2(operand_a_ex_i[30]), .ZN(n169) );
  INV_X1 U252 ( .A(n169), .ZN(n131) );
  AOI21_X1 U253 ( .B1(n162), .B2(n170), .A(n131), .ZN(n132) );
  OAI21_X1 U254 ( .B1(n341), .B2(n133), .A(n132), .ZN(n134) );
  AOI21_X1 U255 ( .B1(n135), .B2(n344), .A(n134), .ZN(n136) );
  OAI21_X1 U256 ( .B1(n263), .B2(n137), .A(n136), .ZN(n143) );
  INV_X1 U257 ( .A(operand_b_ex_i[31]), .ZN(n138) );
  NOR2_X1 U258 ( .A1(n769), .A2(n138), .ZN(n139) );
  OR2_X1 U259 ( .A1(n139), .A2(operand_a_ex_i[31]), .ZN(n141) );
  NAND2_X1 U260 ( .A1(n139), .A2(operand_a_ex_i[31]), .ZN(n140) );
  NAND2_X1 U261 ( .A1(n141), .A2(n140), .ZN(n142) );
  XNOR2_X1 U262 ( .A(n143), .B(n142), .ZN(data_addr_o[31]) );
  INV_X1 U263 ( .A(n255), .ZN(n144) );
  NAND2_X1 U264 ( .A1(n144), .A2(n254), .ZN(n145) );
  XOR2_X1 U265 ( .A(n299), .B(n145), .Z(data_addr_o[8]) );
  INV_X1 U266 ( .A(n148), .ZN(n150) );
  NAND2_X1 U267 ( .A1(n150), .A2(n149), .ZN(n151) );
  XOR2_X1 U268 ( .A(n263), .B(n151), .Z(data_addr_o[16]) );
  INV_X1 U269 ( .A(n153), .ZN(data_addr_o[0]) );
  INV_X1 U270 ( .A(n337), .ZN(n155) );
  NAND2_X1 U271 ( .A1(n338), .A2(n155), .ZN(n157) );
  INV_X1 U272 ( .A(n341), .ZN(n154) );
  AOI21_X1 U273 ( .B1(n344), .B2(n155), .A(n154), .ZN(n156) );
  OAI21_X1 U274 ( .B1(n263), .B2(n157), .A(n156), .ZN(n160) );
  INV_X1 U275 ( .A(n340), .ZN(n158) );
  NAND2_X1 U276 ( .A1(n158), .A2(n339), .ZN(n159) );
  XNOR2_X1 U277 ( .A(n160), .B(n159), .ZN(data_addr_o[28]) );
  INV_X1 U278 ( .A(n161), .ZN(n164) );
  NOR2_X1 U279 ( .A1(n337), .A2(n164), .ZN(n166) );
  NAND2_X1 U280 ( .A1(n338), .A2(n166), .ZN(n168) );
  INV_X1 U281 ( .A(n162), .ZN(n163) );
  OAI21_X1 U282 ( .B1(n341), .B2(n164), .A(n163), .ZN(n165) );
  AOI21_X1 U283 ( .B1(n344), .B2(n166), .A(n165), .ZN(n167) );
  OAI21_X1 U284 ( .B1(n263), .B2(n168), .A(n167), .ZN(n172) );
  NAND2_X1 U285 ( .A1(n170), .A2(n169), .ZN(n171) );
  XNOR2_X1 U286 ( .A(n172), .B(n171), .ZN(data_addr_o[30]) );
  INV_X1 U287 ( .A(n262), .ZN(n305) );
  NAND2_X1 U288 ( .A1(n305), .A2(n210), .ZN(n174) );
  INV_X1 U289 ( .A(n261), .ZN(n309) );
  AOI21_X1 U290 ( .B1(n309), .B2(n210), .A(n212), .ZN(n173) );
  OAI21_X1 U291 ( .B1(n263), .B2(n174), .A(n173), .ZN(n177) );
  INV_X1 U292 ( .A(n214), .ZN(n175) );
  NAND2_X1 U293 ( .A1(n175), .A2(n213), .ZN(n176) );
  XNOR2_X1 U294 ( .A(n177), .B(n176), .ZN(data_addr_o[22]) );
  INV_X1 U295 ( .A(n338), .ZN(n179) );
  INV_X1 U296 ( .A(n344), .ZN(n178) );
  OAI21_X1 U297 ( .B1(n263), .B2(n179), .A(n178), .ZN(n182) );
  INV_X1 U298 ( .A(n180), .ZN(n194) );
  NAND2_X1 U299 ( .A1(n194), .A2(n192), .ZN(n181) );
  XNOR2_X1 U300 ( .A(n182), .B(n181), .ZN(data_addr_o[24]) );
  INV_X1 U301 ( .A(n183), .ZN(n207) );
  NAND2_X1 U302 ( .A1(n202), .A2(n207), .ZN(n186) );
  INV_X1 U303 ( .A(n206), .ZN(n184) );
  AOI21_X1 U304 ( .B1(n203), .B2(n207), .A(n184), .ZN(n185) );
  OAI21_X1 U305 ( .B1(n263), .B2(n186), .A(n185), .ZN(n191) );
  INV_X1 U306 ( .A(n187), .ZN(n189) );
  NAND2_X1 U307 ( .A1(n189), .A2(n188), .ZN(n190) );
  XNOR2_X1 U308 ( .A(n191), .B(n190), .ZN(data_addr_o[19]) );
  NAND2_X1 U309 ( .A1(n338), .A2(n194), .ZN(n196) );
  INV_X1 U310 ( .A(n192), .ZN(n193) );
  AOI21_X1 U311 ( .B1(n344), .B2(n194), .A(n193), .ZN(n195) );
  OAI21_X1 U312 ( .B1(n263), .B2(n196), .A(n195), .ZN(n201) );
  INV_X1 U313 ( .A(n197), .ZN(n199) );
  NAND2_X1 U314 ( .A1(n199), .A2(n198), .ZN(n200) );
  XNOR2_X1 U315 ( .A(n201), .B(n200), .ZN(data_addr_o[25]) );
  INV_X1 U316 ( .A(n202), .ZN(n205) );
  INV_X1 U317 ( .A(n203), .ZN(n204) );
  OAI21_X1 U318 ( .B1(n263), .B2(n205), .A(n204), .ZN(n209) );
  NAND2_X1 U319 ( .A1(n207), .A2(n206), .ZN(n208) );
  XNOR2_X1 U320 ( .A(n209), .B(n208), .ZN(data_addr_o[18]) );
  INV_X1 U321 ( .A(n210), .ZN(n211) );
  NOR2_X1 U322 ( .A1(n211), .A2(n214), .ZN(n217) );
  NAND2_X1 U323 ( .A1(n217), .A2(n305), .ZN(n219) );
  INV_X1 U324 ( .A(n212), .ZN(n215) );
  OAI21_X1 U325 ( .B1(n215), .B2(n214), .A(n213), .ZN(n216) );
  AOI21_X1 U326 ( .B1(n217), .B2(n309), .A(n216), .ZN(n218) );
  OAI21_X1 U327 ( .B1(n263), .B2(n219), .A(n218), .ZN(n224) );
  INV_X1 U328 ( .A(n220), .ZN(n222) );
  NAND2_X1 U329 ( .A1(n222), .A2(n221), .ZN(n223) );
  XNOR2_X1 U330 ( .A(n224), .B(n223), .ZN(data_addr_o[23]) );
  INV_X1 U331 ( .A(n235), .ZN(n225) );
  NOR2_X1 U332 ( .A1(n225), .A2(n237), .ZN(n228) );
  INV_X1 U333 ( .A(n234), .ZN(n226) );
  OAI21_X1 U334 ( .B1(n226), .B2(n237), .A(n238), .ZN(n227) );
  AOI21_X1 U335 ( .B1(n228), .B2(n236), .A(n227), .ZN(n233) );
  INV_X1 U336 ( .A(n229), .ZN(n231) );
  NAND2_X1 U337 ( .A1(n231), .A2(n230), .ZN(n232) );
  XOR2_X1 U338 ( .A(n233), .B(n232), .Z(data_addr_o[7]) );
  AOI21_X1 U339 ( .B1(n236), .B2(n235), .A(n234), .ZN(n241) );
  INV_X1 U340 ( .A(n237), .ZN(n239) );
  NAND2_X1 U341 ( .A1(n239), .A2(n238), .ZN(n240) );
  XOR2_X1 U342 ( .A(n241), .B(n240), .Z(data_addr_o[6]) );
  NAND2_X1 U343 ( .A1(n242), .A2(n245), .ZN(n248) );
  INV_X1 U344 ( .A(n243), .ZN(n244) );
  AOI21_X1 U345 ( .B1(n246), .B2(n245), .A(n244), .ZN(n247) );
  OAI21_X1 U346 ( .B1(n299), .B2(n248), .A(n247), .ZN(n253) );
  INV_X1 U347 ( .A(n249), .ZN(n251) );
  NAND2_X1 U348 ( .A1(n251), .A2(n250), .ZN(n252) );
  XNOR2_X1 U349 ( .A(n253), .B(n252), .ZN(data_addr_o[11]) );
  OAI21_X1 U350 ( .B1(n299), .B2(n255), .A(n254), .ZN(n260) );
  INV_X1 U351 ( .A(n256), .ZN(n258) );
  NAND2_X1 U352 ( .A1(n258), .A2(n257), .ZN(n259) );
  XNOR2_X1 U353 ( .A(n260), .B(n259), .ZN(data_addr_o[9]) );
  OAI21_X1 U354 ( .B1(n263), .B2(n262), .A(n261), .ZN(n266) );
  INV_X1 U355 ( .A(n264), .ZN(n308) );
  NAND2_X1 U356 ( .A1(n308), .A2(n306), .ZN(n265) );
  XNOR2_X1 U357 ( .A(n266), .B(n265), .ZN(data_addr_o[20]) );
  OAI21_X1 U358 ( .B1(n299), .B2(n271), .A(n267), .ZN(n270) );
  INV_X1 U359 ( .A(n268), .ZN(n274) );
  NAND2_X1 U360 ( .A1(n274), .A2(n272), .ZN(n269) );
  XNOR2_X1 U361 ( .A(n270), .B(n269), .ZN(data_addr_o[12]) );
  INV_X1 U362 ( .A(n271), .ZN(n289) );
  NAND2_X1 U363 ( .A1(n289), .A2(n274), .ZN(n276) );
  INV_X1 U364 ( .A(n267), .ZN(n295) );
  INV_X1 U365 ( .A(n272), .ZN(n273) );
  AOI21_X1 U366 ( .B1(n295), .B2(n274), .A(n273), .ZN(n275) );
  OAI21_X1 U367 ( .B1(n299), .B2(n276), .A(n275), .ZN(n281) );
  INV_X1 U368 ( .A(n277), .ZN(n279) );
  NAND2_X1 U369 ( .A1(n279), .A2(n278), .ZN(n280) );
  NAND2_X1 U371 ( .A1(n289), .A2(n287), .ZN(n283) );
  AOI21_X1 U372 ( .B1(n295), .B2(n287), .A(n290), .ZN(n282) );
  OAI21_X1 U373 ( .B1(n299), .B2(n283), .A(n282), .ZN(n286) );
  INV_X1 U374 ( .A(n292), .ZN(n284) );
  NAND2_X1 U375 ( .A1(n284), .A2(n291), .ZN(n285) );
  XNOR2_X1 U376 ( .A(n286), .B(n285), .ZN(data_addr_o[14]) );
  INV_X1 U377 ( .A(n287), .ZN(n288) );
  NOR2_X1 U378 ( .A1(n288), .A2(n292), .ZN(n296) );
  NAND2_X1 U379 ( .A1(n296), .A2(n289), .ZN(n298) );
  INV_X1 U380 ( .A(n290), .ZN(n293) );
  OAI21_X1 U381 ( .B1(n293), .B2(n292), .A(n291), .ZN(n294) );
  AOI21_X1 U382 ( .B1(n296), .B2(n295), .A(n294), .ZN(n297) );
  OAI21_X1 U383 ( .B1(n299), .B2(n298), .A(n297), .ZN(n304) );
  INV_X1 U384 ( .A(n300), .ZN(n302) );
  NAND2_X1 U385 ( .A1(n302), .A2(n301), .ZN(n303) );
  XNOR2_X1 U386 ( .A(n304), .B(n303), .ZN(data_addr_o[15]) );
  NAND2_X1 U387 ( .A1(n305), .A2(n308), .ZN(n311) );
  INV_X1 U388 ( .A(n306), .ZN(n307) );
  AOI21_X1 U389 ( .B1(n309), .B2(n308), .A(n307), .ZN(n310) );
  OAI21_X1 U390 ( .B1(n263), .B2(n311), .A(n310), .ZN(n316) );
  INV_X1 U391 ( .A(n312), .ZN(n314) );
  NAND2_X1 U392 ( .A1(n314), .A2(n313), .ZN(n315) );
  XNOR2_X1 U393 ( .A(n316), .B(n315), .ZN(data_addr_o[21]) );
  NAND2_X1 U394 ( .A1(n338), .A2(n322), .ZN(n318) );
  AOI21_X1 U395 ( .B1(n344), .B2(n322), .A(n324), .ZN(n317) );
  OAI21_X1 U396 ( .B1(n263), .B2(n318), .A(n317), .ZN(n321) );
  INV_X1 U397 ( .A(n326), .ZN(n319) );
  NAND2_X1 U398 ( .A1(n319), .A2(n325), .ZN(n320) );
  INV_X1 U400 ( .A(n322), .ZN(n323) );
  NOR2_X1 U401 ( .A1(n323), .A2(n326), .ZN(n329) );
  NAND2_X1 U402 ( .A1(n338), .A2(n329), .ZN(n331) );
  INV_X1 U403 ( .A(n324), .ZN(n327) );
  OAI21_X1 U404 ( .B1(n327), .B2(n326), .A(n325), .ZN(n328) );
  AOI21_X1 U405 ( .B1(n344), .B2(n329), .A(n328), .ZN(n330) );
  OAI21_X1 U406 ( .B1(n263), .B2(n331), .A(n330), .ZN(n336) );
  INV_X1 U407 ( .A(n332), .ZN(n334) );
  NAND2_X1 U408 ( .A1(n334), .A2(n333), .ZN(n335) );
  XNOR2_X1 U409 ( .A(n336), .B(n335), .ZN(data_addr_o[27]) );
  NOR2_X1 U410 ( .A1(n337), .A2(n340), .ZN(n343) );
  NAND2_X1 U411 ( .A1(n338), .A2(n343), .ZN(n346) );
  OAI21_X1 U412 ( .B1(n341), .B2(n340), .A(n339), .ZN(n342) );
  AOI21_X1 U413 ( .B1(n344), .B2(n343), .A(n342), .ZN(n345) );
  OAI21_X1 U414 ( .B1(n263), .B2(n346), .A(n345), .ZN(n351) );
  INV_X1 U415 ( .A(n347), .ZN(n349) );
  NAND2_X1 U416 ( .A1(n349), .A2(n348), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n351), .B(n350), .ZN(data_addr_o[29]) );
  AND2_X1 U418 ( .A1(n730), .A2(rdata_offset_q[0]), .ZN(n374) );
  NAND2_X1 U419 ( .A1(n374), .A2(n509), .ZN(n508) );
  INV_X1 U420 ( .A(data_rdata_i[19]), .ZN(n608) );
  AND2_X1 U421 ( .A1(n731), .A2(rdata_offset_q[1]), .ZN(n448) );
  INV_X1 U422 ( .A(n509), .ZN(n352) );
  NAND2_X1 U423 ( .A1(n448), .A2(n352), .ZN(n452) );
  OAI22_X1 U424 ( .A1(n508), .A2(n744), .B1(n608), .B2(n452), .ZN(n356) );
  AND2_X1 U425 ( .A1(n448), .A2(n509), .ZN(n566) );
  INV_X1 U426 ( .A(n566), .ZN(n544) );
  NOR2_X2 U427 ( .A1(rdata_offset_q[1]), .A2(rdata_offset_q[0]), .ZN(n522) );
  INV_X1 U428 ( .A(n374), .ZN(n445) );
  NOR2_X1 U429 ( .A1(n509), .A2(n445), .ZN(n453) );
  AOI22_X1 U430 ( .A1(n522), .A2(data_rdata_i[3]), .B1(data_rdata_i[11]), .B2(
        n453), .ZN(n354) );
  AND2_X1 U431 ( .A1(rdata_offset_q[1]), .A2(rdata_offset_q[0]), .ZN(n523) );
  AND2_X1 U432 ( .A1(n523), .A2(data_type_q[1]), .ZN(n454) );
  INV_X1 U433 ( .A(n523), .ZN(n373) );
  NOR2_X1 U434 ( .A1(n373), .A2(data_type_q[1]), .ZN(n513) );
  AOI22_X1 U435 ( .A1(n454), .A2(data_rdata_i[27]), .B1(rdata_q[27]), .B2(n513), .ZN(n353) );
  OAI211_X1 U436 ( .C1(n544), .C2(n752), .A(n354), .B(n353), .ZN(n355) );
  NOR2_X1 U437 ( .A1(n356), .A2(n355), .ZN(n719) );
  MUX2_X1 U438 ( .A(n719), .B(n763), .S(n459), .Z(n357) );
  INV_X1 U439 ( .A(data_rdata_i[22]), .ZN(n623) );
  OAI22_X1 U440 ( .A1(n508), .A2(n747), .B1(n623), .B2(n452), .ZN(n361) );
  AOI22_X1 U441 ( .A1(n522), .A2(data_rdata_i[6]), .B1(data_rdata_i[14]), .B2(
        n453), .ZN(n359) );
  AOI22_X1 U442 ( .A1(n454), .A2(data_rdata_i[30]), .B1(rdata_q[30]), .B2(n513), .ZN(n358) );
  OAI211_X1 U443 ( .C1(n544), .C2(n755), .A(n359), .B(n358), .ZN(n360) );
  NOR2_X1 U444 ( .A1(n361), .A2(n360), .ZN(n713) );
  MUX2_X1 U445 ( .A(n713), .B(n766), .S(n459), .Z(n362) );
  INV_X1 U446 ( .A(data_rdata_i[16]), .ZN(n592) );
  OAI22_X1 U447 ( .A1(n592), .A2(n452), .B1(n508), .B2(n741), .ZN(n366) );
  AOI22_X1 U448 ( .A1(n522), .A2(data_rdata_i[0]), .B1(data_rdata_i[8]), .B2(
        n453), .ZN(n364) );
  AOI22_X1 U449 ( .A1(n454), .A2(data_rdata_i[24]), .B1(rdata_q[24]), .B2(n513), .ZN(n363) );
  OAI211_X1 U450 ( .C1(n544), .C2(n749), .A(n364), .B(n363), .ZN(n365) );
  NOR2_X1 U451 ( .A1(n366), .A2(n365), .ZN(n727) );
  MUX2_X1 U452 ( .A(n727), .B(n760), .S(n459), .Z(n367) );
  AND2_X1 U453 ( .A1(n522), .A2(n509), .ZN(n589) );
  NAND2_X1 U454 ( .A1(data_rvalid_i), .A2(n589), .ZN(n548) );
  INV_X1 U455 ( .A(data_rdata_i[28]), .ZN(n380) );
  INV_X1 U456 ( .A(n508), .ZN(n561) );
  INV_X1 U457 ( .A(data_rdata_i[12]), .ZN(n610) );
  NAND2_X1 U458 ( .A1(n509), .A2(n523), .ZN(n564) );
  INV_X1 U459 ( .A(data_rdata_i[20]), .ZN(n613) );
  OAI22_X1 U460 ( .A1(n544), .A2(n610), .B1(n564), .B2(n613), .ZN(n378) );
  NAND2_X1 U461 ( .A1(data_rdata_i[15]), .A2(n374), .ZN(n370) );
  NAND2_X1 U462 ( .A1(data_rdata_i[7]), .A2(n522), .ZN(n369) );
  NAND2_X1 U463 ( .A1(data_rdata_i[23]), .A2(n448), .ZN(n368) );
  AND3_X1 U464 ( .A1(n370), .A2(n369), .A3(n368), .ZN(n510) );
  NAND2_X1 U465 ( .A1(data_rdata_i[31]), .A2(n454), .ZN(n507) );
  OAI21_X1 U466 ( .B1(n510), .B2(n729), .A(n507), .ZN(n371) );
  NAND2_X1 U467 ( .A1(n371), .A2(data_sign_ext_q_0_), .ZN(n526) );
  NAND2_X1 U468 ( .A1(n526), .A2(data_type_q[1]), .ZN(n531) );
  INV_X1 U469 ( .A(data_rdata_i[7]), .ZN(n633) );
  AOI22_X1 U470 ( .A1(data_rdata_i[31]), .A2(n448), .B1(data_rdata_i[15]), 
        .B2(n522), .ZN(n372) );
  OAI21_X1 U471 ( .B1(n373), .B2(n633), .A(n372), .ZN(n376) );
  AND2_X1 U472 ( .A1(n374), .A2(data_type_q[0]), .ZN(n525) );
  AND2_X1 U473 ( .A1(data_rdata_i[23]), .A2(n525), .ZN(n375) );
  AOI21_X1 U474 ( .B1(n376), .B2(data_type_q[0]), .A(n375), .ZN(n518) );
  OAI21_X1 U475 ( .B1(n518), .B2(n759), .A(n526), .ZN(n377) );
  NAND2_X1 U476 ( .A1(n531), .A2(n377), .ZN(n562) );
  INV_X1 U477 ( .A(n562), .ZN(n545) );
  AOI211_X1 U478 ( .C1(data_rdata_i[4]), .C2(n561), .A(n378), .B(n545), .ZN(
        n612) );
  MUX2_X1 U479 ( .A(n737), .B(n612), .S(data_rvalid_i), .Z(n379) );
  OAI21_X1 U480 ( .B1(n548), .B2(n380), .A(n379), .ZN(data_rdata_ex_o[28]) );
  INV_X1 U481 ( .A(data_rdata_i[30]), .ZN(n383) );
  INV_X1 U482 ( .A(data_rdata_i[14]), .ZN(n620) );
  OAI22_X1 U483 ( .A1(n544), .A2(n620), .B1(n564), .B2(n623), .ZN(n381) );
  AOI211_X1 U484 ( .C1(data_rdata_i[6]), .C2(n561), .A(n381), .B(n545), .ZN(
        n622) );
  MUX2_X1 U485 ( .A(n739), .B(n622), .S(data_rvalid_i), .Z(n382) );
  OAI21_X1 U486 ( .B1(n548), .B2(n383), .A(n382), .ZN(data_rdata_ex_o[30]) );
  INV_X1 U487 ( .A(data_rdata_i[27]), .ZN(n386) );
  INV_X1 U488 ( .A(data_rdata_i[11]), .ZN(n605) );
  OAI22_X1 U489 ( .A1(n544), .A2(n605), .B1(n564), .B2(n608), .ZN(n384) );
  AOI211_X1 U490 ( .C1(data_rdata_i[3]), .C2(n561), .A(n384), .B(n545), .ZN(
        n607) );
  MUX2_X1 U491 ( .A(n736), .B(n607), .S(data_rvalid_i), .Z(n385) );
  OAI21_X1 U492 ( .B1(n548), .B2(n386), .A(n385), .ZN(data_rdata_ex_o[27]) );
  OAI22_X1 U493 ( .A1(n508), .A2(n745), .B1(n613), .B2(n452), .ZN(n423) );
  AOI22_X1 U494 ( .A1(n522), .A2(data_rdata_i[4]), .B1(data_rdata_i[12]), .B2(
        n453), .ZN(n388) );
  AOI22_X1 U495 ( .A1(n454), .A2(data_rdata_i[28]), .B1(rdata_q[28]), .B2(n513), .ZN(n387) );
  OAI211_X1 U496 ( .C1(n544), .C2(n753), .A(n388), .B(n387), .ZN(n389) );
  NOR2_X1 U497 ( .A1(n423), .A2(n389), .ZN(n717) );
  MUX2_X1 U498 ( .A(n717), .B(n764), .S(n459), .Z(n431) );
  INV_X1 U499 ( .A(data_rdata_i[21]), .ZN(n618) );
  OAI22_X1 U500 ( .A1(n508), .A2(n746), .B1(n618), .B2(n452), .ZN(n435) );
  AOI22_X1 U501 ( .A1(n522), .A2(data_rdata_i[5]), .B1(data_rdata_i[13]), .B2(
        n453), .ZN(n433) );
  AOI22_X1 U502 ( .A1(n454), .A2(data_rdata_i[29]), .B1(rdata_q[29]), .B2(n513), .ZN(n432) );
  OAI211_X1 U503 ( .C1(n544), .C2(n754), .A(n433), .B(n432), .ZN(n434) );
  NOR2_X1 U504 ( .A1(n435), .A2(n434), .ZN(n715) );
  MUX2_X1 U505 ( .A(n715), .B(n765), .S(n459), .Z(n436) );
  INV_X1 U506 ( .A(data_rdata_i[29]), .ZN(n439) );
  INV_X1 U507 ( .A(data_rdata_i[13]), .ZN(n615) );
  OAI22_X1 U508 ( .A1(n544), .A2(n615), .B1(n564), .B2(n618), .ZN(n437) );
  AOI211_X1 U509 ( .C1(data_rdata_i[5]), .C2(n561), .A(n437), .B(n545), .ZN(
        n617) );
  MUX2_X1 U510 ( .A(n738), .B(n617), .S(data_rvalid_i), .Z(n438) );
  OAI21_X1 U511 ( .B1(n548), .B2(n439), .A(n438), .ZN(data_rdata_ex_o[29]) );
  INV_X1 U512 ( .A(data_rdata_i[18]), .ZN(n603) );
  OAI22_X1 U513 ( .A1(n508), .A2(n743), .B1(n603), .B2(n452), .ZN(n443) );
  AOI22_X1 U514 ( .A1(n522), .A2(data_rdata_i[2]), .B1(data_rdata_i[10]), .B2(
        n453), .ZN(n441) );
  AOI22_X1 U515 ( .A1(n454), .A2(data_rdata_i[26]), .B1(rdata_q[26]), .B2(n513), .ZN(n440) );
  OAI211_X1 U516 ( .C1(n544), .C2(n751), .A(n441), .B(n440), .ZN(n442) );
  NOR2_X1 U517 ( .A1(n443), .A2(n442), .ZN(n721) );
  MUX2_X1 U518 ( .A(n721), .B(n762), .S(n459), .Z(n444) );
  AOI22_X1 U519 ( .A1(n523), .A2(data_rdata_i[3]), .B1(n522), .B2(
        data_rdata_i[11]), .ZN(n447) );
  NOR2_X1 U520 ( .A1(n445), .A2(data_type_q[0]), .ZN(n524) );
  AOI22_X1 U521 ( .A1(data_rdata_i[19]), .A2(n525), .B1(rdata_q[19]), .B2(n524), .ZN(n446) );
  NAND3_X1 U522 ( .A1(n447), .A2(n446), .A3(n526), .ZN(n450) );
  NAND2_X1 U523 ( .A1(n448), .A2(n756), .ZN(n530) );
  NAND2_X1 U524 ( .A1(n448), .A2(data_type_q[0]), .ZN(n529) );
  OAI22_X1 U525 ( .A1(n736), .A2(n530), .B1(n386), .B2(n529), .ZN(n449) );
  OAI21_X1 U526 ( .B1(n450), .B2(n449), .A(n531), .ZN(n606) );
  INV_X1 U527 ( .A(n606), .ZN(n451) );
  INV_X1 U528 ( .A(data_rdata_i[17]), .ZN(n598) );
  OAI22_X1 U529 ( .A1(n508), .A2(n742), .B1(n598), .B2(n452), .ZN(n458) );
  AOI22_X1 U530 ( .A1(n522), .A2(data_rdata_i[1]), .B1(data_rdata_i[9]), .B2(
        n453), .ZN(n456) );
  AOI22_X1 U531 ( .A1(n454), .A2(data_rdata_i[25]), .B1(rdata_q[25]), .B2(n513), .ZN(n455) );
  OAI211_X1 U532 ( .C1(n544), .C2(n750), .A(n456), .B(n455), .ZN(n457) );
  NOR2_X1 U533 ( .A1(n458), .A2(n457), .ZN(n723) );
  MUX2_X1 U534 ( .A(n723), .B(n761), .S(n459), .Z(n460) );
  AOI22_X1 U535 ( .A1(n523), .A2(data_rdata_i[1]), .B1(n522), .B2(
        data_rdata_i[9]), .ZN(n462) );
  AOI22_X1 U536 ( .A1(data_rdata_i[17]), .A2(n525), .B1(rdata_q[17]), .B2(n524), .ZN(n461) );
  NAND3_X1 U537 ( .A1(n462), .A2(n461), .A3(n526), .ZN(n464) );
  INV_X1 U538 ( .A(data_rdata_i[25]), .ZN(n596) );
  OAI22_X1 U539 ( .A1(n734), .A2(n530), .B1(n596), .B2(n529), .ZN(n463) );
  OAI21_X1 U540 ( .B1(n464), .B2(n463), .A(n531), .ZN(n595) );
  INV_X1 U541 ( .A(n595), .ZN(n465) );
  AOI22_X1 U542 ( .A1(n523), .A2(data_rdata_i[0]), .B1(n522), .B2(
        data_rdata_i[8]), .ZN(n467) );
  AOI22_X1 U543 ( .A1(data_rdata_i[16]), .A2(n525), .B1(rdata_q[16]), .B2(n524), .ZN(n466) );
  NAND3_X1 U544 ( .A1(n467), .A2(n466), .A3(n526), .ZN(n469) );
  INV_X1 U545 ( .A(data_rdata_i[24]), .ZN(n590) );
  OAI22_X1 U546 ( .A1(n733), .A2(n530), .B1(n590), .B2(n529), .ZN(n468) );
  OAI21_X1 U547 ( .B1(n469), .B2(n468), .A(n531), .ZN(n587) );
  INV_X1 U548 ( .A(n587), .ZN(n470) );
  AOI22_X1 U549 ( .A1(n589), .A2(data_rdata_i[20]), .B1(n561), .B2(rdata_q[28]), .ZN(n471) );
  OAI211_X1 U550 ( .C1(n564), .C2(n610), .A(n471), .B(n562), .ZN(n472) );
  AOI21_X1 U551 ( .B1(n566), .B2(data_rdata_i[4]), .A(n472), .ZN(n614) );
  INV_X1 U552 ( .A(n614), .ZN(n473) );
  INV_X1 U553 ( .A(n564), .ZN(n504) );
  AOI22_X1 U554 ( .A1(data_rdata_i[23]), .A2(n589), .B1(n561), .B2(rdata_q[31]), .ZN(n474) );
  OAI211_X1 U555 ( .C1(n633), .C2(n544), .A(n474), .B(n562), .ZN(n475) );
  AOI21_X1 U556 ( .B1(data_rdata_i[15]), .B2(n504), .A(n475), .ZN(n629) );
  INV_X1 U557 ( .A(n629), .ZN(n476) );
  AOI22_X1 U558 ( .A1(n523), .A2(data_rdata_i[4]), .B1(n522), .B2(
        data_rdata_i[12]), .ZN(n478) );
  AOI22_X1 U559 ( .A1(data_rdata_i[20]), .A2(n525), .B1(rdata_q[20]), .B2(n524), .ZN(n477) );
  NAND3_X1 U560 ( .A1(n478), .A2(n477), .A3(n526), .ZN(n480) );
  OAI22_X1 U561 ( .A1(n737), .A2(n530), .B1(n380), .B2(n529), .ZN(n479) );
  OAI21_X1 U562 ( .B1(n480), .B2(n479), .A(n531), .ZN(n611) );
  INV_X1 U563 ( .A(n611), .ZN(n481) );
  INV_X1 U564 ( .A(data_rdata_i[9]), .ZN(n594) );
  AOI22_X1 U565 ( .A1(n589), .A2(data_rdata_i[17]), .B1(n561), .B2(rdata_q[25]), .ZN(n482) );
  OAI211_X1 U566 ( .C1(n564), .C2(n594), .A(n482), .B(n562), .ZN(n483) );
  AOI21_X1 U567 ( .B1(data_rdata_i[1]), .B2(n566), .A(n483), .ZN(n599) );
  INV_X1 U568 ( .A(n599), .ZN(n484) );
  MUX2_X2 U569 ( .A(rdata_q[17]), .B(n484), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[17]) );
  AOI22_X1 U570 ( .A1(n523), .A2(data_rdata_i[5]), .B1(n522), .B2(
        data_rdata_i[13]), .ZN(n486) );
  AOI22_X1 U571 ( .A1(data_rdata_i[21]), .A2(n525), .B1(rdata_q[21]), .B2(n524), .ZN(n485) );
  NAND3_X1 U572 ( .A1(n486), .A2(n485), .A3(n526), .ZN(n488) );
  OAI22_X1 U573 ( .A1(n738), .A2(n530), .B1(n439), .B2(n529), .ZN(n487) );
  OAI21_X1 U574 ( .B1(n488), .B2(n487), .A(n531), .ZN(n616) );
  INV_X1 U575 ( .A(n616), .ZN(n489) );
  AOI22_X1 U576 ( .A1(n589), .A2(data_rdata_i[19]), .B1(n561), .B2(rdata_q[27]), .ZN(n490) );
  OAI211_X1 U577 ( .C1(n564), .C2(n605), .A(n490), .B(n562), .ZN(n491) );
  AOI21_X1 U578 ( .B1(n566), .B2(data_rdata_i[3]), .A(n491), .ZN(n609) );
  INV_X1 U579 ( .A(n609), .ZN(n492) );
  INV_X1 U580 ( .A(data_rdata_i[26]), .ZN(n495) );
  INV_X1 U581 ( .A(data_rdata_i[10]), .ZN(n600) );
  OAI22_X1 U582 ( .A1(n544), .A2(n600), .B1(n564), .B2(n603), .ZN(n493) );
  AOI211_X1 U583 ( .C1(data_rdata_i[2]), .C2(n561), .A(n493), .B(n545), .ZN(
        n602) );
  MUX2_X1 U584 ( .A(n735), .B(n602), .S(data_rvalid_i), .Z(n494) );
  OAI21_X1 U585 ( .B1(n548), .B2(n495), .A(n494), .ZN(data_rdata_ex_o[26]) );
  AOI22_X1 U586 ( .A1(n523), .A2(data_rdata_i[2]), .B1(n522), .B2(
        data_rdata_i[10]), .ZN(n497) );
  AOI22_X1 U587 ( .A1(data_rdata_i[18]), .A2(n525), .B1(rdata_q[18]), .B2(n524), .ZN(n496) );
  NAND3_X1 U588 ( .A1(n497), .A2(n496), .A3(n526), .ZN(n499) );
  OAI22_X1 U589 ( .A1(n735), .A2(n530), .B1(n495), .B2(n529), .ZN(n498) );
  OAI21_X1 U590 ( .B1(n499), .B2(n498), .A(n531), .ZN(n601) );
  INV_X1 U591 ( .A(n601), .ZN(n500) );
  INV_X1 U592 ( .A(data_rdata_i[8]), .ZN(n586) );
  OAI22_X1 U593 ( .A1(n544), .A2(n586), .B1(n564), .B2(n592), .ZN(n501) );
  AOI211_X1 U594 ( .C1(data_rdata_i[0]), .C2(n561), .A(n501), .B(n545), .ZN(
        n591) );
  MUX2_X1 U595 ( .A(n733), .B(n591), .S(data_rvalid_i), .Z(n502) );
  OAI21_X2 U596 ( .B1(n548), .B2(n590), .A(n502), .ZN(data_rdata_ex_o[24]) );
  INV_X1 U597 ( .A(data_rdata_i[31]), .ZN(n506) );
  INV_X1 U598 ( .A(data_rdata_i[15]), .ZN(n626) );
  OAI22_X1 U599 ( .A1(n626), .A2(n544), .B1(n633), .B2(n508), .ZN(n503) );
  AOI211_X1 U600 ( .C1(data_rdata_i[23]), .C2(n504), .A(n503), .B(n545), .ZN(
        n631) );
  MUX2_X1 U601 ( .A(n757), .B(n631), .S(data_rvalid_i), .Z(n505) );
  OAI21_X1 U602 ( .B1(n548), .B2(n506), .A(n505), .ZN(data_rdata_ex_o[31]) );
  OAI21_X1 U603 ( .B1(n508), .B2(n748), .A(n507), .ZN(n512) );
  OAI22_X1 U604 ( .A1(n510), .A2(n509), .B1(n740), .B2(n544), .ZN(n511) );
  AOI211_X1 U605 ( .C1(n513), .C2(rdata_q[31]), .A(n512), .B(n511), .ZN(n635)
         );
  MUX2_X1 U606 ( .A(n758), .B(n635), .S(data_rvalid_i), .Z(n514) );
  OAI21_X1 U607 ( .B1(n548), .B2(n633), .A(n514), .ZN(data_rdata_ex_o[7]) );
  INV_X1 U608 ( .A(n548), .ZN(n520) );
  AOI22_X1 U609 ( .A1(n566), .A2(rdata_q[31]), .B1(n561), .B2(rdata_q[23]), 
        .ZN(n515) );
  OAI21_X1 U610 ( .B1(n564), .B2(n633), .A(n515), .ZN(n516) );
  INV_X1 U611 ( .A(n516), .ZN(n517) );
  OAI211_X1 U612 ( .C1(n518), .C2(data_type_q[1]), .A(n517), .B(n526), .ZN(
        n625) );
  MUX2_X1 U613 ( .A(rdata_q[15]), .B(n625), .S(data_rvalid_i), .Z(n519) );
  AOI21_X1 U614 ( .B1(n520), .B2(data_rdata_i[15]), .A(n519), .ZN(n521) );
  INV_X2 U615 ( .A(n521), .ZN(data_rdata_ex_o[15]) );
  AOI22_X1 U616 ( .A1(n523), .A2(data_rdata_i[6]), .B1(n522), .B2(
        data_rdata_i[14]), .ZN(n528) );
  AOI22_X1 U617 ( .A1(data_rdata_i[22]), .A2(n525), .B1(rdata_q[22]), .B2(n524), .ZN(n527) );
  NAND3_X1 U618 ( .A1(n528), .A2(n527), .A3(n526), .ZN(n533) );
  OAI22_X1 U619 ( .A1(n739), .A2(n530), .B1(n383), .B2(n529), .ZN(n532) );
  OAI21_X1 U620 ( .B1(n533), .B2(n532), .A(n531), .ZN(n621) );
  INV_X1 U621 ( .A(n621), .ZN(n534) );
  AOI22_X1 U622 ( .A1(n589), .A2(data_rdata_i[22]), .B1(n561), .B2(rdata_q[30]), .ZN(n535) );
  OAI211_X1 U623 ( .C1(n564), .C2(n620), .A(n535), .B(n562), .ZN(n536) );
  AOI21_X1 U624 ( .B1(n566), .B2(data_rdata_i[6]), .A(n536), .ZN(n624) );
  INV_X1 U625 ( .A(n624), .ZN(n537) );
  AOI22_X1 U626 ( .A1(n589), .A2(data_rdata_i[18]), .B1(n561), .B2(rdata_q[26]), .ZN(n538) );
  OAI211_X1 U627 ( .C1(n564), .C2(n600), .A(n538), .B(n562), .ZN(n539) );
  AOI21_X1 U628 ( .B1(n566), .B2(data_rdata_i[2]), .A(n539), .ZN(n604) );
  INV_X1 U629 ( .A(n604), .ZN(n540) );
  MUX2_X2 U630 ( .A(rdata_q[18]), .B(n540), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[18]) );
  AOI22_X1 U631 ( .A1(n589), .A2(data_rdata_i[21]), .B1(n561), .B2(rdata_q[29]), .ZN(n541) );
  OAI211_X1 U632 ( .C1(n564), .C2(n615), .A(n541), .B(n562), .ZN(n542) );
  AOI21_X1 U633 ( .B1(n566), .B2(data_rdata_i[5]), .A(n542), .ZN(n619) );
  INV_X1 U634 ( .A(n619), .ZN(n543) );
  MUX2_X2 U635 ( .A(rdata_q[21]), .B(n543), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[21]) );
  OAI22_X1 U636 ( .A1(n544), .A2(n594), .B1(n564), .B2(n598), .ZN(n546) );
  AOI211_X1 U637 ( .C1(data_rdata_i[1]), .C2(n561), .A(n546), .B(n545), .ZN(
        n597) );
  MUX2_X1 U638 ( .A(n734), .B(n597), .S(data_rvalid_i), .Z(n547) );
  OAI21_X1 U639 ( .B1(n548), .B2(n596), .A(n547), .ZN(data_rdata_ex_o[25]) );
  NOR2_X1 U640 ( .A1(n732), .A2(CS[1]), .ZN(n549) );
  NAND2_X1 U641 ( .A1(n459), .A2(n549), .ZN(lsu_ready_wb_o) );
  NOR3_X1 U642 ( .A1(data_addr_o[1]), .A2(data_addr_o[0]), .A3(
        data_type_ex_i[0]), .ZN(n553) );
  INV_X1 U643 ( .A(data_type_ex_i[1]), .ZN(n550) );
  NAND2_X1 U644 ( .A1(n774), .A2(n550), .ZN(n552) );
  INV_X1 U645 ( .A(n552), .ZN(n555) );
  NOR2_X1 U646 ( .A1(data_addr_o[0]), .A2(n555), .ZN(n557) );
  INV_X1 U647 ( .A(n557), .ZN(n551) );
  OAI22_X1 U648 ( .A1(n553), .A2(n552), .B1(data_addr_o[1]), .B2(n551), .ZN(
        data_be_o[0]) );
  INV_X1 U649 ( .A(data_addr_o[1]), .ZN(n638) );
  AOI21_X1 U650 ( .B1(data_addr_o[0]), .B2(data_type_ex_i[1]), .A(n570), .ZN(
        n556) );
  INV_X1 U651 ( .A(n570), .ZN(n554) );
  OAI22_X1 U652 ( .A1(n638), .A2(n556), .B1(data_type_ex_i[0]), .B2(n554), 
        .ZN(data_be_o[3]) );
  NAND3_X1 U653 ( .A1(data_addr_o[1]), .A2(n569), .A3(n555), .ZN(n560) );
  OAI21_X1 U654 ( .B1(data_addr_o[1]), .B2(n556), .A(n560), .ZN(data_be_o[1])
         );
  NAND3_X1 U655 ( .A1(n638), .A2(n570), .A3(n568), .ZN(n559) );
  NAND2_X1 U656 ( .A1(data_addr_o[1]), .A2(n557), .ZN(n558) );
  OAI211_X1 U657 ( .C1(n560), .C2(n153), .A(n559), .B(n558), .ZN(data_be_o[2])
         );
  AOI22_X1 U658 ( .A1(data_rdata_i[16]), .A2(n589), .B1(n561), .B2(rdata_q[24]), .ZN(n563) );
  OAI211_X1 U659 ( .C1(n586), .C2(n564), .A(n563), .B(n562), .ZN(n565) );
  AOI21_X1 U660 ( .B1(n566), .B2(data_rdata_i[0]), .A(n565), .ZN(n593) );
  INV_X1 U661 ( .A(n593), .ZN(n567) );
  MUX2_X2 U662 ( .A(rdata_q[16]), .B(n567), .S(data_rvalid_i), .Z(
        data_rdata_ex_o[16]) );
  NAND2_X1 U663 ( .A1(data_addr_o[1]), .A2(n568), .ZN(n573) );
  AOI21_X1 U664 ( .B1(n584), .B2(data_req_ex_i), .A(CS[1]), .ZN(n574) );
  NOR3_X1 U665 ( .A1(n574), .A2(data_rvalid_i), .A3(CS[0]), .ZN(n575) );
  AOI21_X1 U666 ( .B1(n584), .B2(n576), .A(n575), .ZN(n579) );
  INV_X1 U667 ( .A(ex_valid_i), .ZN(n581) );
  OAI21_X1 U668 ( .B1(ex_valid_i), .B2(n728), .A(lsu_ready_wb_o), .ZN(n580) );
  NAND2_X1 U669 ( .A1(n580), .A2(CS[0]), .ZN(n578) );
  NAND3_X1 U670 ( .A1(n581), .A2(CS[1]), .A3(data_rvalid_i), .ZN(n577) );
  OAI211_X1 U671 ( .C1(n579), .C2(n581), .A(n578), .B(n577), .ZN(n430) );
  INV_X1 U672 ( .A(n580), .ZN(n583) );
  NAND3_X1 U673 ( .A1(n581), .A2(n584), .A3(data_req_o), .ZN(n582) );
  OAI21_X1 U674 ( .B1(n583), .B2(n728), .A(n582), .ZN(n429) );
  INV_X1 U707 ( .A(n625), .ZN(n627) );
  INV_X1 U709 ( .A(data_rdata_i[23]), .ZN(n628) );
  INV_X1 U713 ( .A(data_req_ex_i), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(busy_o) );
  NOR2_X1 U715 ( .A1(n638), .A2(data_addr_o[0]), .ZN(n678) );
  CLKBUF_X1 U716 ( .A(n678), .Z(n688) );
  NOR2_X1 U717 ( .A1(data_addr_o[0]), .A2(data_addr_o[1]), .ZN(n651) );
  CLKBUF_X1 U718 ( .A(n651), .Z(n706) );
  AOI22_X1 U719 ( .A1(n688), .A2(data_wdata_ex_i[8]), .B1(n706), .B2(
        data_wdata_ex_i[24]), .ZN(n640) );
  NOR2_X1 U720 ( .A1(n153), .A2(data_addr_o[1]), .ZN(n683) );
  CLKBUF_X1 U721 ( .A(n683), .Z(n708) );
  AND2_X1 U722 ( .A1(data_addr_o[0]), .A2(data_addr_o[1]), .ZN(n707) );
  CLKBUF_X1 U723 ( .A(n707), .Z(n703) );
  AOI22_X1 U724 ( .A1(n708), .A2(data_wdata_ex_i[16]), .B1(data_wdata_ex_i[0]), 
        .B2(n703), .ZN(n639) );
  NAND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(data_wdata_o[24]) );
  AOI22_X1 U726 ( .A1(n688), .A2(data_wdata_ex_i[0]), .B1(n706), .B2(
        data_wdata_ex_i[16]), .ZN(n642) );
  AOI22_X1 U727 ( .A1(n708), .A2(data_wdata_ex_i[8]), .B1(data_wdata_ex_i[24]), 
        .B2(n703), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n642), .A2(n641), .ZN(data_wdata_o[16]) );
  AOI22_X1 U729 ( .A1(n688), .A2(data_wdata_ex_i[24]), .B1(n651), .B2(
        data_wdata_ex_i[8]), .ZN(n644) );
  AOI22_X1 U730 ( .A1(n708), .A2(data_wdata_ex_i[0]), .B1(data_wdata_ex_i[16]), 
        .B2(n703), .ZN(n643) );
  NAND2_X1 U731 ( .A1(n644), .A2(n643), .ZN(data_wdata_o[8]) );
  AOI22_X1 U732 ( .A1(n688), .A2(data_wdata_ex_i[16]), .B1(n651), .B2(
        data_wdata_ex_i[0]), .ZN(n646) );
  AOI22_X1 U733 ( .A1(n708), .A2(data_wdata_ex_i[24]), .B1(data_wdata_ex_i[8]), 
        .B2(n703), .ZN(n645) );
  NAND2_X1 U734 ( .A1(n646), .A2(n645), .ZN(data_wdata_o[0]) );
  AOI22_X1 U735 ( .A1(n688), .A2(data_wdata_ex_i[9]), .B1(n651), .B2(
        data_wdata_ex_i[25]), .ZN(n648) );
  AOI22_X1 U736 ( .A1(n708), .A2(data_wdata_ex_i[17]), .B1(data_wdata_ex_i[1]), 
        .B2(n703), .ZN(n647) );
  NAND2_X1 U737 ( .A1(n648), .A2(n647), .ZN(data_wdata_o[25]) );
  AOI22_X1 U738 ( .A1(n688), .A2(data_wdata_ex_i[1]), .B1(n651), .B2(
        data_wdata_ex_i[17]), .ZN(n650) );
  AOI22_X1 U739 ( .A1(n708), .A2(data_wdata_ex_i[9]), .B1(data_wdata_ex_i[25]), 
        .B2(n703), .ZN(n649) );
  NAND2_X1 U740 ( .A1(n650), .A2(n649), .ZN(data_wdata_o[17]) );
  AOI22_X1 U741 ( .A1(n688), .A2(data_wdata_ex_i[25]), .B1(n651), .B2(
        data_wdata_ex_i[9]), .ZN(n653) );
  AOI22_X1 U742 ( .A1(n708), .A2(data_wdata_ex_i[1]), .B1(data_wdata_ex_i[17]), 
        .B2(n703), .ZN(n652) );
  NAND2_X1 U743 ( .A1(n653), .A2(n652), .ZN(data_wdata_o[9]) );
  AOI22_X1 U744 ( .A1(n688), .A2(data_wdata_ex_i[17]), .B1(n706), .B2(
        data_wdata_ex_i[1]), .ZN(n655) );
  AOI22_X1 U745 ( .A1(n708), .A2(data_wdata_ex_i[25]), .B1(data_wdata_ex_i[9]), 
        .B2(n703), .ZN(n654) );
  NAND2_X1 U746 ( .A1(n655), .A2(n654), .ZN(data_wdata_o[1]) );
  AOI22_X1 U747 ( .A1(n688), .A2(data_wdata_ex_i[10]), .B1(n651), .B2(
        data_wdata_ex_i[26]), .ZN(n657) );
  AOI22_X1 U748 ( .A1(n708), .A2(data_wdata_ex_i[18]), .B1(data_wdata_ex_i[2]), 
        .B2(n703), .ZN(n656) );
  NAND2_X1 U749 ( .A1(n657), .A2(n656), .ZN(data_wdata_o[26]) );
  AOI22_X1 U750 ( .A1(n688), .A2(data_wdata_ex_i[2]), .B1(n651), .B2(
        data_wdata_ex_i[18]), .ZN(n659) );
  AOI22_X1 U751 ( .A1(n708), .A2(data_wdata_ex_i[10]), .B1(data_wdata_ex_i[26]), .B2(n707), .ZN(n658) );
  NAND2_X1 U752 ( .A1(n659), .A2(n658), .ZN(data_wdata_o[18]) );
  AOI22_X1 U753 ( .A1(n688), .A2(data_wdata_ex_i[26]), .B1(n651), .B2(
        data_wdata_ex_i[10]), .ZN(n661) );
  AOI22_X1 U754 ( .A1(n683), .A2(data_wdata_ex_i[2]), .B1(data_wdata_ex_i[18]), 
        .B2(n707), .ZN(n660) );
  NAND2_X1 U755 ( .A1(n661), .A2(n660), .ZN(data_wdata_o[10]) );
  AOI22_X1 U756 ( .A1(n688), .A2(data_wdata_ex_i[18]), .B1(n651), .B2(
        data_wdata_ex_i[2]), .ZN(n663) );
  AOI22_X1 U757 ( .A1(n683), .A2(data_wdata_ex_i[26]), .B1(data_wdata_ex_i[10]), .B2(n707), .ZN(n662) );
  NAND2_X1 U758 ( .A1(n663), .A2(n662), .ZN(data_wdata_o[2]) );
  AOI22_X1 U759 ( .A1(n688), .A2(data_wdata_ex_i[11]), .B1(n651), .B2(
        data_wdata_ex_i[27]), .ZN(n665) );
  AOI22_X1 U760 ( .A1(n683), .A2(data_wdata_ex_i[19]), .B1(data_wdata_ex_i[3]), 
        .B2(n707), .ZN(n664) );
  NAND2_X1 U761 ( .A1(n665), .A2(n664), .ZN(data_wdata_o[27]) );
  AOI22_X1 U762 ( .A1(n688), .A2(data_wdata_ex_i[3]), .B1(n706), .B2(
        data_wdata_ex_i[19]), .ZN(n667) );
  AOI22_X1 U763 ( .A1(n683), .A2(data_wdata_ex_i[11]), .B1(data_wdata_ex_i[27]), .B2(n707), .ZN(n666) );
  NAND2_X1 U764 ( .A1(n667), .A2(n666), .ZN(data_wdata_o[19]) );
  AOI22_X1 U765 ( .A1(n688), .A2(data_wdata_ex_i[27]), .B1(n706), .B2(
        data_wdata_ex_i[11]), .ZN(n669) );
  AOI22_X1 U766 ( .A1(n683), .A2(data_wdata_ex_i[3]), .B1(data_wdata_ex_i[19]), 
        .B2(n707), .ZN(n668) );
  NAND2_X1 U767 ( .A1(n669), .A2(n668), .ZN(data_wdata_o[11]) );
  AOI22_X1 U768 ( .A1(n688), .A2(data_wdata_ex_i[19]), .B1(n706), .B2(
        data_wdata_ex_i[3]), .ZN(n671) );
  AOI22_X1 U769 ( .A1(n683), .A2(data_wdata_ex_i[27]), .B1(data_wdata_ex_i[11]), .B2(n707), .ZN(n670) );
  NAND2_X1 U770 ( .A1(n671), .A2(n670), .ZN(data_wdata_o[3]) );
  AOI22_X1 U771 ( .A1(n688), .A2(data_wdata_ex_i[12]), .B1(n706), .B2(
        data_wdata_ex_i[28]), .ZN(n673) );
  AOI22_X1 U772 ( .A1(n683), .A2(data_wdata_ex_i[20]), .B1(data_wdata_ex_i[4]), 
        .B2(n707), .ZN(n672) );
  NAND2_X1 U773 ( .A1(n673), .A2(n672), .ZN(data_wdata_o[28]) );
  AOI22_X1 U774 ( .A1(n688), .A2(data_wdata_ex_i[4]), .B1(n706), .B2(
        data_wdata_ex_i[20]), .ZN(n675) );
  AOI22_X1 U775 ( .A1(n683), .A2(data_wdata_ex_i[12]), .B1(data_wdata_ex_i[28]), .B2(n707), .ZN(n674) );
  NAND2_X1 U776 ( .A1(n675), .A2(n674), .ZN(data_wdata_o[20]) );
  AOI22_X1 U777 ( .A1(n688), .A2(data_wdata_ex_i[28]), .B1(n706), .B2(
        data_wdata_ex_i[12]), .ZN(n677) );
  AOI22_X1 U778 ( .A1(n708), .A2(data_wdata_ex_i[4]), .B1(data_wdata_ex_i[20]), 
        .B2(n707), .ZN(n676) );
  NAND2_X1 U779 ( .A1(n677), .A2(n676), .ZN(data_wdata_o[12]) );
  AOI22_X1 U780 ( .A1(n678), .A2(data_wdata_ex_i[20]), .B1(n706), .B2(
        data_wdata_ex_i[4]), .ZN(n680) );
  AOI22_X1 U781 ( .A1(n683), .A2(data_wdata_ex_i[28]), .B1(data_wdata_ex_i[12]), .B2(n707), .ZN(n679) );
  NAND2_X1 U782 ( .A1(n680), .A2(n679), .ZN(data_wdata_o[4]) );
  AOI22_X1 U783 ( .A1(n688), .A2(data_wdata_ex_i[13]), .B1(n706), .B2(
        data_wdata_ex_i[29]), .ZN(n682) );
  AOI22_X1 U784 ( .A1(n708), .A2(data_wdata_ex_i[21]), .B1(data_wdata_ex_i[5]), 
        .B2(n707), .ZN(n681) );
  NAND2_X1 U785 ( .A1(n682), .A2(n681), .ZN(data_wdata_o[29]) );
  AOI22_X1 U786 ( .A1(n688), .A2(data_wdata_ex_i[5]), .B1(n706), .B2(
        data_wdata_ex_i[21]), .ZN(n685) );
  AOI22_X1 U787 ( .A1(n683), .A2(data_wdata_ex_i[13]), .B1(data_wdata_ex_i[29]), .B2(n707), .ZN(n684) );
  NAND2_X1 U788 ( .A1(n685), .A2(n684), .ZN(data_wdata_o[21]) );
  AOI22_X1 U789 ( .A1(n688), .A2(data_wdata_ex_i[29]), .B1(n706), .B2(
        data_wdata_ex_i[13]), .ZN(n687) );
  AOI22_X1 U790 ( .A1(n708), .A2(data_wdata_ex_i[5]), .B1(data_wdata_ex_i[21]), 
        .B2(n707), .ZN(n686) );
  NAND2_X1 U791 ( .A1(n687), .A2(n686), .ZN(data_wdata_o[13]) );
  AOI22_X1 U792 ( .A1(n688), .A2(data_wdata_ex_i[21]), .B1(n706), .B2(
        data_wdata_ex_i[5]), .ZN(n690) );
  AOI22_X1 U793 ( .A1(n708), .A2(data_wdata_ex_i[29]), .B1(data_wdata_ex_i[13]), .B2(n707), .ZN(n689) );
  NAND2_X1 U794 ( .A1(n690), .A2(n689), .ZN(data_wdata_o[5]) );
  AOI22_X1 U795 ( .A1(n678), .A2(data_wdata_ex_i[14]), .B1(n706), .B2(
        data_wdata_ex_i[30]), .ZN(n692) );
  AOI22_X1 U796 ( .A1(n708), .A2(data_wdata_ex_i[22]), .B1(data_wdata_ex_i[6]), 
        .B2(n707), .ZN(n691) );
  NAND2_X1 U797 ( .A1(n692), .A2(n691), .ZN(data_wdata_o[30]) );
  AOI22_X1 U798 ( .A1(n678), .A2(data_wdata_ex_i[6]), .B1(n706), .B2(
        data_wdata_ex_i[22]), .ZN(n694) );
  AOI22_X1 U799 ( .A1(n708), .A2(data_wdata_ex_i[14]), .B1(data_wdata_ex_i[30]), .B2(n707), .ZN(n693) );
  NAND2_X1 U800 ( .A1(n694), .A2(n693), .ZN(data_wdata_o[22]) );
  AOI22_X1 U801 ( .A1(n678), .A2(data_wdata_ex_i[30]), .B1(n706), .B2(
        data_wdata_ex_i[14]), .ZN(n696) );
  AOI22_X1 U802 ( .A1(n708), .A2(data_wdata_ex_i[6]), .B1(data_wdata_ex_i[22]), 
        .B2(n707), .ZN(n695) );
  NAND2_X1 U803 ( .A1(n696), .A2(n695), .ZN(data_wdata_o[14]) );
  AOI22_X1 U804 ( .A1(n678), .A2(data_wdata_ex_i[22]), .B1(n706), .B2(
        data_wdata_ex_i[6]), .ZN(n698) );
  AOI22_X1 U805 ( .A1(n708), .A2(data_wdata_ex_i[30]), .B1(data_wdata_ex_i[14]), .B2(n707), .ZN(n697) );
  NAND2_X1 U806 ( .A1(n698), .A2(n697), .ZN(data_wdata_o[6]) );
  AOI22_X1 U807 ( .A1(n678), .A2(data_wdata_ex_i[15]), .B1(n706), .B2(
        data_wdata_ex_i[31]), .ZN(n700) );
  AOI22_X1 U808 ( .A1(n708), .A2(data_wdata_ex_i[23]), .B1(data_wdata_ex_i[7]), 
        .B2(n707), .ZN(n699) );
  NAND2_X1 U809 ( .A1(n700), .A2(n699), .ZN(data_wdata_o[31]) );
  AOI22_X1 U810 ( .A1(n678), .A2(data_wdata_ex_i[7]), .B1(n706), .B2(
        data_wdata_ex_i[23]), .ZN(n702) );
  AOI22_X1 U811 ( .A1(n708), .A2(data_wdata_ex_i[15]), .B1(data_wdata_ex_i[31]), .B2(n703), .ZN(n701) );
  NAND2_X1 U812 ( .A1(n702), .A2(n701), .ZN(data_wdata_o[23]) );
  AOI22_X1 U813 ( .A1(n678), .A2(data_wdata_ex_i[31]), .B1(n706), .B2(
        data_wdata_ex_i[15]), .ZN(n705) );
  AOI22_X1 U814 ( .A1(n708), .A2(data_wdata_ex_i[7]), .B1(data_wdata_ex_i[23]), 
        .B2(n703), .ZN(n704) );
  NAND2_X1 U815 ( .A1(n705), .A2(n704), .ZN(data_wdata_o[15]) );
  AOI22_X1 U816 ( .A1(n678), .A2(data_wdata_ex_i[23]), .B1(n706), .B2(
        data_wdata_ex_i[7]), .ZN(n710) );
  AOI22_X1 U817 ( .A1(n708), .A2(data_wdata_ex_i[31]), .B1(data_wdata_ex_i[15]), .B2(n707), .ZN(n709) );
  NAND2_X1 U818 ( .A1(n710), .A2(n709), .ZN(data_wdata_o[7]) );
  SDFFR_X1 data_we_q_reg ( .D(data_we_ex_i), .SI(1'b0), .SE(1'b0), .CK(n874), 
        .RN(rst_n), .QN(n767) );
  SDFFR_X1 data_type_q_reg_1_ ( .D(data_type_ex_i[1]), .SI(1'b0), .SE(1'b0), 
        .CK(n874), .RN(rst_n), .Q(data_type_q[1]), .QN(n729) );
  SDFFR_X1 data_type_q_reg_0_ ( .D(data_type_ex_i[0]), .SI(1'b0), .SE(1'b0), 
        .CK(n874), .RN(rst_n), .Q(data_type_q[0]), .QN(n756) );
  SDFFR_X1 rdata_offset_q_reg_1_ ( .D(data_addr_o[1]), .SI(1'b0), .SE(1'b0), 
        .CK(n874), .RN(rst_n), .Q(rdata_offset_q[1]), .QN(n730) );
  SDFFR_X1 rdata_offset_q_reg_0_ ( .D(data_addr_o[0]), .SI(1'b0), .SE(1'b0), 
        .CK(n874), .RN(rst_n), .Q(rdata_offset_q[0]), .QN(n731) );
  SDFFR_X1 data_sign_ext_q_reg_0_ ( .D(data_sign_ext_ex_i[0]), .SI(1'b0), .SE(
        1'b0), .CK(n874), .RN(rst_n), .Q(data_sign_ext_q_0_), .QN(n759) );
  SDFFR_X1 rdata_q_reg_31_ ( .D(n876), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[31]), .QN(n757) );
  SDFFR_X1 rdata_q_reg_30_ ( .D(n877), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[30]), .QN(n739) );
  SDFFR_X1 rdata_q_reg_29_ ( .D(n878), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[29]), .QN(n738) );
  SDFFR_X1 rdata_q_reg_28_ ( .D(n879), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[28]), .QN(n737) );
  SDFFR_X1 rdata_q_reg_27_ ( .D(n880), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[27]), .QN(n736) );
  SDFFR_X1 rdata_q_reg_26_ ( .D(n881), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[26]), .QN(n735) );
  SDFFR_X1 rdata_q_reg_25_ ( .D(n882), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[25]), .QN(n734) );
  SDFFR_X1 rdata_q_reg_24_ ( .D(n883), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[24]), .QN(n733) );
  SDFFR_X1 rdata_q_reg_23_ ( .D(n884), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[23]), .QN(n740) );
  SDFFR_X1 rdata_q_reg_22_ ( .D(n885), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[22]), .QN(n755) );
  SDFFR_X1 rdata_q_reg_21_ ( .D(n886), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[21]), .QN(n754) );
  SDFFR_X1 rdata_q_reg_20_ ( .D(n887), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[20]), .QN(n753) );
  SDFFR_X1 rdata_q_reg_19_ ( .D(n888), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[19]), .QN(n752) );
  SDFFR_X1 rdata_q_reg_18_ ( .D(n889), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[18]), .QN(n751) );
  SDFFR_X1 rdata_q_reg_17_ ( .D(n890), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[17]), .QN(n750) );
  SDFFR_X1 rdata_q_reg_16_ ( .D(n891), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[16]), .QN(n749) );
  SDFFR_X1 rdata_q_reg_15_ ( .D(n892), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[15]), .QN(n748) );
  SDFFR_X1 rdata_q_reg_14_ ( .D(n893), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[14]), .QN(n747) );
  SDFFR_X1 rdata_q_reg_13_ ( .D(n894), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[13]), .QN(n746) );
  SDFFR_X1 rdata_q_reg_12_ ( .D(n895), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[12]), .QN(n745) );
  SDFFR_X1 rdata_q_reg_11_ ( .D(n896), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[11]), .QN(n744) );
  SDFFR_X1 rdata_q_reg_10_ ( .D(n897), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[10]), .QN(n743) );
  SDFFR_X1 rdata_q_reg_9_ ( .D(n898), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[9]), .QN(n742) );
  SDFFR_X1 rdata_q_reg_8_ ( .D(n899), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .Q(rdata_q[8]), .QN(n741) );
  SDFFR_X1 rdata_q_reg_7_ ( .D(n900), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .QN(n758) );
  SDFFR_X1 rdata_q_reg_6_ ( .D(n901), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .QN(n766) );
  SDFFR_X1 rdata_q_reg_5_ ( .D(n902), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .QN(n765) );
  SDFFR_X1 rdata_q_reg_4_ ( .D(n903), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .QN(n764) );
  SDFFR_X1 rdata_q_reg_3_ ( .D(n904), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .QN(n763) );
  SDFFR_X1 rdata_q_reg_2_ ( .D(n905), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .QN(n762) );
  SDFFR_X1 rdata_q_reg_1_ ( .D(n906), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .QN(n761) );
  SDFFR_X1 rdata_q_reg_0_ ( .D(n907), .SI(1'b0), .SE(1'b0), .CK(n908), .RN(
        rst_n), .QN(n760) );
  SDFFR_X1 CS_reg_0_ ( .D(n430), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(rst_n), 
        .Q(CS[0]), .QN(n732) );
  SDFFR_X1 CS_reg_1_ ( .D(n429), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(rst_n), 
        .Q(CS[1]), .QN(n728) );
  SNPS_CLOCK_GATE_HIGH_riscv_load_store_unit_0 clk_gate_rdata_q_reg_0_ ( .CLK(
        clk), .EN(n630), .ENCLK(n908), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_load_store_unit_1 clk_gate_data_sign_ext_q_reg_0_ ( 
        .CLK(clk), .EN(n584), .ENCLK(n874), .TE(1'b0) );
  NOR2_X1 U77 ( .A1(n28), .A2(operand_a_ex_i[5]), .ZN(n48) );
  NOR2_X1 U133 ( .A1(n73), .A2(operand_a_ex_i[11]), .ZN(n249) );
  OAI21_X1 U240 ( .B1(n261), .B2(n121), .A(n120), .ZN(n344) );
  NOR2_X1 U199 ( .A1(n262), .A2(n121), .ZN(n338) );
  INV_X4 U6 ( .A(data_rvalid_i), .ZN(n459) );
  CLKBUF_X1 U3 ( .A(n773), .Z(n768) );
  CLKBUF_X1 U5 ( .A(n773), .Z(n769) );
  BUF_X2 U8 ( .A(n773), .Z(n770) );
  INV_X1 U9 ( .A(addr_useincr_ex_i), .ZN(n773) );
  XNOR2_X1 U10 ( .A(n321), .B(n320), .ZN(data_addr_o[26]) );
  XNOR2_X1 U31 ( .A(n281), .B(n280), .ZN(data_addr_o[13]) );
  INV_X1 U44 ( .A(n772), .ZN(n771) );
  NOR2_X1 U59 ( .A1(n20), .A2(operand_a_ex_i[3]), .ZN(n57) );
  NOR2_X1 U81 ( .A1(n29), .A2(operand_a_ex_i[6]), .ZN(n237) );
  NOR2_X1 U142 ( .A1(n38), .A2(operand_a_ex_i[9]), .ZN(n256) );
  NOR2_X1 U370 ( .A1(n268), .A2(n277), .ZN(n287) );
  AND3_X1 U399 ( .A1(data_rvalid_i), .A2(data_req_ex_i), .A3(n728), .ZN(n576)
         );
  AND2_X1 U675 ( .A1(data_rvalid_i), .A2(n767), .ZN(n630) );
  OR2_X1 U676 ( .A1(data_misaligned_o), .A2(n774), .ZN(n772) );
  INV_X1 U677 ( .A(data_misaligned_ex_i), .ZN(n774) );
  OAI22_X1 U866 ( .A1(n506), .A2(n855), .B1(n631), .B2(n772), .ZN(n876) );
  NOR2_X1 U867 ( .A1(n589), .A2(n772), .ZN(n855) );
  OAI22_X1 U868 ( .A1(n383), .A2(n856), .B1(n622), .B2(n859), .ZN(n877) );
  OAI22_X1 U869 ( .A1(n439), .A2(n856), .B1(n617), .B2(n772), .ZN(n878) );
  NOR2_X1 U870 ( .A1(n589), .A2(n772), .ZN(n856) );
  OAI22_X1 U871 ( .A1(n380), .A2(n857), .B1(n612), .B2(n772), .ZN(n879) );
  OAI22_X1 U872 ( .A1(n386), .A2(n857), .B1(n607), .B2(n772), .ZN(n880) );
  NOR2_X1 U873 ( .A1(n589), .A2(n772), .ZN(n857) );
  OAI22_X1 U874 ( .A1(n495), .A2(n858), .B1(n602), .B2(n859), .ZN(n881) );
  OAI22_X1 U875 ( .A1(n596), .A2(n858), .B1(n597), .B2(n772), .ZN(n882) );
  NOR2_X1 U876 ( .A1(n589), .A2(n772), .ZN(n858) );
  OAI22_X1 U877 ( .A1(n590), .A2(n860), .B1(n591), .B2(n859), .ZN(n883) );
  AOI22_X1 U878 ( .A1(n771), .A2(n629), .B1(n628), .B2(n772), .ZN(n884) );
  AOI22_X1 U879 ( .A1(n771), .A2(n624), .B1(n623), .B2(n859), .ZN(n885) );
  AOI22_X1 U880 ( .A1(n771), .A2(n619), .B1(n618), .B2(n859), .ZN(n886) );
  INV_X1 U881 ( .A(n771), .ZN(n859) );
  AOI22_X1 U882 ( .A1(n771), .A2(n614), .B1(n613), .B2(n859), .ZN(n887) );
  AOI22_X1 U883 ( .A1(n771), .A2(n609), .B1(n608), .B2(n772), .ZN(n888) );
  AOI22_X1 U884 ( .A1(n771), .A2(n604), .B1(n603), .B2(n772), .ZN(n889) );
  AOI22_X1 U885 ( .A1(n771), .A2(n599), .B1(n598), .B2(n772), .ZN(n890) );
  AOI22_X1 U886 ( .A1(n771), .A2(n593), .B1(n592), .B2(n859), .ZN(n891) );
  OAI22_X1 U887 ( .A1(n626), .A2(n860), .B1(n627), .B2(n772), .ZN(n892) );
  NOR2_X1 U888 ( .A1(n589), .A2(n772), .ZN(n860) );
  AOI22_X1 U889 ( .A1(n771), .A2(n621), .B1(n620), .B2(n859), .ZN(n893) );
  AOI22_X1 U890 ( .A1(n771), .A2(n616), .B1(n615), .B2(n772), .ZN(n894) );
  AOI22_X1 U891 ( .A1(n771), .A2(n611), .B1(n610), .B2(n859), .ZN(n895) );
  AOI22_X1 U892 ( .A1(n771), .A2(n606), .B1(n605), .B2(n859), .ZN(n896) );
  AOI22_X1 U893 ( .A1(n771), .A2(n601), .B1(n600), .B2(n772), .ZN(n897) );
  AOI22_X1 U894 ( .A1(n771), .A2(n595), .B1(n594), .B2(n859), .ZN(n898) );
  AOI22_X1 U895 ( .A1(n771), .A2(n587), .B1(n586), .B2(n772), .ZN(n899) );
  OAI21_X1 U896 ( .B1(n771), .B2(n633), .A(n861), .ZN(n900) );
  AOI22_X1 U897 ( .A1(n771), .A2(n862), .B1(n509), .B2(n863), .ZN(n861) );
  OAI22_X1 U898 ( .A1(n633), .A2(n864), .B1(n865), .B2(n772), .ZN(n863) );
  INV_X1 U899 ( .A(n522), .ZN(n864) );
  AOI21_X1 U900 ( .B1(n865), .B2(n510), .A(n509), .ZN(n862) );
  AOI211_X1 U901 ( .C1(rdata_q[31]), .C2(n513), .A(n512), .B(n866), .ZN(n865)
         );
  NOR2_X1 U902 ( .A1(n544), .A2(n740), .ZN(n866) );
  OAI21_X1 U903 ( .B1(n859), .B2(n713), .A(n867), .ZN(n901) );
  NAND2_X1 U904 ( .A1(n859), .A2(data_rdata_i[6]), .ZN(n867) );
  OAI21_X1 U905 ( .B1(n859), .B2(n715), .A(n868), .ZN(n902) );
  NAND2_X1 U906 ( .A1(n859), .A2(data_rdata_i[5]), .ZN(n868) );
  OAI21_X1 U907 ( .B1(n859), .B2(n717), .A(n869), .ZN(n903) );
  NAND2_X1 U908 ( .A1(n859), .A2(data_rdata_i[4]), .ZN(n869) );
  OAI21_X1 U909 ( .B1(n859), .B2(n719), .A(n870), .ZN(n904) );
  NAND2_X1 U910 ( .A1(n859), .A2(data_rdata_i[3]), .ZN(n870) );
  OAI21_X1 U911 ( .B1(n859), .B2(n721), .A(n871), .ZN(n905) );
  NAND2_X1 U912 ( .A1(n772), .A2(data_rdata_i[2]), .ZN(n871) );
  OAI21_X1 U913 ( .B1(n859), .B2(n723), .A(n872), .ZN(n906) );
  NAND2_X1 U914 ( .A1(n859), .A2(data_rdata_i[1]), .ZN(n872) );
  OAI21_X1 U915 ( .B1(n772), .B2(n727), .A(n873), .ZN(n907) );
  NAND2_X1 U916 ( .A1(n859), .A2(data_rdata_i[0]), .ZN(n873) );
endmodule



    module riscv_ex_stage_FPU0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_DIV0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5 ( 
        clk, rst_n, alu_operator_i, alu_operand_a_i, alu_operand_b_i, 
        alu_operand_c_i, bmask_a_i, bmask_b_i, imm_vec_ext_i, alu_vec_mode_i, 
        alu_is_clpx_i, alu_is_subrot_i, alu_clpx_shift_i, mult_operator_i, 
        mult_operand_a_i, mult_operand_b_i, mult_operand_c_i, mult_en_i, 
        mult_signed_mode_i, mult_imm_i, mult_dot_op_a_i, mult_dot_op_b_i, 
        mult_dot_op_c_i, mult_dot_signed_i, mult_is_clpx_i, mult_clpx_shift_i, 
        mult_clpx_img_i, mult_multicycle_o, fpu_prec_i, fpu_fflags_o, 
        fpu_fflags_we_o, apu_en_i, apu_op_i, apu_lat_i, apu_operands_i, 
        apu_waddr_i, apu_flags_i, apu_read_regs_i, apu_read_regs_valid_i, 
        apu_read_dep_o, apu_write_regs_i, apu_write_regs_valid_i, 
        apu_write_dep_o, apu_perf_type_o, apu_perf_cont_o, apu_perf_wb_o, 
        apu_busy_o, apu_ready_wb_o, apu_master_req_o, apu_master_ready_o, 
        apu_master_gnt_i, apu_master_operands_o, apu_master_op_o, 
        apu_master_valid_i, apu_master_result_i, lsu_en_i, lsu_rdata_i, 
        branch_in_ex_i, regfile_alu_waddr_i, regfile_we_i, regfile_waddr_i, 
        csr_rdata_i, regfile_waddr_wb_o, regfile_we_wb_o, regfile_wdata_wb_o, 
        regfile_alu_waddr_fw_o, regfile_alu_we_fw_o, regfile_alu_wdata_fw_o, 
        jump_target_o, branch_decision_o, lsu_ready_ex_i, ex_ready_o, 
        ex_valid_o, wb_ready_i, lsu_err_i_BAR, regfile_alu_we_i, alu_en_i_BAR, 
        mult_sel_subword_i_BAR, csr_access_i_BAR );
  input [6:0] alu_operator_i;
  input [31:0] alu_operand_a_i;
  input [31:0] alu_operand_b_i;
  input [31:0] alu_operand_c_i;
  input [4:0] bmask_a_i;
  input [4:0] bmask_b_i;
  input [1:0] imm_vec_ext_i;
  input [1:0] alu_vec_mode_i;
  input [1:0] alu_clpx_shift_i;
  input [2:0] mult_operator_i;
  input [31:0] mult_operand_a_i;
  input [31:0] mult_operand_b_i;
  input [31:0] mult_operand_c_i;
  input [1:0] mult_signed_mode_i;
  input [4:0] mult_imm_i;
  input [31:0] mult_dot_op_a_i;
  input [31:0] mult_dot_op_b_i;
  input [31:0] mult_dot_op_c_i;
  input [1:0] mult_dot_signed_i;
  input [1:0] mult_clpx_shift_i;
  input [4:0] fpu_prec_i;
  output [4:0] fpu_fflags_o;
  input [5:0] apu_op_i;
  input [1:0] apu_lat_i;
  input [95:0] apu_operands_i;
  input [5:0] apu_waddr_i;
  input [14:0] apu_flags_i;
  input [17:0] apu_read_regs_i;
  input [2:0] apu_read_regs_valid_i;
  input [11:0] apu_write_regs_i;
  input [1:0] apu_write_regs_valid_i;
  output [95:0] apu_master_operands_o;
  output [5:0] apu_master_op_o;
  input [31:0] apu_master_result_i;
  input [31:0] lsu_rdata_i;
  input [5:0] regfile_alu_waddr_i;
  input [5:0] regfile_waddr_i;
  input [31:0] csr_rdata_i;
  output [5:0] regfile_waddr_wb_o;
  output [31:0] regfile_wdata_wb_o;
  output [5:0] regfile_alu_waddr_fw_o;
  output [31:0] regfile_alu_wdata_fw_o;
  output [31:0] jump_target_o;
  input clk, rst_n, alu_is_clpx_i, alu_is_subrot_i, mult_en_i, mult_is_clpx_i,
         mult_clpx_img_i, apu_en_i, apu_master_gnt_i, apu_master_valid_i,
         lsu_en_i, branch_in_ex_i, regfile_we_i, lsu_ready_ex_i, wb_ready_i,
         lsu_err_i_BAR, regfile_alu_we_i, alu_en_i_BAR, mult_sel_subword_i_BAR,
         csr_access_i_BAR;
  output mult_multicycle_o, fpu_fflags_we_o, apu_read_dep_o, apu_write_dep_o,
         apu_perf_type_o, apu_perf_cont_o, apu_perf_wb_o, apu_busy_o,
         apu_ready_wb_o, apu_master_req_o, apu_master_ready_o, regfile_we_wb_o,
         regfile_alu_we_fw_o, branch_decision_o, ex_ready_o, ex_valid_o;
  wire   regfile_alu_we_i, csr_access_i, alu_ready, mult_ready, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n167, n168, n169, n170, n171, n172, n173,
         n184, n185, n186, n199, n201;
  wire   [31:0] alu_result;
  wire   [31:0] mult_result;
  assign regfile_wdata_wb_o[31] = lsu_rdata_i[31];
  assign regfile_wdata_wb_o[30] = lsu_rdata_i[30];
  assign regfile_wdata_wb_o[29] = lsu_rdata_i[29];
  assign regfile_wdata_wb_o[28] = lsu_rdata_i[28];
  assign regfile_wdata_wb_o[27] = lsu_rdata_i[27];
  assign regfile_wdata_wb_o[26] = lsu_rdata_i[26];
  assign regfile_wdata_wb_o[25] = lsu_rdata_i[25];
  assign regfile_wdata_wb_o[24] = lsu_rdata_i[24];
  assign regfile_wdata_wb_o[23] = lsu_rdata_i[23];
  assign regfile_wdata_wb_o[22] = lsu_rdata_i[22];
  assign regfile_wdata_wb_o[21] = lsu_rdata_i[21];
  assign regfile_wdata_wb_o[20] = lsu_rdata_i[20];
  assign regfile_wdata_wb_o[19] = lsu_rdata_i[19];
  assign regfile_wdata_wb_o[18] = lsu_rdata_i[18];
  assign regfile_wdata_wb_o[17] = lsu_rdata_i[17];
  assign regfile_wdata_wb_o[16] = lsu_rdata_i[16];
  assign regfile_wdata_wb_o[15] = lsu_rdata_i[15];
  assign regfile_wdata_wb_o[14] = lsu_rdata_i[14];
  assign regfile_wdata_wb_o[13] = lsu_rdata_i[13];
  assign regfile_wdata_wb_o[12] = lsu_rdata_i[12];
  assign regfile_wdata_wb_o[11] = lsu_rdata_i[11];
  assign regfile_wdata_wb_o[10] = lsu_rdata_i[10];
  assign regfile_wdata_wb_o[9] = lsu_rdata_i[9];
  assign regfile_wdata_wb_o[8] = lsu_rdata_i[8];
  assign regfile_wdata_wb_o[7] = lsu_rdata_i[7];
  assign regfile_wdata_wb_o[6] = lsu_rdata_i[6];
  assign regfile_wdata_wb_o[5] = lsu_rdata_i[5];
  assign regfile_wdata_wb_o[4] = lsu_rdata_i[4];
  assign regfile_wdata_wb_o[3] = lsu_rdata_i[3];
  assign regfile_wdata_wb_o[2] = lsu_rdata_i[2];
  assign regfile_wdata_wb_o[1] = lsu_rdata_i[1];
  assign regfile_wdata_wb_o[0] = lsu_rdata_i[0];
  assign regfile_alu_waddr_fw_o[4] = regfile_alu_waddr_i[4];
  assign regfile_alu_waddr_fw_o[3] = regfile_alu_waddr_i[3];
  assign regfile_alu_waddr_fw_o[2] = regfile_alu_waddr_i[2];
  assign regfile_alu_waddr_fw_o[1] = regfile_alu_waddr_i[1];
  assign regfile_alu_waddr_fw_o[0] = regfile_alu_waddr_i[0];
  assign regfile_alu_we_fw_o = regfile_alu_we_i;
  assign csr_access_i = csr_access_i_BAR;
  assign jump_target_o[31] = alu_operand_c_i[31];
  assign jump_target_o[30] = alu_operand_c_i[30];
  assign jump_target_o[29] = alu_operand_c_i[29];
  assign jump_target_o[28] = alu_operand_c_i[28];
  assign jump_target_o[27] = alu_operand_c_i[27];
  assign jump_target_o[26] = alu_operand_c_i[26];
  assign jump_target_o[25] = alu_operand_c_i[25];
  assign jump_target_o[24] = alu_operand_c_i[24];
  assign jump_target_o[23] = alu_operand_c_i[23];
  assign jump_target_o[22] = alu_operand_c_i[22];
  assign jump_target_o[21] = alu_operand_c_i[21];
  assign jump_target_o[20] = alu_operand_c_i[20];
  assign jump_target_o[19] = alu_operand_c_i[19];
  assign jump_target_o[18] = alu_operand_c_i[18];
  assign jump_target_o[17] = alu_operand_c_i[17];
  assign jump_target_o[16] = alu_operand_c_i[16];
  assign jump_target_o[15] = alu_operand_c_i[15];
  assign jump_target_o[14] = alu_operand_c_i[14];
  assign jump_target_o[13] = alu_operand_c_i[13];
  assign jump_target_o[12] = alu_operand_c_i[12];
  assign jump_target_o[11] = alu_operand_c_i[11];
  assign jump_target_o[10] = alu_operand_c_i[10];
  assign jump_target_o[9] = alu_operand_c_i[9];
  assign jump_target_o[8] = alu_operand_c_i[8];
  assign jump_target_o[7] = alu_operand_c_i[7];
  assign jump_target_o[6] = alu_operand_c_i[6];
  assign jump_target_o[5] = alu_operand_c_i[5];
  assign jump_target_o[4] = alu_operand_c_i[4];
  assign jump_target_o[3] = alu_operand_c_i[3];
  assign jump_target_o[2] = alu_operand_c_i[2];
  assign jump_target_o[1] = alu_operand_c_i[1];

  INV_X1 U89 ( .A(rst_n) );
  NAND2_X2 U7 ( .A1(n133), .A2(n132), .ZN(regfile_alu_wdata_fw_o[17]) );
  NAND2_X2 U15 ( .A1(n123), .A2(n122), .ZN(regfile_alu_wdata_fw_o[13]) );
  AND2_X1 U25 ( .A1(csr_rdata_i[7]), .A2(n186), .ZN(n101) );
  AOI21_X1 U27 ( .B1(mult_result[7]), .B2(n163), .A(n101), .ZN(n91) );
  NAND2_X1 U28 ( .A1(n92), .A2(n153), .ZN(regfile_alu_wdata_fw_o[3]) );
  NAND2_X1 U29 ( .A1(alu_result[3]), .A2(n184), .ZN(n92) );
  INV_X1 U30 ( .A(alu_en_i_BAR), .ZN(n93) );
  CLKBUF_X1 U33 ( .A(ex_ready_o), .Z(n172) );
  AOI22_X1 U34 ( .A1(mult_result[15]), .A2(n167), .B1(csr_rdata_i[15]), .B2(
        n185), .ZN(n94) );
  INV_X1 U35 ( .A(mult_en_i), .ZN(n98) );
  NOR2_X1 U37 ( .A1(n98), .A2(n186), .ZN(n167) );
  AOI21_X1 U38 ( .B1(mult_result[5]), .B2(n163), .A(n115), .ZN(n116) );
  AND3_X1 U40 ( .A1(wb_ready_i), .A2(alu_ready), .A3(mult_ready), .ZN(n95) );
  NAND2_X1 U41 ( .A1(lsu_ready_ex_i), .A2(n95), .ZN(n114) );
  NOR4_X1 U42 ( .A1(n93), .A2(mult_en_i), .A3(n185), .A4(lsu_en_i), .ZN(n96)
         );
  NOR2_X1 U43 ( .A1(n114), .A2(n96), .ZN(ex_valid_o) );
  NAND3_X1 U44 ( .A1(ex_valid_o), .A2(regfile_we_i), .A3(lsu_err_i_BAR), .ZN(
        n170) );
  OAI21_X1 U45 ( .B1(wb_ready_i), .B2(n173), .A(n170), .ZN(n97) );
  INV_X1 U46 ( .A(n97), .ZN(n171) );
  AOI22_X1 U47 ( .A1(mult_result[0]), .A2(n163), .B1(n185), .B2(csr_rdata_i[0]), .ZN(n100) );
  NAND2_X1 U48 ( .A1(alu_result[0]), .A2(n184), .ZN(n99) );
  NAND2_X1 U49 ( .A1(alu_result[7]), .A2(n184), .ZN(n102) );
  NAND2_X1 U50 ( .A1(alu_result[29]), .A2(n184), .ZN(n105) );
  AOI22_X1 U51 ( .A1(mult_result[29]), .A2(n167), .B1(n185), .B2(
        csr_rdata_i[29]), .ZN(n104) );
  NAND2_X1 U52 ( .A1(alu_result[23]), .A2(n184), .ZN(n107) );
  AOI22_X1 U53 ( .A1(mult_result[23]), .A2(n163), .B1(n185), .B2(
        csr_rdata_i[23]), .ZN(n106) );
  NAND2_X1 U54 ( .A1(alu_result[9]), .A2(n184), .ZN(n109) );
  AOI22_X1 U55 ( .A1(mult_result[9]), .A2(n163), .B1(n185), .B2(csr_rdata_i[9]), .ZN(n108) );
  NAND2_X1 U57 ( .A1(alu_result[6]), .A2(n184), .ZN(n112) );
  NAND2_X1 U58 ( .A1(mult_result[6]), .A2(n163), .ZN(n111) );
  NAND2_X1 U59 ( .A1(csr_rdata_i[6]), .A2(n186), .ZN(n110) );
  INV_X1 U60 ( .A(branch_in_ex_i), .ZN(n113) );
  NAND2_X1 U61 ( .A1(n114), .A2(n113), .ZN(ex_ready_o) );
  NAND2_X1 U62 ( .A1(alu_result[5]), .A2(n184), .ZN(n117) );
  AND2_X1 U63 ( .A1(csr_rdata_i[5]), .A2(n186), .ZN(n115) );
  NAND2_X1 U64 ( .A1(n117), .A2(n116), .ZN(regfile_alu_wdata_fw_o[5]) );
  NAND2_X1 U65 ( .A1(alu_result[18]), .A2(n184), .ZN(n119) );
  AOI22_X1 U66 ( .A1(mult_result[18]), .A2(n163), .B1(n186), .B2(
        csr_rdata_i[18]), .ZN(n118) );
  NAND2_X1 U67 ( .A1(alu_result[14]), .A2(n184), .ZN(n121) );
  AOI22_X1 U68 ( .A1(mult_result[14]), .A2(n167), .B1(n185), .B2(
        csr_rdata_i[14]), .ZN(n120) );
  NAND2_X1 U69 ( .A1(alu_result[13]), .A2(n184), .ZN(n123) );
  AOI22_X1 U70 ( .A1(mult_result[13]), .A2(n167), .B1(n185), .B2(
        csr_rdata_i[13]), .ZN(n122) );
  NAND2_X1 U71 ( .A1(alu_result[28]), .A2(n184), .ZN(n125) );
  AOI22_X1 U72 ( .A1(mult_result[28]), .A2(n163), .B1(n185), .B2(
        csr_rdata_i[28]), .ZN(n124) );
  NAND2_X1 U73 ( .A1(alu_result[30]), .A2(n184), .ZN(n127) );
  AOI22_X1 U74 ( .A1(mult_result[30]), .A2(n167), .B1(n185), .B2(
        csr_rdata_i[30]), .ZN(n126) );
  NAND2_X1 U75 ( .A1(alu_result[27]), .A2(n184), .ZN(n129) );
  AOI22_X1 U76 ( .A1(mult_result[27]), .A2(n167), .B1(n186), .B2(
        csr_rdata_i[27]), .ZN(n128) );
  NAND2_X1 U77 ( .A1(alu_result[20]), .A2(n184), .ZN(n131) );
  AOI22_X1 U78 ( .A1(mult_result[20]), .A2(n163), .B1(n186), .B2(
        csr_rdata_i[20]), .ZN(n130) );
  NAND2_X1 U79 ( .A1(alu_result[17]), .A2(n184), .ZN(n133) );
  AOI22_X1 U80 ( .A1(mult_result[17]), .A2(n163), .B1(n185), .B2(
        csr_rdata_i[17]), .ZN(n132) );
  NAND2_X1 U81 ( .A1(alu_result[19]), .A2(n184), .ZN(n135) );
  AOI22_X1 U82 ( .A1(mult_result[19]), .A2(n163), .B1(n186), .B2(
        csr_rdata_i[19]), .ZN(n134) );
  NAND2_X1 U83 ( .A1(alu_result[26]), .A2(n184), .ZN(n137) );
  AOI22_X1 U84 ( .A1(mult_result[26]), .A2(n163), .B1(n186), .B2(
        csr_rdata_i[26]), .ZN(n136) );
  NAND2_X1 U85 ( .A1(n137), .A2(n136), .ZN(regfile_alu_wdata_fw_o[26]) );
  NAND2_X1 U86 ( .A1(alu_result[10]), .A2(n184), .ZN(n139) );
  AOI22_X1 U87 ( .A1(mult_result[10]), .A2(n163), .B1(n185), .B2(
        csr_rdata_i[10]), .ZN(n138) );
  NAND2_X1 U88 ( .A1(alu_result[31]), .A2(n184), .ZN(n141) );
  AOI22_X1 U90 ( .A1(mult_result[31]), .A2(n167), .B1(n186), .B2(
        csr_rdata_i[31]), .ZN(n140) );
  NAND2_X1 U91 ( .A1(alu_result[15]), .A2(n184), .ZN(n142) );
  NAND2_X1 U92 ( .A1(alu_result[22]), .A2(n184), .ZN(n144) );
  AOI22_X1 U93 ( .A1(mult_result[22]), .A2(n163), .B1(n185), .B2(
        csr_rdata_i[22]), .ZN(n143) );
  NAND2_X1 U94 ( .A1(alu_result[25]), .A2(n184), .ZN(n146) );
  NAND2_X1 U96 ( .A1(alu_result[2]), .A2(n184), .ZN(n148) );
  AOI22_X1 U97 ( .A1(mult_result[2]), .A2(n163), .B1(n186), .B2(csr_rdata_i[2]), .ZN(n147) );
  NAND2_X1 U98 ( .A1(n148), .A2(n147), .ZN(regfile_alu_wdata_fw_o[2]) );
  NAND2_X1 U99 ( .A1(alu_result[4]), .A2(n184), .ZN(n150) );
  AOI22_X1 U100 ( .A1(mult_result[4]), .A2(n163), .B1(n185), .B2(
        csr_rdata_i[4]), .ZN(n149) );
  NAND2_X1 U101 ( .A1(n150), .A2(n149), .ZN(regfile_alu_wdata_fw_o[4]) );
  NAND2_X1 U102 ( .A1(alu_result[1]), .A2(n184), .ZN(n152) );
  AOI22_X1 U103 ( .A1(mult_result[1]), .A2(n163), .B1(n185), .B2(
        csr_rdata_i[1]), .ZN(n151) );
  NAND2_X1 U104 ( .A1(n152), .A2(n151), .ZN(regfile_alu_wdata_fw_o[1]) );
  AOI22_X1 U105 ( .A1(mult_result[3]), .A2(n163), .B1(n185), .B2(
        csr_rdata_i[3]), .ZN(n153) );
  NAND2_X1 U106 ( .A1(alu_result[8]), .A2(n184), .ZN(n155) );
  AOI22_X1 U107 ( .A1(mult_result[8]), .A2(n163), .B1(n185), .B2(
        csr_rdata_i[8]), .ZN(n154) );
  NAND2_X1 U108 ( .A1(alu_result[11]), .A2(n184), .ZN(n158) );
  AOI22_X1 U109 ( .A1(mult_result[11]), .A2(n163), .B1(n185), .B2(
        csr_rdata_i[11]), .ZN(n157) );
  NAND2_X1 U110 ( .A1(n158), .A2(n157), .ZN(regfile_alu_wdata_fw_o[11]) );
  NAND2_X1 U111 ( .A1(alu_result[12]), .A2(n184), .ZN(n160) );
  AOI22_X1 U112 ( .A1(mult_result[12]), .A2(n167), .B1(n185), .B2(
        csr_rdata_i[12]), .ZN(n159) );
  NAND2_X1 U113 ( .A1(alu_result[16]), .A2(n184), .ZN(n162) );
  AOI22_X1 U114 ( .A1(mult_result[16]), .A2(n163), .B1(n185), .B2(
        csr_rdata_i[16]), .ZN(n161) );
  NAND2_X1 U115 ( .A1(n162), .A2(n161), .ZN(regfile_alu_wdata_fw_o[16]) );
  NAND2_X1 U116 ( .A1(alu_result[21]), .A2(n184), .ZN(n165) );
  AOI22_X1 U117 ( .A1(mult_result[21]), .A2(n163), .B1(n185), .B2(
        csr_rdata_i[21]), .ZN(n164) );
  NAND2_X1 U118 ( .A1(alu_result[24]), .A2(n184), .ZN(n169) );
  AOI22_X1 U119 ( .A1(mult_result[24]), .A2(n167), .B1(n185), .B2(
        csr_rdata_i[24]), .ZN(n168) );
  SDFFR_X1 regfile_waddr_lsu_reg_4_ ( .D(regfile_waddr_i[4]), .SI(1'b0), .SE(
        1'b0), .CK(n199), .RN(rst_n), .Q(regfile_waddr_wb_o[4]) );
  SDFFR_X1 regfile_waddr_lsu_reg_3_ ( .D(regfile_waddr_i[3]), .SI(1'b0), .SE(
        1'b0), .CK(n199), .RN(rst_n), .Q(regfile_waddr_wb_o[3]) );
  SDFFR_X1 regfile_waddr_lsu_reg_2_ ( .D(regfile_waddr_i[2]), .SI(1'b0), .SE(
        1'b0), .CK(n199), .RN(rst_n), .Q(regfile_waddr_wb_o[2]) );
  SDFFR_X1 regfile_waddr_lsu_reg_1_ ( .D(regfile_waddr_i[1]), .SI(1'b0), .SE(
        1'b0), .CK(n199), .RN(rst_n), .Q(regfile_waddr_wb_o[1]) );
  SDFFR_X1 regfile_waddr_lsu_reg_0_ ( .D(regfile_waddr_i[0]), .SI(1'b0), .SE(
        1'b0), .CK(n199), .RN(rst_n), .Q(regfile_waddr_wb_o[0]) );
  SDFFS_X1 regfile_we_lsu_reg ( .D(n171), .SI(1'b0), .SE(1'b0), .CK(clk), .SN(
        rst_n), .Q(n173), .QN(regfile_we_wb_o) );
  riscv_alu_SHARED_INT_DIV0_FPU0 alu_i ( .clk(clk), .rst_n(rst_n), 
        .operator_i(alu_operator_i), .operand_a_i(alu_operand_a_i), 
        .operand_b_i(alu_operand_b_i), .operand_c_i(alu_operand_c_i), 
        .vector_mode_i(alu_vec_mode_i), .bmask_a_i(bmask_a_i), .bmask_b_i(
        bmask_b_i), .imm_vec_ext_i(imm_vec_ext_i), .is_clpx_i(alu_is_clpx_i), 
        .is_subrot_i(alu_is_subrot_i), .clpx_shift_i(alu_clpx_shift_i), 
        .result_o(alu_result), .comparison_result_o(branch_decision_o), 
        .ready_o(alu_ready), .ex_ready_i(n172), .enable_i_BAR(alu_en_i_BAR) );
  riscv_mult_SHARED_DSP_MULT0 mult_i ( .clk(clk), .rst_n(rst_n), .enable_i(
        mult_en_i), .operator_i(mult_operator_i), .short_signed_i(
        mult_signed_mode_i), .op_a_i(mult_operand_a_i), .op_b_i(
        mult_operand_b_i), .op_c_i(mult_operand_c_i), .imm_i(mult_imm_i), 
        .dot_signed_i(mult_dot_signed_i), .dot_op_a_i(mult_dot_op_a_i), 
        .dot_op_b_i(mult_dot_op_b_i), .dot_op_c_i(mult_dot_op_c_i), 
        .is_clpx_i(mult_is_clpx_i), .clpx_shift_i(mult_clpx_shift_i), 
        .clpx_img_i(mult_clpx_img_i), .result_o(mult_result), .multicycle_o(
        mult_multicycle_o), .ready_o(mult_ready), .ex_ready_i(n172), 
        .short_subword_i_BAR(mult_sel_subword_i_BAR) );
  SNPS_CLOCK_GATE_HIGH_riscv_ex_stage_FPU0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_DIV0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_0 clk_gate_regfile_waddr_lsu_reg_0_ ( 
        .CLK(clk), .EN(n201), .ENCLK(n199), .TE(1'b0) );
  NAND2_X1 U5 ( .A1(n144), .A2(n143), .ZN(regfile_alu_wdata_fw_o[22]) );
  NAND2_X1 U8 ( .A1(n135), .A2(n134), .ZN(regfile_alu_wdata_fw_o[19]) );
  NAND2_X1 U20 ( .A1(n169), .A2(n168), .ZN(regfile_alu_wdata_fw_o[24]) );
  NAND2_X1 U9 ( .A1(n107), .A2(n106), .ZN(regfile_alu_wdata_fw_o[23]) );
  NAND2_X1 U18 ( .A1(n139), .A2(n138), .ZN(regfile_alu_wdata_fw_o[10]) );
  NAND2_X1 U16 ( .A1(n121), .A2(n120), .ZN(regfile_alu_wdata_fw_o[14]) );
  NAND2_X2 U19 ( .A1(n102), .A2(n91), .ZN(regfile_alu_wdata_fw_o[7]) );
  NAND2_X2 U4 ( .A1(n146), .A2(n145), .ZN(regfile_alu_wdata_fw_o[25]) );
  INV_X2 U3 ( .A(n103), .ZN(n184) );
  NAND2_X1 U6 ( .A1(n105), .A2(n104), .ZN(regfile_alu_wdata_fw_o[29]) );
  NAND2_X1 U10 ( .A1(n141), .A2(n140), .ZN(regfile_alu_wdata_fw_o[31]) );
  NAND3_X1 U11 ( .A1(n112), .A2(n111), .A3(n110), .ZN(
        regfile_alu_wdata_fw_o[6]) );
  CLKBUF_X1 U12 ( .A(n167), .Z(n163) );
  AOI22_X1 U13 ( .A1(mult_result[25]), .A2(n167), .B1(n185), .B2(
        csr_rdata_i[25]), .ZN(n145) );
  NAND2_X1 U14 ( .A1(n127), .A2(n126), .ZN(regfile_alu_wdata_fw_o[30]) );
  NAND2_X1 U17 ( .A1(n160), .A2(n159), .ZN(regfile_alu_wdata_fw_o[12]) );
  NAND2_X1 U21 ( .A1(n99), .A2(n100), .ZN(regfile_alu_wdata_fw_o[0]) );
  NAND2_X1 U22 ( .A1(n129), .A2(n128), .ZN(regfile_alu_wdata_fw_o[27]) );
  NAND2_X1 U23 ( .A1(n119), .A2(n118), .ZN(regfile_alu_wdata_fw_o[18]) );
  NAND2_X1 U24 ( .A1(n125), .A2(n124), .ZN(regfile_alu_wdata_fw_o[28]) );
  NAND2_X1 U26 ( .A1(n131), .A2(n130), .ZN(regfile_alu_wdata_fw_o[20]) );
  NAND2_X2 U31 ( .A1(n155), .A2(n154), .ZN(regfile_alu_wdata_fw_o[8]) );
  NAND2_X1 U32 ( .A1(n142), .A2(n94), .ZN(regfile_alu_wdata_fw_o[15]) );
  NAND2_X1 U36 ( .A1(n109), .A2(n108), .ZN(regfile_alu_wdata_fw_o[9]) );
  OR3_X1 U39 ( .A1(alu_en_i_BAR), .A2(n186), .A3(mult_en_i), .ZN(n103) );
  INV_X1 U56 ( .A(csr_access_i), .ZN(n185) );
  INV_X1 U95 ( .A(csr_access_i), .ZN(n186) );
  NAND2_X2 U120 ( .A1(n165), .A2(n164), .ZN(regfile_alu_wdata_fw_o[21]) );
  INV_X1 U134 ( .A(n170), .ZN(n201) );
endmodule



    module riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5 ( 
        clk, rst_n, test_en_i, fregfile_disable_i, fetch_enable_i, ctrl_busy_o, 
        core_ctrl_firstfetch_o, hwlp_dec_cnt_i, is_hwlp_i, instr_valid_i, 
        instr_rdata_i, instr_req_o, branch_in_ex_o, branch_decision_i, 
        jump_target_o, clear_instr_valid_o, pc_set_o, pc_mux_o, exc_pc_mux_o, 
        trap_addr_mux_o, illegal_c_insn_i, is_compressed_i, is_fetch_failed_i, 
        pc_if_i, pc_id_i, halt_if_o, ex_ready_i, wb_ready_i, id_valid_o, 
        ex_valid_i, pc_ex_o, alu_operand_a_ex_o, alu_operand_b_ex_o, 
        alu_operand_c_ex_o, bmask_a_ex_o, bmask_b_ex_o, imm_vec_ext_ex_o, 
        alu_vec_mode_ex_o, regfile_waddr_ex_o, regfile_we_ex_o, 
        regfile_alu_waddr_ex_o, alu_operator_ex_o, alu_is_clpx_ex_o, 
        alu_is_subrot_ex_o, alu_clpx_shift_ex_o, mult_operator_ex_o, 
        mult_operand_a_ex_o, mult_operand_b_ex_o, mult_operand_c_ex_o, 
        mult_en_ex_o, mult_signed_mode_ex_o, mult_imm_ex_o, mult_dot_op_a_ex_o, 
        mult_dot_op_b_ex_o, mult_dot_op_c_ex_o, mult_dot_signed_ex_o, 
        mult_is_clpx_ex_o, mult_clpx_shift_ex_o, mult_clpx_img_ex_o, 
        apu_en_ex_o, apu_type_ex_o, apu_op_ex_o, apu_lat_ex_o, 
        apu_operands_ex_o, apu_flags_ex_o, apu_waddr_ex_o, apu_read_regs_o, 
        apu_read_regs_valid_o, apu_read_dep_i, apu_write_regs_o, 
        apu_write_regs_valid_o, apu_write_dep_i, apu_perf_dep_o, apu_busy_i, 
        frm_i, csr_op_ex_o, current_priv_lvl_i, csr_irq_sec_o, csr_save_if_o, 
        csr_save_id_o, csr_restore_mret_id_o, csr_restore_uret_id_o, 
        csr_restore_dret_id_o, csr_save_cause_o, hwlp_start_o, hwlp_end_o, 
        hwlp_cnt_o, csr_hwlp_regid_i, csr_hwlp_we_i, csr_hwlp_data_i, 
        data_req_ex_o, data_we_ex_o, data_type_ex_o, data_sign_ext_ex_o, 
        data_reg_offset_ex_o, data_load_event_ex_o, data_misaligned_i, irq_i, 
        irq_sec_i, irq_id_i, m_irq_enable_i, u_irq_enable_i, irq_id_o, 
        exc_cause_o, debug_mode_o, debug_cause_o, debug_csr_save_o, 
        debug_req_i, debug_single_step_i, debug_ebreakm_i, debug_ebreaku_i, 
        regfile_waddr_wb_i, regfile_we_wb_i, regfile_wdata_wb_i, 
        regfile_alu_waddr_fw_i, regfile_alu_we_fw_i, regfile_alu_wdata_fw_i, 
        mult_multicycle_i, perf_jump_o, perf_jr_stall_o, perf_ld_stall_o, 
        perf_pipeline_stall_o, irq_ack_o_BAR, csr_cause_o_5__BAR, 
        csr_cause_o_4_, csr_cause_o_3_, csr_cause_o_2_, csr_cause_o_0_, 
        id_ready_o_BAR, data_err_ack_o_BAR, csr_save_ex_o_BAR, data_err_i_BAR, 
        regfile_alu_we_ex_o, alu_en_ex_o_BAR, mult_sel_subword_ex_o_BAR, 
        csr_cause_o_1__BAR, is_decoding_o, csr_access_ex_o_BAR, 
        data_misaligned_ex_o_BAR, prepost_useincr_ex_o );
  input [1:0] hwlp_dec_cnt_i;
  input [31:0] instr_rdata_i;
  output [31:0] jump_target_o;
  output [2:0] pc_mux_o;
  output [2:0] exc_pc_mux_o;
  input [31:0] pc_if_i;
  input [31:0] pc_id_i;
  output [31:0] pc_ex_o;
  output [31:0] alu_operand_a_ex_o;
  output [31:0] alu_operand_b_ex_o;
  output [31:0] alu_operand_c_ex_o;
  output [4:0] bmask_a_ex_o;
  output [4:0] bmask_b_ex_o;
  output [1:0] imm_vec_ext_ex_o;
  output [1:0] alu_vec_mode_ex_o;
  output [5:0] regfile_waddr_ex_o;
  output [5:0] regfile_alu_waddr_ex_o;
  output [6:0] alu_operator_ex_o;
  output [1:0] alu_clpx_shift_ex_o;
  output [2:0] mult_operator_ex_o;
  output [31:0] mult_operand_a_ex_o;
  output [31:0] mult_operand_b_ex_o;
  output [31:0] mult_operand_c_ex_o;
  output [1:0] mult_signed_mode_ex_o;
  output [4:0] mult_imm_ex_o;
  output [31:0] mult_dot_op_a_ex_o;
  output [31:0] mult_dot_op_b_ex_o;
  output [31:0] mult_dot_op_c_ex_o;
  output [1:0] mult_dot_signed_ex_o;
  output [1:0] mult_clpx_shift_ex_o;
  output [1:2] apu_type_ex_o;
  output [5:0] apu_op_ex_o;
  output [1:0] apu_lat_ex_o;
  output [95:0] apu_operands_ex_o;
  output [14:0] apu_flags_ex_o;
  output [5:0] apu_waddr_ex_o;
  output [17:0] apu_read_regs_o;
  output [2:0] apu_read_regs_valid_o;
  output [11:0] apu_write_regs_o;
  output [1:0] apu_write_regs_valid_o;
  input [2:0] frm_i;
  output [1:0] csr_op_ex_o;
  input [1:0] current_priv_lvl_i;
  output [63:0] hwlp_start_o;
  output [63:0] hwlp_end_o;
  output [63:0] hwlp_cnt_o;
  input [0:0] csr_hwlp_regid_i;
  input [2:0] csr_hwlp_we_i;
  input [31:0] csr_hwlp_data_i;
  output [1:0] data_type_ex_o;
  output [1:0] data_sign_ext_ex_o;
  output [1:0] data_reg_offset_ex_o;
  input [4:0] irq_id_i;
  output [4:0] irq_id_o;
  output [5:0] exc_cause_o;
  output [2:0] debug_cause_o;
  input [5:0] regfile_waddr_wb_i;
  input [31:0] regfile_wdata_wb_i;
  input [5:0] regfile_alu_waddr_fw_i;
  input [31:0] regfile_alu_wdata_fw_i;
  input clk, rst_n, test_en_i, fregfile_disable_i, fetch_enable_i, is_hwlp_i,
         instr_valid_i, branch_decision_i, illegal_c_insn_i, is_compressed_i,
         is_fetch_failed_i, ex_ready_i, wb_ready_i, ex_valid_i, apu_read_dep_i,
         apu_write_dep_i, apu_busy_i, data_misaligned_i, irq_i, irq_sec_i,
         m_irq_enable_i, u_irq_enable_i, debug_req_i, debug_single_step_i,
         debug_ebreakm_i, debug_ebreaku_i, regfile_we_wb_i,
         regfile_alu_we_fw_i, mult_multicycle_i, data_err_i_BAR;
  output ctrl_busy_o, core_ctrl_firstfetch_o, instr_req_o, branch_in_ex_o,
         clear_instr_valid_o, pc_set_o, trap_addr_mux_o, halt_if_o, id_valid_o,
         regfile_we_ex_o, alu_is_clpx_ex_o, alu_is_subrot_ex_o, mult_en_ex_o,
         mult_is_clpx_ex_o, mult_clpx_img_ex_o, apu_en_ex_o, apu_perf_dep_o,
         csr_irq_sec_o, csr_save_if_o, csr_save_id_o, csr_restore_mret_id_o,
         csr_restore_uret_id_o, csr_restore_dret_id_o, csr_save_cause_o,
         data_req_ex_o, data_we_ex_o, data_load_event_ex_o, debug_mode_o,
         debug_csr_save_o, perf_jump_o, perf_jr_stall_o, perf_ld_stall_o,
         perf_pipeline_stall_o, irq_ack_o_BAR, csr_cause_o_5__BAR,
         csr_cause_o_4_, csr_cause_o_3_, csr_cause_o_2_, csr_cause_o_0_,
         id_ready_o_BAR, data_err_ack_o_BAR, csr_save_ex_o_BAR,
         regfile_alu_we_ex_o, alu_en_ex_o_BAR, mult_sel_subword_ex_o_BAR,
         csr_cause_o_1__BAR, is_decoding_o, csr_access_ex_o_BAR,
         data_misaligned_ex_o_BAR, prepost_useincr_ex_o;
  wire   is_decoding_o_BAR, csr_access_ex_o, regfile_alu_waddr_mux_sel,
         rega_used_dec, reg_d_ex_is_reg_a_id, regb_used_dec,
         reg_d_ex_is_reg_b_id, regc_used_dec, reg_d_ex_is_reg_c_id,
         reg_d_wb_is_reg_a_id, reg_d_wb_is_reg_b_id, reg_d_wb_is_reg_c_id,
         reg_d_alu_is_reg_a_id, reg_d_alu_is_reg_b_id, reg_d_alu_is_reg_c_id,
         branch_taken_ex, mult_int_en, mult_dot_en, hwloop_start_mux_sel,
         hwloop_cnt_mux_sel, hwloop_regid_0_, imm_a_mux_sel_0_,
         scalar_replication, bmask_a_mux_0_, alu_bmask_a_mux_sel,
         alu_bmask_b_mux_sel, mult_imm_mux_0_, csr_access, deassert_we,
         illegal_insn_dec, mret_insn_dec, uret_insn_dec, dret_insn_dec,
         mret_dec, dret_dec, ecall_insn_dec, pipe_flush_dec, fencei_insn_dec,
         alu_en, is_clpx, is_subrot, mult_sel_subword, regfile_we_id,
         regfile_alu_we_id, regfile_alu_we_dec_id, csr_status, data_req_id,
         data_we_id, prepost_useincr, data_sign_ext_id_0_, data_load_event_id,
         irq_req_ctrl, irq_sec_ctrl, exc_ack, exc_kill, jr_stall, load_stall,
         hwloop_valid, n1276, n1352, n1353, n1626, n1634, n1635, n1636, n1637,
         n1638, n13, n16, n21, n22, n23, n24, n25, n31, n32, n33, n38, n44,
         n47, n48, n53, n55, n67, n68, n71, n72, n74, n75, n76, n77, n78, n79,
         n80, n90, n91, n94, n95, n96, n99, n100, n101, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n113, n114, n116, n117, n118, n119,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n168, n169,
         n171, n172, n173, n174, n175, n176, n177, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n627, n628, n629, n630, n631, n632,
         n634, n635, n636, n638, n640, n641, n642, n643, n646, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n778, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1328, n1396, n1632, n1633, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2434, n2435, n2448,
         n2451, n2452, n2453, n2455, n2456, n2457, n2458, n2459, n2462, n2463,
         n2467, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2480, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2517, n2518, n2519, n2520, n2521, n2523,
         n2524, n2525, n2526, n2527, n2528, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2577, n2597, n2599,
         n2604, n2627, n2631, n2644, n2645, n2647, n2648, n2649, n2650, n2651,
         n2652, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2678, n2681, n2682, n2683, n2684, n2685, n2686, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3481, n3483, n3484, n3486, n3487, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3506, n3507, n3509, n3510, n3511, n3512,
         n3513, n3515, n3517, n3518, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3540;
  wire   [1:0] regc_mux;
  wire   [4:0] regfile_alu_waddr_id;
  wire   [2:0] hwloop_we_int;
  wire   [31:0] hwloop_start;
  wire   [31:0] hwloop_end;
  wire   [31:0] hwloop_cnt;
  wire   [2:0] hwloop_we;
  wire   [1:0] jump_target_mux_sel;
  wire   [31:0] regfile_data_ra_id;
  wire   [2:0] alu_op_a_mux_sel;
  wire   [1:0] operand_a_fw_mux_sel;
  wire   [3:0] imm_b_mux_sel;
  wire   [2:0] alu_op_b_mux_sel;
  wire   [1:0] alu_vec_mode;
  wire   [1:0] operand_b_fw_mux_sel;
  wire   [31:0] regfile_data_rb_id;
  wire   [1:0] alu_op_c_mux_sel;
  wire   [1:0] operand_c_fw_mux_sel;
  wire   [31:0] regfile_data_rc_id;
  wire   [1:0] bmask_b_mux;
  wire   [6:0] alu_operator;
  wire   [2:0] mult_operator;
  wire   [1:0] mult_signed_mode;
  wire   [1:0] mult_dot_signed;
  wire   [1:0] csr_op;
  wire   [1:0] data_type_id;
  wire   [1:0] jump_in_dec;
  wire   [1:0] jump_in_id;
  wire   [4:0] irq_id_ctrl;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign is_decoding_o = is_decoding_o_BAR;
  assign data_reg_offset_ex_o[0] = 1'b0;
  assign data_reg_offset_ex_o[1] = 1'b0;
  assign data_sign_ext_ex_o[1] = 1'b0;
  assign apu_en_ex_o = 1'b0;
  assign regfile_alu_waddr_ex_o[5] = 1'b0;
  assign regfile_waddr_ex_o[5] = 1'b0;
  assign exc_pc_mux_o[2] = 1'b0;
  assign data_misaligned_ex_o_BAR = n2597;

  INV_X1 U15 ( .A(regfile_data_ra_id[16]), .ZN(n2274) );
  CLKBUF_X1 U16 ( .A(regfile_data_ra_id[11]), .Z(n25) );
  CLKBUF_X1 U17 ( .A(regfile_data_ra_id[8]), .Z(n24) );
  OAI21_X2 U18 ( .B1(n445), .B2(n334), .A(n333), .ZN(n368) );
  INV_X1 U19 ( .A(n90), .ZN(n23) );
  NAND2_X1 U26 ( .A1(n220), .A2(n79), .ZN(n246) );
  NAND2_X1 U27 ( .A1(n460), .A2(n327), .ZN(n446) );
  BUF_X1 U29 ( .A(n367), .Z(n399) );
  INV_X1 U30 ( .A(regfile_data_ra_id[19]), .ZN(n1933) );
  NAND2_X1 U31 ( .A1(n315), .A2(n13), .ZN(n325) );
  NAND2_X1 U32 ( .A1(regfile_data_ra_id[19]), .A2(n23), .ZN(n13) );
  NOR2_X2 U34 ( .A1(n224), .A2(n223), .ZN(n515) );
  NAND2_X1 U35 ( .A1(n310), .A2(n16), .ZN(n320) );
  NAND2_X1 U36 ( .A1(regfile_data_ra_id[16]), .A2(n23), .ZN(n16) );
  NOR2_X2 U39 ( .A1(n149), .A2(n266), .ZN(n562) );
  NAND2_X1 U40 ( .A1(n2062), .A2(n21), .ZN(n2510) );
  OR2_X1 U41 ( .A1(n2059), .A2(n1848), .ZN(n21) );
  NAND2_X1 U42 ( .A1(n302), .A2(n22), .ZN(n329) );
  NAND2_X1 U43 ( .A1(regfile_data_ra_id[20]), .A2(n23), .ZN(n22) );
  BUF_X1 U48 ( .A(regfile_data_ra_id[6]), .Z(n32) );
  BUF_X1 U49 ( .A(instr_rdata_i[18]), .Z(n33) );
  INV_X1 U53 ( .A(n2274), .ZN(n38) );
  NOR2_X2 U55 ( .A1(n495), .A2(n501), .ZN(n487) );
  NOR2_X2 U56 ( .A1(n440), .A2(n434), .ZN(n426) );
  AND2_X1 U60 ( .A1(n2209), .A2(n1130), .ZN(n1195) );
  OR2_X1 U62 ( .A1(n2126), .A2(n1848), .ZN(n44) );
  NOR2_X1 U73 ( .A1(n490), .A2(n481), .ZN(n243) );
  AND2_X1 U74 ( .A1(scalar_replication), .A2(n1732), .ZN(n1848) );
  BUF_X1 U79 ( .A(instr_rdata_i[15]), .Z(n113) );
  BUF_X1 U80 ( .A(instr_rdata_i[31]), .Z(n352) );
  AND2_X1 U83 ( .A1(n2011), .A2(n2010), .ZN(n75) );
  AOI21_X1 U86 ( .B1(regfile_alu_wdata_fw_i[8]), .B2(n2205), .A(n632), .ZN(
        n2198) );
  INV_X2 U94 ( .A(n94), .ZN(n53) );
  NOR2_X1 U95 ( .A1(hwloop_start_mux_sel), .A2(n211), .ZN(n995) );
  AND2_X1 U96 ( .A1(n1939), .A2(n1937), .ZN(n71) );
  NOR2_X2 U100 ( .A1(n1901), .A2(n1900), .ZN(n2084) );
  BUF_X1 U101 ( .A(n367), .Z(n584) );
  NOR2_X1 U102 ( .A1(n515), .A2(n511), .ZN(n247) );
  OR2_X1 U103 ( .A1(regc_mux[1]), .A2(regc_mux[0]), .ZN(n743) );
  NOR2_X1 U104 ( .A1(n222), .A2(instr_rdata_i[30]), .ZN(n511) );
  AND2_X1 U105 ( .A1(n78), .A2(n76), .ZN(n528) );
  AND3_X1 U106 ( .A1(n121), .A2(n229), .A3(n120), .ZN(n501) );
  AND3_X1 U107 ( .A1(n119), .A2(n226), .A3(n118), .ZN(n495) );
  CLKBUF_X1 U108 ( .A(regfile_data_ra_id[0]), .Z(n114) );
  AND2_X1 U109 ( .A1(regfile_data_ra_id[17]), .A2(n23), .ZN(n104) );
  INV_X1 U110 ( .A(regfile_data_ra_id[17]), .ZN(n1888) );
  INV_X1 U111 ( .A(alu_op_b_mux_sel[2]), .ZN(n1853) );
  NOR2_X1 U112 ( .A1(n77), .A2(instr_rdata_i[29]), .ZN(n76) );
  INV_X1 U113 ( .A(n160), .ZN(n77) );
  OR2_X1 U117 ( .A1(jump_target_mux_sel[1]), .A2(n215), .ZN(n318) );
  NAND2_X1 U118 ( .A1(n247), .A2(n520), .ZN(n506) );
  NAND2_X1 U119 ( .A1(n2664), .A2(n44), .ZN(n2514) );
  NAND3_X1 U121 ( .A1(n2062), .A2(n2060), .A3(n2061), .ZN(n2527) );
  NAND2_X1 U122 ( .A1(n1925), .A2(n1848), .ZN(n2062) );
  NAND2_X1 U123 ( .A1(n68), .A2(n67), .ZN(n149) );
  NAND2_X1 U124 ( .A1(n277), .A2(pc_id_i[3]), .ZN(n67) );
  NAND2_X1 U125 ( .A1(regfile_data_ra_id[3]), .A2(n23), .ZN(n68) );
  NAND3_X1 U126 ( .A1(n1938), .A2(n72), .A3(n71), .ZN(n2519) );
  NAND2_X1 U127 ( .A1(n1925), .A2(scalar_replication), .ZN(n72) );
  NOR2_X1 U130 ( .A1(n328), .A2(n352), .ZN(n440) );
  NAND3_X1 U131 ( .A1(n74), .A2(n2013), .A3(n75), .ZN(n2525) );
  NAND2_X1 U132 ( .A1(n2012), .A2(n2033), .ZN(n74) );
  OAI21_X1 U133 ( .B1(n580), .B2(n402), .A(n401), .ZN(n407) );
  AND2_X4 U134 ( .A1(n290), .A2(n289), .ZN(n580) );
  NAND2_X1 U135 ( .A1(n246), .A2(n2668), .ZN(n597) );
  NAND2_X1 U136 ( .A1(n78), .A2(n160), .ZN(n221) );
  NAND2_X1 U137 ( .A1(regfile_data_ra_id[9]), .A2(n23), .ZN(n78) );
  NAND2_X1 U138 ( .A1(regfile_data_ra_id[8]), .A2(n23), .ZN(n79) );
  INV_X2 U143 ( .A(instr_rdata_i[24]), .ZN(n1904) );
  INV_X1 U145 ( .A(n55), .ZN(n91) );
  NOR2_X1 U146 ( .A1(n596), .A2(n528), .ZN(n520) );
  INV_X1 U147 ( .A(n311), .ZN(n317) );
  OAI21_X1 U148 ( .B1(n2673), .B2(n738), .A(n227), .ZN(n311) );
  NOR2_X1 U149 ( .A1(n1863), .A2(n154), .ZN(n153) );
  INV_X1 U150 ( .A(regfile_data_ra_id[13]), .ZN(n154) );
  AOI21_X1 U151 ( .B1(n1038), .B2(n146), .A(n1779), .ZN(n145) );
  INV_X1 U152 ( .A(n1228), .ZN(n146) );
  AOI21_X1 U153 ( .B1(n1036), .B2(n1882), .A(n1684), .ZN(n142) );
  AOI21_X1 U154 ( .B1(n135), .B2(n1865), .A(n1719), .ZN(n127) );
  AND2_X1 U155 ( .A1(n132), .A2(n604), .ZN(n124) );
  INV_X1 U156 ( .A(n133), .ZN(n132) );
  OAI21_X1 U157 ( .B1(n604), .B2(n2205), .A(n134), .ZN(n133) );
  INV_X1 U158 ( .A(n31), .ZN(n1727) );
  OR2_X1 U162 ( .A1(n2148), .A2(n1684), .ZN(n172) );
  AOI21_X1 U163 ( .B1(regfile_alu_wdata_fw_i[9]), .B2(n2205), .A(n636), .ZN(
        n2204) );
  OAI211_X1 U164 ( .C1(n2106), .C2(n2125), .A(n2105), .B(n2107), .ZN(n2531) );
  OR2_X1 U165 ( .A1(n2126), .A2(n2125), .ZN(n151) );
  NOR2_X1 U166 ( .A1(n158), .A2(n157), .ZN(n159) );
  INV_X1 U167 ( .A(n2455), .ZN(n157) );
  INV_X1 U168 ( .A(n2671), .ZN(n158) );
  INV_X1 U169 ( .A(n234), .ZN(n118) );
  INV_X1 U170 ( .A(pc_id_i[9]), .ZN(n161) );
  INV_X1 U172 ( .A(n236), .ZN(n120) );
  NOR2_X1 U173 ( .A1(n1863), .A2(n137), .ZN(n1796) );
  INV_X1 U174 ( .A(n1038), .ZN(n147) );
  INV_X1 U175 ( .A(n1036), .ZN(n143) );
  NOR2_X1 U176 ( .A1(n95), .A2(n153), .ZN(n152) );
  AND2_X1 U177 ( .A1(regfile_wdata_wb_i[6]), .A2(n2179), .ZN(n135) );
  OAI21_X1 U178 ( .B1(n580), .B2(n576), .A(n577), .ZN(n472) );
  NOR2_X1 U179 ( .A1(n282), .A2(instr_rdata_i[25]), .ZN(n552) );
  INV_X1 U180 ( .A(regfile_data_ra_id[12]), .ZN(n1806) );
  OAI21_X1 U181 ( .B1(n838), .B2(n205), .A(n204), .ZN(n840) );
  NOR2_X1 U182 ( .A1(n862), .A2(n206), .ZN(n864) );
  NOR2_X1 U183 ( .A1(n873), .A2(n207), .ZN(n875) );
  INV_X1 U184 ( .A(pc_id_i[27]), .ZN(n888) );
  XNOR2_X1 U185 ( .A(n891), .B(pc_id_i[28]), .ZN(n991) );
  NOR2_X1 U186 ( .A1(n891), .A2(n209), .ZN(n893) );
  AND2_X1 U187 ( .A1(n1101), .A2(n1103), .ZN(n1073) );
  CLKBUF_X1 U188 ( .A(branch_taken_ex), .Z(n185) );
  AND2_X1 U189 ( .A1(n684), .A2(n156), .ZN(n155) );
  AOI21_X1 U190 ( .B1(regfile_alu_wdata_fw_i[0]), .B2(n99), .A(n138), .ZN(n148) );
  OR2_X1 U191 ( .A1(n129), .A2(n132), .ZN(n125) );
  OR2_X1 U192 ( .A1(n126), .A2(n124), .ZN(n123) );
  INV_X1 U198 ( .A(n1779), .ZN(n131) );
  OR2_X1 U199 ( .A1(n719), .A2(n2130), .ZN(n94) );
  INV_X2 U200 ( .A(hwloop_we_int[2]), .ZN(n615) );
  AND2_X1 U201 ( .A1(n1860), .A2(instr_rdata_i[13]), .ZN(n95) );
  OR2_X1 U202 ( .A1(n2092), .A2(n1848), .ZN(n96) );
  OR2_X1 U206 ( .A1(n145), .A2(n142), .ZN(n99) );
  INV_X1 U207 ( .A(n173), .ZN(n171) );
  NAND2_X1 U208 ( .A1(n1924), .A2(n1922), .ZN(n173) );
  AND2_X1 U209 ( .A1(n184), .A2(n2455), .ZN(n100) );
  OR2_X1 U210 ( .A1(n1798), .A2(n2177), .ZN(n101) );
  OAI21_X1 U211 ( .B1(n104), .B2(n103), .A(n321), .ZN(n469) );
  INV_X1 U212 ( .A(n313), .ZN(n103) );
  NOR2_X1 U213 ( .A1(n105), .A2(n104), .ZN(n468) );
  NAND2_X1 U214 ( .A1(n313), .A2(n106), .ZN(n105) );
  INV_X1 U215 ( .A(n321), .ZN(n106) );
  OAI211_X2 U216 ( .C1(n743), .C2(n735), .A(n734), .B(n733), .ZN(n1637) );
  OAI211_X2 U217 ( .C1(n2431), .C2(n743), .A(n730), .B(n729), .ZN(n1636) );
  INV_X1 U218 ( .A(n1881), .ZN(n134) );
  INV_X2 U219 ( .A(n1103), .ZN(n1194) );
  INV_X2 U220 ( .A(n2273), .ZN(n2410) );
  NAND2_X1 U222 ( .A1(n286), .A2(n544), .ZN(n108) );
  NAND2_X1 U223 ( .A1(n109), .A2(n278), .ZN(n284) );
  NAND2_X1 U224 ( .A1(regfile_data_ra_id[7]), .A2(n23), .ZN(n109) );
  NAND2_X1 U225 ( .A1(n275), .A2(n111), .ZN(n282) );
  NAND2_X1 U226 ( .A1(regfile_data_ra_id[5]), .A2(n23), .ZN(n111) );
  OR2_X1 U229 ( .A1(n292), .A2(n161), .ZN(n160) );
  OAI21_X1 U230 ( .B1(n1042), .B2(n572), .A(n573), .ZN(n561) );
  NAND2_X1 U231 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  INV_X2 U232 ( .A(n1904), .ZN(n2604) );
  NAND2_X1 U233 ( .A1(n117), .A2(n96), .ZN(n2512) );
  NAND2_X1 U234 ( .A1(n117), .A2(n2094), .ZN(n2530) );
  NAND2_X1 U235 ( .A1(n1971), .A2(n1848), .ZN(n117) );
  NAND2_X1 U236 ( .A1(n119), .A2(n226), .ZN(n235) );
  NAND2_X1 U237 ( .A1(regfile_data_ra_id[12]), .A2(n215), .ZN(n119) );
  NAND2_X1 U238 ( .A1(n121), .A2(n229), .ZN(n237) );
  NAND2_X1 U239 ( .A1(regfile_data_ra_id[13]), .A2(n23), .ZN(n121) );
  AOI21_X1 U241 ( .B1(regfile_alu_wdata_fw_i[6]), .B2(n125), .A(n123), .ZN(
        n1822) );
  AOI21_X1 U242 ( .B1(regfile_alu_wdata_fw_i[6]), .B2(n1228), .A(n1072), .ZN(
        n2176) );
  AOI21_X1 U243 ( .B1(regfile_alu_wdata_fw_i[6]), .B2(n1879), .A(n135), .ZN(
        n2171) );
  AOI21_X1 U244 ( .B1(regfile_alu_wdata_fw_i[6]), .B2(n2205), .A(n604), .ZN(
        n2173) );
  NAND2_X1 U245 ( .A1(n128), .A2(n127), .ZN(n126) );
  NAND2_X1 U246 ( .A1(n1072), .A2(n131), .ZN(n128) );
  NAND2_X1 U247 ( .A1(n130), .A2(n101), .ZN(n129) );
  NAND2_X1 U248 ( .A1(n1228), .A2(n131), .ZN(n130) );
  NAND2_X1 U249 ( .A1(n136), .A2(n217), .ZN(n224) );
  NAND2_X1 U250 ( .A1(regfile_data_ra_id[11]), .A2(n23), .ZN(n136) );
  INV_X1 U251 ( .A(n25), .ZN(n137) );
  NAND3_X1 U252 ( .A1(n140), .A2(n139), .A3(n1225), .ZN(n138) );
  NAND2_X1 U253 ( .A1(n142), .A2(n143), .ZN(n139) );
  NAND2_X1 U254 ( .A1(n145), .A2(n147), .ZN(n140) );
  NAND2_X1 U255 ( .A1(n141), .A2(n1036), .ZN(n1205) );
  NAND2_X1 U256 ( .A1(regfile_alu_wdata_fw_i[0]), .A2(n2205), .ZN(n141) );
  NAND2_X1 U257 ( .A1(n144), .A2(n1038), .ZN(n1206) );
  NAND2_X1 U258 ( .A1(regfile_alu_wdata_fw_i[0]), .A2(n1228), .ZN(n144) );
  NAND2_X1 U259 ( .A1(n1226), .A2(n148), .ZN(n1872) );
  NAND2_X1 U260 ( .A1(n149), .A2(n266), .ZN(n563) );
  NAND3_X1 U264 ( .A1(n2124), .A2(n2123), .A3(n151), .ZN(n150) );
  NAND2_X1 U265 ( .A1(n1816), .A2(n152), .ZN(n1817) );
  NAND2_X1 U266 ( .A1(n685), .A2(n155), .ZN(hwloop_cnt[13]) );
  NAND2_X1 U267 ( .A1(n53), .A2(regfile_data_ra_id[13]), .ZN(n156) );
  NAND2_X1 U268 ( .A1(ex_ready_i), .A2(n100), .ZN(id_ready_o_BAR) );
  NAND2_X1 U269 ( .A1(n159), .A2(n2434), .ZN(n810) );
  INV_X1 U270 ( .A(regfile_data_ra_id[9]), .ZN(n1754) );
  NAND2_X1 U271 ( .A1(n215), .A2(n352), .ZN(n227) );
  NAND3_X1 U275 ( .A1(n2048), .A2(n2046), .A3(n2047), .ZN(n162) );
  AND2_X1 U276 ( .A1(n1923), .A2(n171), .ZN(n169) );
  NAND2_X1 U278 ( .A1(n169), .A2(n168), .ZN(n2518) );
  NAND2_X1 U279 ( .A1(n1912), .A2(scalar_replication), .ZN(n168) );
  NAND2_X1 U280 ( .A1(n1653), .A2(n172), .ZN(n1912) );
  AOI21_X1 U281 ( .B1(regfile_alu_wdata_fw_i[2]), .B2(n1228), .A(n1054), .ZN(
        n1647) );
  OR2_X1 U282 ( .A1(n1005), .A2(n212), .ZN(n174) );
  OR2_X1 U283 ( .A1(n1202), .A2(n1884), .ZN(n175) );
  INV_X1 U284 ( .A(pc_id_i[28]), .ZN(n209) );
  AND2_X1 U285 ( .A1(n831), .A2(pc_id_i[6]), .ZN(n176) );
  OR2_X1 U286 ( .A1(n831), .A2(pc_id_i[6]), .ZN(n177) );
  AND2_X1 U287 ( .A1(n213), .A2(n174), .ZN(n179) );
  AND2_X1 U288 ( .A1(n1948), .A2(n1947), .ZN(n180) );
  OR2_X1 U289 ( .A1(n2063), .A2(n1848), .ZN(n181) );
  OR2_X1 U290 ( .A1(n2045), .A2(n1848), .ZN(n182) );
  OR2_X1 U291 ( .A1(n2106), .A2(n1848), .ZN(n183) );
  OR2_X1 U292 ( .A1(n191), .A2(n190), .ZN(n192) );
  OR2_X1 U293 ( .A1(n821), .A2(pc_id_i[3]), .ZN(n201) );
  INV_X1 U294 ( .A(pc_id_i[7]), .ZN(n835) );
  OR2_X1 U295 ( .A1(n1849), .A2(n1884), .ZN(n1850) );
  XNOR2_X1 U296 ( .A(n821), .B(pc_id_i[3]), .ZN(n822) );
  AOI21_X1 U297 ( .B1(n833), .B2(n177), .A(n176), .ZN(n838) );
  NOR2_X1 U298 ( .A1(n882), .A2(n208), .ZN(n884) );
  XNOR2_X1 U299 ( .A(n859), .B(n858), .ZN(n940) );
  XNOR2_X1 U300 ( .A(n880), .B(n879), .ZN(n971) );
  OR2_X1 U301 ( .A1(n2427), .A2(n186), .ZN(n605) );
  OR2_X1 U302 ( .A1(n2161), .A2(n1684), .ZN(n1667) );
  OR2_X1 U303 ( .A1(n1685), .A2(n1684), .ZN(n1686) );
  NAND2_X1 U304 ( .A1(n2205), .A2(n2269), .ZN(n2424) );
  INV_X1 U305 ( .A(mult_multicycle_i), .ZN(n2434) );
  INV_X1 U306 ( .A(n2427), .ZN(n1032) );
  NAND2_X1 U307 ( .A1(id_valid_o), .A2(n2434), .ZN(n2427) );
  NOR2_X1 U308 ( .A1(n2577), .A2(n91), .ZN(id_valid_o) );
  INV_X1 U309 ( .A(data_misaligned_i), .ZN(n2455) );
  NOR2_X1 U310 ( .A1(load_stall), .A2(jr_stall), .ZN(n184) );
  AND2_X1 U311 ( .A1(branch_decision_i), .A2(branch_in_ex_o), .ZN(
        branch_taken_ex) );
  NOR2_X1 U312 ( .A1(n185), .A2(alu_en), .ZN(n186) );
  NOR2_X1 U314 ( .A1(id_valid_o), .A2(n810), .ZN(n187) );
  AOI21_X1 U317 ( .B1(n1032), .B2(n185), .A(n187), .ZN(n2448) );
  INV_X1 U321 ( .A(instr_rdata_i[17]), .ZN(n770) );
  INV_X1 U322 ( .A(n113), .ZN(n768) );
  INV_X1 U323 ( .A(n80), .ZN(n1008) );
  NAND3_X1 U324 ( .A1(n770), .A2(n768), .A3(n1008), .ZN(n191) );
  INV_X1 U325 ( .A(n33), .ZN(n1914) );
  INV_X1 U326 ( .A(n116), .ZN(n1010) );
  NAND2_X1 U327 ( .A1(n1914), .A2(n1010), .ZN(n190) );
  NAND2_X1 U328 ( .A1(rega_used_dec), .A2(n192), .ZN(n809) );
  XOR2_X1 U329 ( .A(n110), .B(regfile_waddr_ex_o[2]), .Z(n195) );
  XOR2_X1 U330 ( .A(n33), .B(regfile_waddr_ex_o[3]), .Z(n194) );
  XOR2_X1 U331 ( .A(n113), .B(regfile_waddr_ex_o[0]), .Z(n193) );
  NOR3_X1 U332 ( .A1(n195), .A2(n194), .A3(n193), .ZN(n198) );
  XNOR2_X1 U333 ( .A(regfile_waddr_ex_o[4]), .B(n116), .ZN(n197) );
  XNOR2_X1 U334 ( .A(regfile_waddr_ex_o[1]), .B(n80), .ZN(n196) );
  NAND3_X1 U335 ( .A1(n198), .A2(n197), .A3(n196), .ZN(n199) );
  NOR2_X1 U336 ( .A1(n809), .A2(n199), .ZN(reg_d_ex_is_reg_a_id) );
  INV_X1 U337 ( .A(instr_rdata_i[31]), .ZN(n738) );
  NOR2_X1 U338 ( .A1(n2631), .A2(n738), .ZN(n853) );
  INV_X1 U339 ( .A(instr_rdata_i[30]), .ZN(n735) );
  NOR2_X1 U340 ( .A1(n2631), .A2(n735), .ZN(n850) );
  INV_X1 U341 ( .A(instr_rdata_i[29]), .ZN(n2431) );
  NOR2_X1 U342 ( .A1(n2631), .A2(n2431), .ZN(n847) );
  INV_X1 U343 ( .A(n2668), .ZN(n2430) );
  NOR2_X1 U344 ( .A1(n2631), .A2(n2430), .ZN(n844) );
  INV_X1 U345 ( .A(n2678), .ZN(n2429) );
  NOR2_X1 U346 ( .A1(n2631), .A2(n2429), .ZN(n841) );
  OAI22_X1 U348 ( .A1(n2657), .A2(n1010), .B1(n2631), .B2(n1904), .ZN(n829) );
  INV_X1 U349 ( .A(instr_rdata_i[23]), .ZN(n1991) );
  OAI22_X1 U350 ( .A1(n2657), .A2(n1914), .B1(n2631), .B2(n1991), .ZN(n826) );
  INV_X1 U351 ( .A(instr_rdata_i[21]), .ZN(n1738) );
  OAI22_X1 U352 ( .A1(n2657), .A2(n1008), .B1(n2631), .B2(n1738), .ZN(n819) );
  INV_X1 U353 ( .A(instr_rdata_i[20]), .ZN(n2467) );
  OAI22_X1 U354 ( .A1(n2657), .A2(n768), .B1(n2631), .B2(n2467), .ZN(n816) );
  AND2_X1 U355 ( .A1(pc_id_i[1]), .A2(n816), .ZN(n818) );
  INV_X1 U356 ( .A(instr_rdata_i[22]), .ZN(n1984) );
  OAI22_X1 U357 ( .A1(n2657), .A2(n770), .B1(n2631), .B2(n1984), .ZN(n821) );
  NAND2_X1 U358 ( .A1(n823), .A2(n201), .ZN(n203) );
  NAND2_X1 U359 ( .A1(n821), .A2(pc_id_i[3]), .ZN(n202) );
  NAND2_X1 U360 ( .A1(n203), .A2(n202), .ZN(n825) );
  INV_X1 U361 ( .A(instr_rdata_i[25]), .ZN(n2463) );
  NOR2_X1 U362 ( .A1(n2631), .A2(n2463), .ZN(n831) );
  INV_X1 U363 ( .A(instr_rdata_i[26]), .ZN(n2428) );
  NOR2_X1 U364 ( .A1(n2631), .A2(n2428), .ZN(n836) );
  NOR2_X1 U365 ( .A1(n836), .A2(pc_id_i[7]), .ZN(n205) );
  NAND2_X1 U366 ( .A1(n836), .A2(pc_id_i[7]), .ZN(n204) );
  NAND2_X1 U367 ( .A1(n859), .A2(pc_id_i[14]), .ZN(n862) );
  INV_X1 U368 ( .A(pc_id_i[15]), .ZN(n206) );
  NAND2_X1 U369 ( .A1(n871), .A2(pc_id_i[19]), .ZN(n873) );
  INV_X1 U370 ( .A(pc_id_i[20]), .ZN(n207) );
  NAND2_X1 U371 ( .A1(n880), .A2(pc_id_i[23]), .ZN(n882) );
  INV_X1 U372 ( .A(pc_id_i[24]), .ZN(n208) );
  NAND2_X1 U373 ( .A1(n889), .A2(pc_id_i[27]), .ZN(n891) );
  XOR2_X1 U374 ( .A(n210), .B(pc_id_i[31]), .Z(n898) );
  INV_X1 U375 ( .A(hwloop_we_int[0]), .ZN(n211) );
  NAND2_X1 U376 ( .A1(n2659), .A2(n1000), .ZN(n214) );
  NAND2_X1 U377 ( .A1(n900), .A2(pc_if_i[31]), .ZN(n213) );
  INV_X1 U379 ( .A(csr_hwlp_data_i[31]), .ZN(n212) );
  NAND2_X1 U380 ( .A1(n214), .A2(n179), .ZN(hwloop_start[31]) );
  INV_X1 U381 ( .A(n47), .ZN(n1773) );
  INV_X1 U382 ( .A(jump_target_mux_sel[0]), .ZN(n215) );
  NAND2_X1 U384 ( .A1(n277), .A2(pc_id_i[10]), .ZN(n216) );
  OAI21_X1 U385 ( .B1(n1773), .B2(n90), .A(n216), .ZN(n222) );
  NAND2_X1 U386 ( .A1(n277), .A2(pc_id_i[11]), .ZN(n217) );
  INV_X1 U387 ( .A(instr_rdata_i[7]), .ZN(n1216) );
  INV_X1 U388 ( .A(n48), .ZN(n218) );
  NAND2_X1 U389 ( .A1(n218), .A2(instr_rdata_i[20]), .ZN(n219) );
  OAI211_X1 U390 ( .C1(n2673), .C2(n1216), .A(n219), .B(n227), .ZN(n223) );
  NAND2_X1 U391 ( .A1(n277), .A2(pc_id_i[8]), .ZN(n220) );
  NAND2_X1 U392 ( .A1(n221), .A2(instr_rdata_i[29]), .ZN(n529) );
  NAND2_X1 U393 ( .A1(n222), .A2(instr_rdata_i[30]), .ZN(n524) );
  NAND2_X1 U394 ( .A1(n224), .A2(n223), .ZN(n516) );
  OAI21_X1 U395 ( .B1(n515), .B2(n524), .A(n516), .ZN(n225) );
  AOI21_X1 U396 ( .B1(n521), .B2(n247), .A(n225), .ZN(n475) );
  NAND2_X1 U397 ( .A1(n349), .A2(pc_id_i[12]), .ZN(n226) );
  INV_X1 U398 ( .A(instr_rdata_i[12]), .ZN(n228) );
  OAI21_X1 U399 ( .B1(n228), .B2(n48), .A(n2669), .ZN(n234) );
  NAND2_X1 U400 ( .A1(n349), .A2(pc_id_i[13]), .ZN(n229) );
  INV_X1 U401 ( .A(instr_rdata_i[13]), .ZN(n230) );
  OAI21_X1 U402 ( .B1(n230), .B2(n48), .A(n317), .ZN(n236) );
  INV_X1 U403 ( .A(regfile_data_ra_id[14]), .ZN(n1828) );
  NAND2_X1 U404 ( .A1(n349), .A2(pc_id_i[14]), .ZN(n231) );
  OAI21_X1 U405 ( .B1(n1828), .B2(n90), .A(n231), .ZN(n239) );
  INV_X1 U406 ( .A(instr_rdata_i[14]), .ZN(n232) );
  OAI21_X1 U407 ( .B1(n232), .B2(n48), .A(n2669), .ZN(n238) );
  INV_X1 U409 ( .A(regfile_data_ra_id[15]), .ZN(n1840) );
  INV_X2 U410 ( .A(n292), .ZN(n349) );
  NAND2_X1 U411 ( .A1(n349), .A2(pc_id_i[15]), .ZN(n233) );
  OAI21_X1 U412 ( .B1(n1840), .B2(n90), .A(n233), .ZN(n241) );
  OAI21_X1 U413 ( .B1(n768), .B2(n48), .A(n2669), .ZN(n240) );
  NOR2_X1 U414 ( .A1(n241), .A2(n240), .ZN(n481) );
  NAND2_X1 U415 ( .A1(n487), .A2(n243), .ZN(n248) );
  NAND2_X1 U416 ( .A1(n235), .A2(n234), .ZN(n507) );
  NAND2_X1 U417 ( .A1(n237), .A2(n236), .ZN(n502) );
  OAI21_X1 U418 ( .B1(n501), .B2(n507), .A(n502), .ZN(n486) );
  NAND2_X1 U419 ( .A1(n239), .A2(n238), .ZN(n491) );
  NAND2_X1 U420 ( .A1(n241), .A2(n240), .ZN(n482) );
  OAI21_X1 U421 ( .B1(n481), .B2(n491), .A(n482), .ZN(n242) );
  AOI21_X1 U422 ( .B1(n243), .B2(n486), .A(n242), .ZN(n244) );
  OAI21_X1 U423 ( .B1(n475), .B2(n248), .A(n244), .ZN(n245) );
  INV_X1 U424 ( .A(n245), .ZN(n290) );
  NOR2_X1 U425 ( .A1(n246), .A2(n2668), .ZN(n596) );
  NOR2_X1 U426 ( .A1(n506), .A2(n248), .ZN(n288) );
  INV_X1 U427 ( .A(regfile_data_ra_id[2]), .ZN(n2152) );
  NAND2_X1 U428 ( .A1(n277), .A2(pc_id_i[2]), .ZN(n249) );
  OAI21_X1 U429 ( .B1(n2152), .B2(n90), .A(n249), .ZN(n265) );
  NOR2_X1 U430 ( .A1(n48), .A2(n1984), .ZN(n252) );
  INV_X1 U431 ( .A(instr_rdata_i[9]), .ZN(n250) );
  OAI22_X1 U432 ( .A1(n2673), .A2(n250), .B1(n90), .B2(n1984), .ZN(n251) );
  OR2_X1 U433 ( .A1(n252), .A2(n251), .ZN(n264) );
  NOR2_X1 U434 ( .A1(n265), .A2(n264), .ZN(n567) );
  NOR2_X1 U435 ( .A1(n48), .A2(n1991), .ZN(n255) );
  INV_X1 U436 ( .A(instr_rdata_i[10]), .ZN(n253) );
  OAI22_X1 U437 ( .A1(n2673), .A2(n253), .B1(n90), .B2(n1991), .ZN(n254) );
  OR2_X1 U438 ( .A1(n255), .A2(n254), .ZN(n266) );
  NOR2_X1 U439 ( .A1(n567), .A2(n562), .ZN(n268) );
  INV_X1 U440 ( .A(regfile_data_ra_id[1]), .ZN(n257) );
  NAND2_X1 U441 ( .A1(n277), .A2(pc_id_i[1]), .ZN(n256) );
  OAI21_X1 U442 ( .B1(n257), .B2(n90), .A(n256), .ZN(n263) );
  NOR2_X1 U443 ( .A1(n48), .A2(n1738), .ZN(n260) );
  INV_X1 U444 ( .A(instr_rdata_i[8]), .ZN(n258) );
  OAI22_X1 U445 ( .A1(n2673), .A2(n258), .B1(n90), .B2(n1738), .ZN(n259) );
  OR2_X1 U446 ( .A1(n260), .A2(n259), .ZN(n262) );
  NOR2_X1 U447 ( .A1(n263), .A2(n262), .ZN(n572) );
  INV_X1 U448 ( .A(regfile_data_ra_id[0]), .ZN(n2134) );
  NAND2_X1 U449 ( .A1(n277), .A2(pc_id_i[0]), .ZN(n261) );
  OAI21_X1 U450 ( .B1(n2134), .B2(n90), .A(n261), .ZN(n1041) );
  NOR2_X1 U451 ( .A1(n90), .A2(n2467), .ZN(n1040) );
  NAND2_X1 U452 ( .A1(n263), .A2(n262), .ZN(n573) );
  NAND2_X1 U453 ( .A1(n265), .A2(n264), .ZN(n568) );
  OAI21_X1 U454 ( .B1(n562), .B2(n568), .A(n563), .ZN(n267) );
  AOI21_X1 U455 ( .B1(n268), .B2(n561), .A(n267), .ZN(n534) );
  INV_X1 U456 ( .A(regfile_data_ra_id[4]), .ZN(n270) );
  NAND2_X1 U457 ( .A1(n277), .A2(pc_id_i[4]), .ZN(n269) );
  OAI21_X1 U458 ( .B1(n270), .B2(n90), .A(n269), .ZN(n281) );
  NOR2_X1 U459 ( .A1(n48), .A2(n1904), .ZN(n274) );
  INV_X1 U460 ( .A(instr_rdata_i[11]), .ZN(n271) );
  OAI22_X1 U461 ( .A1(n2673), .A2(n271), .B1(n90), .B2(n1904), .ZN(n273) );
  OR2_X1 U462 ( .A1(n274), .A2(n273), .ZN(n280) );
  NOR2_X1 U463 ( .A1(n281), .A2(n280), .ZN(n550) );
  NAND2_X1 U464 ( .A1(n277), .A2(pc_id_i[5]), .ZN(n275) );
  NOR2_X1 U465 ( .A1(n550), .A2(n552), .ZN(n544) );
  INV_X1 U466 ( .A(regfile_data_ra_id[6]), .ZN(n1718) );
  NAND2_X1 U467 ( .A1(n277), .A2(pc_id_i[6]), .ZN(n276) );
  OAI21_X1 U468 ( .B1(n1718), .B2(n90), .A(n276), .ZN(n283) );
  NOR2_X1 U469 ( .A1(n283), .A2(instr_rdata_i[26]), .ZN(n545) );
  NAND2_X1 U470 ( .A1(n277), .A2(pc_id_i[7]), .ZN(n278) );
  NOR2_X1 U471 ( .A1(n284), .A2(n2678), .ZN(n538) );
  NOR2_X1 U472 ( .A1(n545), .A2(n538), .ZN(n286) );
  NAND2_X1 U473 ( .A1(n281), .A2(n280), .ZN(n557) );
  NAND2_X1 U474 ( .A1(n282), .A2(instr_rdata_i[25]), .ZN(n553) );
  OAI21_X1 U475 ( .B1(n552), .B2(n557), .A(n553), .ZN(n543) );
  NAND2_X1 U476 ( .A1(n283), .A2(instr_rdata_i[26]), .ZN(n546) );
  NAND2_X1 U477 ( .A1(n284), .A2(n2678), .ZN(n539) );
  OAI21_X1 U478 ( .B1(n538), .B2(n546), .A(n539), .ZN(n285) );
  AOI21_X1 U479 ( .B1(n286), .B2(n543), .A(n285), .ZN(n287) );
  INV_X1 U481 ( .A(regfile_data_ra_id[28]), .ZN(n2069) );
  OAI22_X1 U482 ( .A1(n2672), .A2(n209), .B1(n90), .B2(n2069), .ZN(n336) );
  NOR2_X1 U483 ( .A1(n336), .A2(n352), .ZN(n373) );
  INV_X1 U484 ( .A(pc_id_i[29]), .ZN(n291) );
  INV_X1 U485 ( .A(regfile_data_ra_id[29]), .ZN(n2080) );
  OAI22_X1 U486 ( .A1(n2672), .A2(n291), .B1(n90), .B2(n2080), .ZN(n335) );
  NOR2_X1 U487 ( .A1(n335), .A2(n352), .ZN(n362) );
  NOR2_X1 U488 ( .A1(n373), .A2(n362), .ZN(n581) );
  AOI22_X1 U489 ( .A1(regfile_data_ra_id[30]), .A2(n23), .B1(pc_id_i[30]), 
        .B2(n349), .ZN(n293) );
  INV_X1 U490 ( .A(n293), .ZN(n337) );
  OR2_X1 U491 ( .A1(n337), .A2(n352), .ZN(n593) );
  NAND2_X1 U492 ( .A1(n581), .A2(n593), .ZN(n301) );
  INV_X1 U493 ( .A(regfile_data_ra_id[24]), .ZN(n295) );
  NAND2_X1 U494 ( .A1(n349), .A2(pc_id_i[24]), .ZN(n294) );
  OAI21_X1 U495 ( .B1(n295), .B2(n90), .A(n294), .ZN(n340) );
  NOR2_X1 U496 ( .A1(n340), .A2(n352), .ZN(n398) );
  INV_X1 U497 ( .A(regfile_data_ra_id[25]), .ZN(n297) );
  NAND2_X1 U498 ( .A1(n349), .A2(pc_id_i[25]), .ZN(n296) );
  OAI21_X1 U499 ( .B1(n297), .B2(n90), .A(n296), .ZN(n339) );
  NOR2_X1 U500 ( .A1(n339), .A2(n352), .ZN(n403) );
  NOR2_X1 U501 ( .A1(n398), .A2(n403), .ZN(n390) );
  INV_X1 U502 ( .A(regfile_data_ra_id[26]), .ZN(n2039) );
  NAND2_X1 U503 ( .A1(n349), .A2(pc_id_i[26]), .ZN(n298) );
  OAI21_X1 U504 ( .B1(n2039), .B2(n90), .A(n298), .ZN(n342) );
  NOR2_X1 U505 ( .A1(n342), .A2(n352), .ZN(n393) );
  INV_X1 U506 ( .A(regfile_data_ra_id[27]), .ZN(n2054) );
  NAND2_X1 U507 ( .A1(n349), .A2(pc_id_i[27]), .ZN(n299) );
  OAI21_X1 U508 ( .B1(n2054), .B2(n90), .A(n299), .ZN(n341) );
  NOR2_X1 U509 ( .A1(n341), .A2(n352), .ZN(n384) );
  NOR2_X1 U510 ( .A1(n393), .A2(n384), .ZN(n300) );
  NAND2_X1 U511 ( .A1(n390), .A2(n300), .ZN(n583) );
  NOR2_X1 U512 ( .A1(n301), .A2(n583), .ZN(n346) );
  NAND2_X1 U513 ( .A1(n349), .A2(pc_id_i[20]), .ZN(n302) );
  NOR2_X1 U514 ( .A1(n329), .A2(n352), .ZN(n434) );
  INV_X1 U515 ( .A(n2644), .ZN(n1958) );
  NAND2_X1 U516 ( .A1(n349), .A2(pc_id_i[21]), .ZN(n304) );
  OAI21_X1 U517 ( .B1(n1958), .B2(n90), .A(n304), .ZN(n328) );
  INV_X1 U518 ( .A(regfile_data_ra_id[22]), .ZN(n306) );
  NAND2_X1 U519 ( .A1(n349), .A2(pc_id_i[22]), .ZN(n305) );
  OAI21_X1 U520 ( .B1(n306), .B2(n90), .A(n305), .ZN(n331) );
  NOR2_X1 U521 ( .A1(n331), .A2(n352), .ZN(n429) );
  INV_X1 U522 ( .A(regfile_data_ra_id[23]), .ZN(n308) );
  NAND2_X1 U523 ( .A1(n349), .A2(pc_id_i[23]), .ZN(n307) );
  OAI21_X1 U524 ( .B1(n308), .B2(n90), .A(n307), .ZN(n330) );
  NOR2_X1 U525 ( .A1(n330), .A2(n352), .ZN(n420) );
  NOR2_X1 U526 ( .A1(n429), .A2(n420), .ZN(n309) );
  NAND2_X1 U527 ( .A1(n426), .A2(n309), .ZN(n334) );
  NAND2_X1 U528 ( .A1(n349), .A2(pc_id_i[16]), .ZN(n310) );
  NOR2_X1 U529 ( .A1(n48), .A2(n1008), .ZN(n312) );
  OR2_X1 U530 ( .A1(n312), .A2(n311), .ZN(n319) );
  NAND2_X1 U532 ( .A1(n277), .A2(pc_id_i[17]), .ZN(n313) );
  OAI21_X1 U533 ( .B1(n770), .B2(n48), .A(n317), .ZN(n321) );
  NOR2_X1 U534 ( .A1(n576), .A2(n468), .ZN(n460) );
  INV_X1 U535 ( .A(regfile_data_ra_id[18]), .ZN(n1919) );
  NAND2_X1 U536 ( .A1(n349), .A2(pc_id_i[18]), .ZN(n314) );
  OAI21_X1 U537 ( .B1(n1919), .B2(n90), .A(n314), .ZN(n323) );
  OAI21_X1 U538 ( .B1(n1914), .B2(n48), .A(n2669), .ZN(n322) );
  NOR2_X1 U539 ( .A1(n323), .A2(n322), .ZN(n451) );
  NAND2_X1 U540 ( .A1(n277), .A2(pc_id_i[19]), .ZN(n315) );
  OAI21_X1 U541 ( .B1(n1010), .B2(n48), .A(n2669), .ZN(n324) );
  NOR2_X1 U542 ( .A1(n325), .A2(n324), .ZN(n455) );
  NOR2_X1 U543 ( .A1(n334), .A2(n446), .ZN(n367) );
  NAND2_X1 U544 ( .A1(n346), .A2(n584), .ZN(n348) );
  NAND2_X1 U545 ( .A1(n320), .A2(n319), .ZN(n577) );
  OAI21_X1 U546 ( .B1(n468), .B2(n577), .A(n469), .ZN(n461) );
  NAND2_X1 U547 ( .A1(n323), .A2(n322), .ZN(n464) );
  NAND2_X1 U548 ( .A1(n325), .A2(n324), .ZN(n456) );
  OAI21_X1 U549 ( .B1(n455), .B2(n464), .A(n456), .ZN(n326) );
  AOI21_X1 U550 ( .B1(n327), .B2(n461), .A(n326), .ZN(n445) );
  NAND2_X1 U551 ( .A1(n328), .A2(instr_rdata_i[31]), .ZN(n441) );
  NAND2_X1 U552 ( .A1(n329), .A2(instr_rdata_i[31]), .ZN(n447) );
  NAND2_X1 U553 ( .A1(n441), .A2(n447), .ZN(n425) );
  NAND2_X1 U554 ( .A1(n330), .A2(instr_rdata_i[31]), .ZN(n421) );
  NAND2_X1 U555 ( .A1(n331), .A2(instr_rdata_i[31]), .ZN(n430) );
  NAND2_X1 U556 ( .A1(n421), .A2(n430), .ZN(n332) );
  NOR2_X1 U557 ( .A1(n425), .A2(n332), .ZN(n333) );
  NAND2_X1 U558 ( .A1(n335), .A2(n352), .ZN(n363) );
  NAND2_X1 U559 ( .A1(n336), .A2(n352), .ZN(n374) );
  NAND2_X1 U560 ( .A1(n363), .A2(n374), .ZN(n585) );
  NAND2_X1 U561 ( .A1(n337), .A2(n352), .ZN(n592) );
  INV_X1 U562 ( .A(n592), .ZN(n338) );
  NOR2_X1 U563 ( .A1(n585), .A2(n338), .ZN(n344) );
  NAND2_X1 U564 ( .A1(n339), .A2(n352), .ZN(n404) );
  NAND2_X1 U565 ( .A1(n340), .A2(instr_rdata_i[31]), .ZN(n410) );
  NAND2_X1 U566 ( .A1(n404), .A2(n410), .ZN(n389) );
  NAND2_X1 U567 ( .A1(n341), .A2(n352), .ZN(n385) );
  NAND2_X1 U568 ( .A1(n342), .A2(instr_rdata_i[31]), .ZN(n394) );
  NAND2_X1 U569 ( .A1(n385), .A2(n394), .ZN(n343) );
  NOR2_X1 U570 ( .A1(n389), .A2(n343), .ZN(n586) );
  NAND2_X1 U571 ( .A1(n344), .A2(n586), .ZN(n345) );
  AOI21_X1 U572 ( .B1(n346), .B2(n368), .A(n345), .ZN(n347) );
  OAI21_X1 U573 ( .B1(n580), .B2(n348), .A(n347), .ZN(n357) );
  AOI22_X1 U574 ( .A1(regfile_data_ra_id[31]), .A2(n23), .B1(pc_id_i[31]), 
        .B2(n349), .ZN(n351) );
  INV_X1 U575 ( .A(n351), .ZN(n353) );
  OR2_X1 U576 ( .A1(n353), .A2(n352), .ZN(n355) );
  NAND2_X1 U577 ( .A1(n353), .A2(n352), .ZN(n354) );
  NAND2_X1 U578 ( .A1(n355), .A2(n354), .ZN(n356) );
  XNOR2_X1 U579 ( .A(n357), .B(n356), .ZN(jump_target_o[31]) );
  NOR2_X1 U580 ( .A1(n583), .A2(n373), .ZN(n359) );
  NAND2_X1 U581 ( .A1(n399), .A2(n359), .ZN(n361) );
  NAND2_X1 U582 ( .A1(n374), .A2(n586), .ZN(n358) );
  AOI21_X1 U583 ( .B1(n368), .B2(n359), .A(n358), .ZN(n360) );
  OAI21_X1 U584 ( .B1(n580), .B2(n361), .A(n360), .ZN(n366) );
  INV_X1 U585 ( .A(n362), .ZN(n364) );
  NAND2_X1 U586 ( .A1(n364), .A2(n363), .ZN(n365) );
  XNOR2_X1 U587 ( .A(n366), .B(n365), .ZN(jump_target_o[29]) );
  INV_X1 U588 ( .A(n583), .ZN(n370) );
  NAND2_X1 U589 ( .A1(n399), .A2(n370), .ZN(n372) );
  INV_X1 U590 ( .A(n586), .ZN(n369) );
  AOI21_X1 U591 ( .B1(n368), .B2(n370), .A(n369), .ZN(n371) );
  OAI21_X1 U592 ( .B1(n580), .B2(n372), .A(n371), .ZN(n377) );
  INV_X1 U593 ( .A(n373), .ZN(n375) );
  NAND2_X1 U594 ( .A1(n375), .A2(n374), .ZN(n376) );
  XNOR2_X1 U595 ( .A(n377), .B(n376), .ZN(jump_target_o[28]) );
  INV_X1 U596 ( .A(n390), .ZN(n378) );
  NOR2_X1 U597 ( .A1(n378), .A2(n393), .ZN(n381) );
  NAND2_X1 U598 ( .A1(n399), .A2(n381), .ZN(n383) );
  INV_X1 U599 ( .A(n389), .ZN(n379) );
  NAND2_X1 U600 ( .A1(n394), .A2(n379), .ZN(n380) );
  AOI21_X1 U601 ( .B1(n368), .B2(n381), .A(n380), .ZN(n382) );
  OAI21_X1 U602 ( .B1(n580), .B2(n383), .A(n382), .ZN(n388) );
  INV_X1 U603 ( .A(n384), .ZN(n386) );
  NAND2_X1 U604 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U605 ( .A(n388), .B(n387), .ZN(jump_target_o[27]) );
  NAND2_X1 U606 ( .A1(n584), .A2(n390), .ZN(n392) );
  AOI21_X1 U607 ( .B1(n368), .B2(n390), .A(n389), .ZN(n391) );
  OAI21_X1 U608 ( .B1(n580), .B2(n392), .A(n391), .ZN(n397) );
  INV_X1 U609 ( .A(n393), .ZN(n395) );
  NAND2_X1 U610 ( .A1(n395), .A2(n394), .ZN(n396) );
  XNOR2_X1 U611 ( .A(n397), .B(n396), .ZN(jump_target_o[26]) );
  INV_X1 U612 ( .A(n398), .ZN(n411) );
  NAND2_X1 U613 ( .A1(n399), .A2(n411), .ZN(n402) );
  INV_X1 U614 ( .A(n410), .ZN(n400) );
  AOI21_X1 U615 ( .B1(n368), .B2(n411), .A(n400), .ZN(n401) );
  INV_X1 U616 ( .A(n403), .ZN(n405) );
  NAND2_X1 U617 ( .A1(n405), .A2(n404), .ZN(n406) );
  XNOR2_X1 U618 ( .A(n407), .B(n406), .ZN(jump_target_o[25]) );
  INV_X1 U619 ( .A(n584), .ZN(n409) );
  INV_X1 U620 ( .A(n368), .ZN(n408) );
  OAI21_X1 U621 ( .B1(n580), .B2(n409), .A(n408), .ZN(n413) );
  NAND2_X1 U622 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U623 ( .A(n413), .B(n412), .ZN(jump_target_o[24]) );
  INV_X1 U624 ( .A(n426), .ZN(n414) );
  NOR2_X1 U625 ( .A1(n414), .A2(n429), .ZN(n417) );
  INV_X1 U626 ( .A(n446), .ZN(n435) );
  NAND2_X1 U627 ( .A1(n417), .A2(n435), .ZN(n419) );
  INV_X1 U628 ( .A(n445), .ZN(n437) );
  INV_X1 U629 ( .A(n425), .ZN(n415) );
  NAND2_X1 U630 ( .A1(n430), .A2(n415), .ZN(n416) );
  AOI21_X1 U631 ( .B1(n417), .B2(n437), .A(n416), .ZN(n418) );
  OAI21_X1 U632 ( .B1(n580), .B2(n419), .A(n418), .ZN(n424) );
  INV_X1 U633 ( .A(n420), .ZN(n422) );
  NAND2_X1 U634 ( .A1(n422), .A2(n421), .ZN(n423) );
  XNOR2_X1 U635 ( .A(n424), .B(n423), .ZN(jump_target_o[23]) );
  NAND2_X1 U636 ( .A1(n435), .A2(n426), .ZN(n428) );
  AOI21_X1 U637 ( .B1(n437), .B2(n426), .A(n425), .ZN(n427) );
  OAI21_X1 U638 ( .B1(n580), .B2(n428), .A(n427), .ZN(n433) );
  INV_X1 U639 ( .A(n429), .ZN(n431) );
  NAND2_X1 U640 ( .A1(n431), .A2(n430), .ZN(n432) );
  XNOR2_X1 U641 ( .A(n433), .B(n432), .ZN(jump_target_o[22]) );
  INV_X1 U642 ( .A(n434), .ZN(n448) );
  NAND2_X1 U643 ( .A1(n435), .A2(n448), .ZN(n439) );
  INV_X1 U644 ( .A(n447), .ZN(n436) );
  AOI21_X1 U645 ( .B1(n437), .B2(n448), .A(n436), .ZN(n438) );
  OAI21_X1 U646 ( .B1(n580), .B2(n439), .A(n438), .ZN(n444) );
  INV_X1 U647 ( .A(n440), .ZN(n442) );
  NAND2_X1 U648 ( .A1(n442), .A2(n441), .ZN(n443) );
  XNOR2_X1 U649 ( .A(n444), .B(n443), .ZN(jump_target_o[21]) );
  OAI21_X1 U650 ( .B1(n580), .B2(n446), .A(n445), .ZN(n450) );
  NAND2_X1 U651 ( .A1(n448), .A2(n447), .ZN(n449) );
  XNOR2_X1 U652 ( .A(n450), .B(n449), .ZN(jump_target_o[20]) );
  INV_X1 U653 ( .A(n451), .ZN(n465) );
  NAND2_X1 U654 ( .A1(n460), .A2(n465), .ZN(n454) );
  INV_X1 U655 ( .A(n464), .ZN(n452) );
  AOI21_X1 U656 ( .B1(n461), .B2(n465), .A(n452), .ZN(n453) );
  OAI21_X1 U657 ( .B1(n580), .B2(n454), .A(n453), .ZN(n459) );
  INV_X1 U658 ( .A(n455), .ZN(n457) );
  NAND2_X1 U659 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U660 ( .A(n459), .B(n458), .ZN(jump_target_o[19]) );
  INV_X1 U661 ( .A(n460), .ZN(n463) );
  INV_X1 U662 ( .A(n461), .ZN(n462) );
  OAI21_X1 U663 ( .B1(n580), .B2(n463), .A(n462), .ZN(n467) );
  NAND2_X1 U664 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U665 ( .A(n467), .B(n466), .ZN(jump_target_o[18]) );
  NAND2_X1 U667 ( .A1(n2670), .A2(n469), .ZN(n471) );
  XNOR2_X1 U668 ( .A(n472), .B(n471), .ZN(jump_target_o[17]) );
  INV_X1 U669 ( .A(n473), .ZN(n600) );
  INV_X1 U670 ( .A(n487), .ZN(n474) );
  NOR2_X1 U671 ( .A1(n474), .A2(n490), .ZN(n478) );
  INV_X1 U672 ( .A(n506), .ZN(n496) );
  NAND2_X1 U673 ( .A1(n478), .A2(n496), .ZN(n480) );
  INV_X1 U674 ( .A(n475), .ZN(n498) );
  INV_X1 U675 ( .A(n486), .ZN(n476) );
  OAI21_X1 U676 ( .B1(n476), .B2(n490), .A(n491), .ZN(n477) );
  AOI21_X1 U677 ( .B1(n478), .B2(n498), .A(n477), .ZN(n479) );
  OAI21_X1 U678 ( .B1(n600), .B2(n480), .A(n479), .ZN(n485) );
  INV_X1 U679 ( .A(n481), .ZN(n483) );
  NAND2_X1 U680 ( .A1(n483), .A2(n482), .ZN(n484) );
  XNOR2_X1 U681 ( .A(n485), .B(n484), .ZN(jump_target_o[15]) );
  NAND2_X1 U682 ( .A1(n496), .A2(n487), .ZN(n489) );
  AOI21_X1 U683 ( .B1(n498), .B2(n487), .A(n486), .ZN(n488) );
  OAI21_X1 U684 ( .B1(n600), .B2(n489), .A(n488), .ZN(n494) );
  INV_X1 U685 ( .A(n490), .ZN(n492) );
  NAND2_X1 U686 ( .A1(n492), .A2(n491), .ZN(n493) );
  XNOR2_X1 U687 ( .A(n494), .B(n493), .ZN(jump_target_o[14]) );
  INV_X1 U688 ( .A(n495), .ZN(n508) );
  NAND2_X1 U689 ( .A1(n496), .A2(n508), .ZN(n500) );
  INV_X1 U690 ( .A(n507), .ZN(n497) );
  AOI21_X1 U691 ( .B1(n498), .B2(n508), .A(n497), .ZN(n499) );
  OAI21_X1 U692 ( .B1(n600), .B2(n500), .A(n499), .ZN(n505) );
  INV_X1 U693 ( .A(n501), .ZN(n503) );
  NAND2_X1 U694 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U695 ( .A(n505), .B(n504), .ZN(jump_target_o[13]) );
  OAI21_X1 U696 ( .B1(n600), .B2(n506), .A(n475), .ZN(n510) );
  NAND2_X1 U697 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U698 ( .A(n510), .B(n509), .ZN(jump_target_o[12]) );
  INV_X1 U699 ( .A(n511), .ZN(n525) );
  NAND2_X1 U700 ( .A1(n520), .A2(n525), .ZN(n514) );
  INV_X1 U701 ( .A(n524), .ZN(n512) );
  AOI21_X1 U702 ( .B1(n521), .B2(n525), .A(n512), .ZN(n513) );
  OAI21_X1 U703 ( .B1(n600), .B2(n514), .A(n513), .ZN(n519) );
  INV_X1 U704 ( .A(n515), .ZN(n517) );
  NAND2_X1 U705 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U706 ( .A(n519), .B(n518), .ZN(jump_target_o[11]) );
  INV_X1 U707 ( .A(n520), .ZN(n523) );
  INV_X1 U708 ( .A(n521), .ZN(n522) );
  OAI21_X1 U709 ( .B1(n600), .B2(n523), .A(n522), .ZN(n527) );
  NAND2_X1 U710 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U711 ( .A(n527), .B(n526), .ZN(jump_target_o[10]) );
  OAI21_X1 U712 ( .B1(n600), .B2(n596), .A(n597), .ZN(n532) );
  INV_X1 U713 ( .A(n528), .ZN(n530) );
  NAND2_X1 U714 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U715 ( .A(n532), .B(n531), .ZN(jump_target_o[9]) );
  INV_X1 U716 ( .A(n544), .ZN(n533) );
  NOR2_X1 U717 ( .A1(n533), .A2(n545), .ZN(n537) );
  INV_X1 U718 ( .A(n534), .ZN(n560) );
  INV_X1 U719 ( .A(n543), .ZN(n535) );
  OAI21_X1 U720 ( .B1(n535), .B2(n545), .A(n546), .ZN(n536) );
  AOI21_X1 U721 ( .B1(n537), .B2(n560), .A(n536), .ZN(n542) );
  INV_X1 U722 ( .A(n538), .ZN(n540) );
  NAND2_X1 U723 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U724 ( .A(n542), .B(n541), .Z(jump_target_o[7]) );
  AOI21_X1 U725 ( .B1(n560), .B2(n544), .A(n543), .ZN(n549) );
  INV_X1 U726 ( .A(n545), .ZN(n547) );
  NAND2_X1 U727 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U728 ( .A(n549), .B(n548), .Z(jump_target_o[6]) );
  INV_X1 U729 ( .A(n550), .ZN(n558) );
  INV_X1 U730 ( .A(n557), .ZN(n551) );
  AOI21_X1 U731 ( .B1(n560), .B2(n558), .A(n551), .ZN(n556) );
  INV_X1 U732 ( .A(n552), .ZN(n554) );
  NAND2_X1 U733 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U734 ( .A(n556), .B(n555), .Z(jump_target_o[5]) );
  NAND2_X1 U735 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U736 ( .A(n560), .B(n559), .ZN(jump_target_o[4]) );
  INV_X1 U737 ( .A(n561), .ZN(n571) );
  OAI21_X1 U738 ( .B1(n571), .B2(n567), .A(n568), .ZN(n566) );
  INV_X1 U739 ( .A(n562), .ZN(n564) );
  NAND2_X1 U740 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U741 ( .A(n566), .B(n565), .ZN(jump_target_o[3]) );
  INV_X1 U742 ( .A(n567), .ZN(n569) );
  NAND2_X1 U743 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U744 ( .A(n571), .B(n570), .Z(jump_target_o[2]) );
  INV_X1 U745 ( .A(n572), .ZN(n574) );
  NAND2_X1 U746 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U747 ( .A(n1042), .B(n575), .Z(jump_target_o[1]) );
  INV_X1 U748 ( .A(n576), .ZN(n578) );
  NAND2_X1 U749 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U750 ( .A(n580), .B(n579), .Z(jump_target_o[16]) );
  INV_X1 U751 ( .A(n581), .ZN(n582) );
  NOR2_X1 U752 ( .A1(n583), .A2(n582), .ZN(n589) );
  NAND2_X1 U753 ( .A1(n584), .A2(n589), .ZN(n591) );
  INV_X1 U754 ( .A(n585), .ZN(n587) );
  NAND2_X1 U755 ( .A1(n587), .A2(n586), .ZN(n588) );
  AOI21_X1 U756 ( .B1(n368), .B2(n589), .A(n588), .ZN(n590) );
  OAI21_X1 U757 ( .B1(n580), .B2(n591), .A(n590), .ZN(n595) );
  NAND2_X1 U758 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U759 ( .A(n595), .B(n594), .ZN(jump_target_o[30]) );
  INV_X1 U760 ( .A(n596), .ZN(n598) );
  NAND2_X1 U761 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U762 ( .A(n600), .B(n599), .Z(jump_target_o[8]) );
  AOI21_X1 U764 ( .B1(n2574), .B2(csr_hwlp_we_i[0]), .A(n1005), .ZN(n601) );
  INV_X1 U765 ( .A(n601), .ZN(hwloop_we[0]) );
  INV_X1 U766 ( .A(operand_b_fw_mux_sel[0]), .ZN(n602) );
  OR2_X1 U767 ( .A1(n602), .A2(operand_b_fw_mux_sel[1]), .ZN(n1882) );
  INV_X1 U768 ( .A(n1882), .ZN(n2205) );
  INV_X1 U769 ( .A(n2207), .ZN(n1764) );
  AOI22_X1 U770 ( .A1(regfile_wdata_wb_i[6]), .A2(n2207), .B1(n2209), .B2(
        regfile_data_rb_id[6]), .ZN(n603) );
  INV_X1 U771 ( .A(n603), .ZN(n604) );
  NAND2_X1 U776 ( .A1(hwloop_we_int[2]), .A2(hwloop_cnt_mux_sel), .ZN(n719) );
  INV_X1 U777 ( .A(operand_a_fw_mux_sel[0]), .ZN(n607) );
  NOR2_X2 U778 ( .A1(n607), .A2(operand_a_fw_mux_sel[1]), .ZN(n1879) );
  INV_X1 U779 ( .A(n1879), .ZN(n2177) );
  NOR2_X1 U780 ( .A1(n719), .A2(n2177), .ZN(n811) );
  AND2_X1 U781 ( .A1(n607), .A2(operand_a_fw_mux_sel[1]), .ZN(n2179) );
  INV_X1 U782 ( .A(n2179), .ZN(n1884) );
  INV_X1 U783 ( .A(regfile_wdata_wb_i[0]), .ZN(n1202) );
  AND2_X1 U784 ( .A1(n2177), .A2(n1884), .ZN(n1649) );
  INV_X1 U785 ( .A(n1649), .ZN(n2130) );
  NAND2_X1 U786 ( .A1(n53), .A2(n114), .ZN(n610) );
  INV_X1 U787 ( .A(hwloop_cnt_mux_sel), .ZN(n608) );
  AND2_X1 U788 ( .A1(hwloop_we_int[2]), .A2(n608), .ZN(n784) );
  AOI22_X1 U789 ( .A1(n784), .A2(instr_rdata_i[20]), .B1(n615), .B2(
        csr_hwlp_data_i[0]), .ZN(n609) );
  OAI211_X1 U790 ( .C1(n814), .C2(n1202), .A(n610), .B(n609), .ZN(n611) );
  AOI21_X1 U791 ( .B1(regfile_alu_wdata_fw_i[0]), .B2(n788), .A(n611), .ZN(
        n612) );
  INV_X1 U792 ( .A(n612), .ZN(hwloop_cnt[0]) );
  INV_X1 U793 ( .A(n814), .ZN(n616) );
  INV_X1 U794 ( .A(regfile_wdata_wb_i[31]), .ZN(n2420) );
  NAND2_X1 U795 ( .A1(regfile_alu_wdata_fw_i[31]), .A2(n811), .ZN(n614) );
  AOI22_X1 U796 ( .A1(n53), .A2(regfile_data_ra_id[31]), .B1(
        csr_hwlp_data_i[31]), .B2(n615), .ZN(n613) );
  OAI211_X1 U797 ( .C1(n814), .C2(n2420), .A(n614), .B(n613), .ZN(
        hwloop_cnt[31]) );
  NAND2_X1 U798 ( .A1(regfile_alu_wdata_fw_i[6]), .A2(n788), .ZN(n620) );
  AOI22_X1 U799 ( .A1(n784), .A2(n2683), .B1(n615), .B2(csr_hwlp_data_i[6]), 
        .ZN(n619) );
  NAND2_X1 U800 ( .A1(n53), .A2(n32), .ZN(n618) );
  NAND2_X1 U801 ( .A1(n616), .A2(regfile_wdata_wb_i[6]), .ZN(n617) );
  NAND4_X1 U802 ( .A1(n620), .A2(n619), .A3(n618), .A4(n617), .ZN(
        hwloop_cnt[6]) );
  INV_X1 U803 ( .A(regfile_wdata_wb_i[27]), .ZN(n2378) );
  NAND2_X1 U804 ( .A1(regfile_alu_wdata_fw_i[27]), .A2(n788), .ZN(n622) );
  AOI22_X1 U805 ( .A1(n53), .A2(regfile_data_ra_id[27]), .B1(
        csr_hwlp_data_i[27]), .B2(n615), .ZN(n621) );
  OAI211_X1 U806 ( .C1(n814), .C2(n2378), .A(n622), .B(n621), .ZN(
        hwloop_cnt[27]) );
  INV_X1 U807 ( .A(regfile_wdata_wb_i[30]), .ZN(n2406) );
  NAND2_X1 U808 ( .A1(regfile_alu_wdata_fw_i[30]), .A2(n788), .ZN(n624) );
  AOI22_X1 U809 ( .A1(n53), .A2(regfile_data_ra_id[30]), .B1(
        csr_hwlp_data_i[30]), .B2(n615), .ZN(n623) );
  OAI211_X1 U810 ( .C1(n814), .C2(n2406), .A(n624), .B(n623), .ZN(
        hwloop_cnt[30]) );
  INV_X1 U811 ( .A(regfile_wdata_wb_i[25]), .ZN(n2360) );
  AOI22_X1 U813 ( .A1(n53), .A2(regfile_data_ra_id[25]), .B1(
        csr_hwlp_data_i[25]), .B2(n615), .ZN(n625) );
  NAND2_X1 U815 ( .A1(regfile_wdata_wb_i[3]), .A2(n2179), .ZN(n628) );
  NAND2_X1 U816 ( .A1(n1649), .A2(regfile_data_ra_id[3]), .ZN(n627) );
  NAND2_X1 U817 ( .A1(n628), .A2(n627), .ZN(n629) );
  AOI21_X1 U818 ( .B1(regfile_alu_wdata_fw_i[3]), .B2(n1879), .A(n629), .ZN(
        n1664) );
  AOI22_X1 U819 ( .A1(n784), .A2(instr_rdata_i[23]), .B1(n615), .B2(
        csr_hwlp_data_i[3]), .ZN(n630) );
  OAI21_X1 U820 ( .B1(n1664), .B2(n719), .A(n630), .ZN(hwloop_cnt[3]) );
  AOI22_X1 U821 ( .A1(regfile_wdata_wb_i[8]), .A2(n2207), .B1(n2209), .B2(
        regfile_data_rb_id[8]), .ZN(n631) );
  INV_X1 U822 ( .A(n631), .ZN(n632) );
  NAND2_X1 U825 ( .A1(regfile_wdata_wb_i[9]), .A2(n2207), .ZN(n635) );
  NAND2_X1 U826 ( .A1(n2209), .A2(regfile_data_rb_id[9]), .ZN(n634) );
  NAND2_X1 U827 ( .A1(n635), .A2(n634), .ZN(n636) );
  INV_X1 U831 ( .A(bmask_b_mux[1]), .ZN(n2462) );
  NAND2_X1 U834 ( .A1(regfile_wdata_wb_i[3]), .A2(n2207), .ZN(n641) );
  NAND2_X1 U835 ( .A1(n2209), .A2(regfile_data_rb_id[3]), .ZN(n640) );
  NAND2_X1 U836 ( .A1(n641), .A2(n640), .ZN(n642) );
  AOI21_X1 U837 ( .B1(regfile_alu_wdata_fw_i[3]), .B2(n2205), .A(n642), .ZN(
        n2161) );
  INV_X1 U838 ( .A(n2161), .ZN(n643) );
  INV_X1 U845 ( .A(regfile_wdata_wb_i[28]), .ZN(n2387) );
  AOI22_X1 U847 ( .A1(n53), .A2(regfile_data_ra_id[28]), .B1(
        csr_hwlp_data_i[28]), .B2(n615), .ZN(n646) );
  INV_X1 U849 ( .A(regfile_wdata_wb_i[2]), .ZN(n1053) );
  NAND2_X1 U850 ( .A1(n53), .A2(n2627), .ZN(n649) );
  AOI22_X1 U851 ( .A1(n784), .A2(instr_rdata_i[22]), .B1(n615), .B2(
        csr_hwlp_data_i[2]), .ZN(n648) );
  OAI211_X1 U852 ( .C1(n814), .C2(n1053), .A(n649), .B(n648), .ZN(n650) );
  AOI21_X1 U853 ( .B1(regfile_alu_wdata_fw_i[2]), .B2(n788), .A(n650), .ZN(
        n651) );
  INV_X1 U854 ( .A(n651), .ZN(hwloop_cnt[2]) );
  INV_X1 U855 ( .A(regfile_wdata_wb_i[11]), .ZN(n1781) );
  NAND2_X1 U856 ( .A1(n53), .A2(n25), .ZN(n653) );
  AOI22_X1 U857 ( .A1(n784), .A2(instr_rdata_i[31]), .B1(n615), .B2(
        csr_hwlp_data_i[11]), .ZN(n652) );
  OAI211_X1 U858 ( .C1(n814), .C2(n1781), .A(n653), .B(n652), .ZN(n654) );
  AOI21_X1 U859 ( .B1(regfile_alu_wdata_fw_i[11]), .B2(n788), .A(n654), .ZN(
        n655) );
  INV_X1 U860 ( .A(n655), .ZN(hwloop_cnt[11]) );
  NAND2_X1 U861 ( .A1(regfile_alu_wdata_fw_i[5]), .A2(n2205), .ZN(n657) );
  AOI22_X1 U862 ( .A1(regfile_wdata_wb_i[5]), .A2(n2207), .B1(n2209), .B2(
        regfile_data_rb_id[5]), .ZN(n656) );
  NAND2_X1 U863 ( .A1(n657), .A2(n656), .ZN(n1692) );
  INV_X1 U864 ( .A(n2660), .ZN(n659) );
  INV_X1 U867 ( .A(regfile_wdata_wb_i[8]), .ZN(n2195) );
  NAND2_X1 U868 ( .A1(n53), .A2(n24), .ZN(n661) );
  AOI22_X1 U869 ( .A1(n784), .A2(n2668), .B1(n615), .B2(csr_hwlp_data_i[8]), 
        .ZN(n660) );
  OAI211_X1 U870 ( .C1(n814), .C2(n2195), .A(n661), .B(n660), .ZN(n662) );
  AOI21_X1 U871 ( .B1(regfile_alu_wdata_fw_i[8]), .B2(n788), .A(n662), .ZN(
        n663) );
  INV_X1 U872 ( .A(n663), .ZN(hwloop_cnt[8]) );
  INV_X1 U873 ( .A(regfile_wdata_wb_i[29]), .ZN(n2396) );
  NAND2_X1 U874 ( .A1(regfile_alu_wdata_fw_i[29]), .A2(n788), .ZN(n665) );
  AOI22_X1 U875 ( .A1(n53), .A2(regfile_data_ra_id[29]), .B1(
        csr_hwlp_data_i[29]), .B2(n615), .ZN(n664) );
  OAI211_X1 U876 ( .C1(n814), .C2(n2396), .A(n665), .B(n664), .ZN(
        hwloop_cnt[29]) );
  INV_X1 U877 ( .A(regfile_wdata_wb_i[9]), .ZN(n2201) );
  NAND2_X1 U878 ( .A1(n53), .A2(regfile_data_ra_id[9]), .ZN(n667) );
  AOI22_X1 U879 ( .A1(n784), .A2(instr_rdata_i[29]), .B1(n615), .B2(
        csr_hwlp_data_i[9]), .ZN(n666) );
  OAI211_X1 U880 ( .C1(n814), .C2(n2201), .A(n667), .B(n666), .ZN(n668) );
  AOI21_X1 U881 ( .B1(regfile_alu_wdata_fw_i[9]), .B2(n788), .A(n668), .ZN(
        n669) );
  INV_X1 U882 ( .A(n669), .ZN(hwloop_cnt[9]) );
  INV_X1 U883 ( .A(regfile_wdata_wb_i[26]), .ZN(n2369) );
  NAND2_X1 U884 ( .A1(regfile_alu_wdata_fw_i[26]), .A2(n788), .ZN(n671) );
  AOI22_X1 U885 ( .A1(n53), .A2(regfile_data_ra_id[26]), .B1(
        csr_hwlp_data_i[26]), .B2(n615), .ZN(n670) );
  OAI211_X1 U886 ( .C1(n814), .C2(n2369), .A(n671), .B(n670), .ZN(
        hwloop_cnt[26]) );
  NAND2_X1 U887 ( .A1(regfile_alu_wdata_fw_i[12]), .A2(n788), .ZN(n673) );
  AOI22_X1 U888 ( .A1(n616), .A2(regfile_wdata_wb_i[12]), .B1(
        csr_hwlp_data_i[12]), .B2(n615), .ZN(n672) );
  OAI211_X1 U889 ( .C1(n94), .C2(n1806), .A(n673), .B(n672), .ZN(
        hwloop_cnt[12]) );
  NAND2_X1 U890 ( .A1(regfile_alu_wdata_fw_i[14]), .A2(n788), .ZN(n675) );
  AOI22_X1 U891 ( .A1(n616), .A2(regfile_wdata_wb_i[14]), .B1(
        csr_hwlp_data_i[14]), .B2(n615), .ZN(n674) );
  OAI211_X1 U892 ( .C1(n94), .C2(n1828), .A(n675), .B(n674), .ZN(
        hwloop_cnt[14]) );
  INV_X1 U893 ( .A(regfile_wdata_wb_i[20]), .ZN(n2315) );
  NAND2_X1 U894 ( .A1(regfile_alu_wdata_fw_i[20]), .A2(n811), .ZN(n677) );
  AOI22_X1 U895 ( .A1(n53), .A2(regfile_data_ra_id[20]), .B1(
        csr_hwlp_data_i[20]), .B2(n615), .ZN(n676) );
  OAI211_X1 U896 ( .C1(n814), .C2(n2315), .A(n677), .B(n676), .ZN(
        hwloop_cnt[20]) );
  NAND2_X1 U897 ( .A1(regfile_alu_wdata_fw_i[1]), .A2(n2205), .ZN(n679) );
  AOI22_X1 U898 ( .A1(regfile_wdata_wb_i[1]), .A2(n2207), .B1(n2209), .B2(
        regfile_data_rb_id[1]), .ZN(n678) );
  NAND2_X1 U899 ( .A1(n679), .A2(n678), .ZN(n1229) );
  NAND2_X1 U903 ( .A1(n2663), .A2(n811), .ZN(n683) );
  AOI22_X1 U904 ( .A1(n616), .A2(regfile_wdata_wb_i[15]), .B1(
        csr_hwlp_data_i[15]), .B2(n615), .ZN(n682) );
  OAI211_X1 U905 ( .C1(n94), .C2(n1840), .A(n683), .B(n682), .ZN(
        hwloop_cnt[15]) );
  NAND2_X1 U906 ( .A1(regfile_alu_wdata_fw_i[13]), .A2(n811), .ZN(n685) );
  AOI22_X1 U907 ( .A1(n616), .A2(regfile_wdata_wb_i[13]), .B1(
        csr_hwlp_data_i[13]), .B2(n615), .ZN(n684) );
  INV_X1 U908 ( .A(regfile_wdata_wb_i[23]), .ZN(n2342) );
  NAND2_X1 U909 ( .A1(regfile_alu_wdata_fw_i[23]), .A2(n811), .ZN(n687) );
  INV_X1 U910 ( .A(csr_hwlp_data_i[23]), .ZN(n974) );
  AOI22_X1 U911 ( .A1(n53), .A2(regfile_data_ra_id[23]), .B1(
        csr_hwlp_data_i[23]), .B2(n615), .ZN(n686) );
  OAI211_X1 U912 ( .C1(n814), .C2(n2342), .A(n687), .B(n686), .ZN(
        hwloop_cnt[23]) );
  INV_X1 U913 ( .A(regfile_wdata_wb_i[17]), .ZN(n2285) );
  NAND2_X1 U914 ( .A1(regfile_alu_wdata_fw_i[17]), .A2(n811), .ZN(n689) );
  AOI22_X1 U915 ( .A1(n53), .A2(regfile_data_ra_id[17]), .B1(
        csr_hwlp_data_i[17]), .B2(n615), .ZN(n688) );
  OAI211_X1 U916 ( .C1(n814), .C2(n2285), .A(n689), .B(n688), .ZN(
        hwloop_cnt[17]) );
  INV_X1 U917 ( .A(regfile_wdata_wb_i[19]), .ZN(n2306) );
  NAND2_X1 U918 ( .A1(regfile_alu_wdata_fw_i[19]), .A2(n811), .ZN(n691) );
  AOI22_X1 U919 ( .A1(n53), .A2(regfile_data_ra_id[19]), .B1(
        csr_hwlp_data_i[19]), .B2(n615), .ZN(n690) );
  OAI211_X1 U920 ( .C1(n814), .C2(n2306), .A(n691), .B(n690), .ZN(
        hwloop_cnt[19]) );
  NAND2_X1 U921 ( .A1(regfile_wdata_wb_i[4]), .A2(n2179), .ZN(n693) );
  NAND2_X1 U922 ( .A1(n1649), .A2(regfile_data_ra_id[4]), .ZN(n692) );
  NAND2_X1 U923 ( .A1(n693), .A2(n692), .ZN(n694) );
  AOI21_X1 U924 ( .B1(regfile_alu_wdata_fw_i[4]), .B2(n1879), .A(n694), .ZN(
        n1681) );
  AOI22_X1 U925 ( .A1(n784), .A2(n2604), .B1(n615), .B2(csr_hwlp_data_i[4]), 
        .ZN(n695) );
  OAI21_X1 U926 ( .B1(n1681), .B2(n719), .A(n695), .ZN(hwloop_cnt[4]) );
  INV_X1 U927 ( .A(regfile_wdata_wb_i[22]), .ZN(n2333) );
  NAND2_X1 U928 ( .A1(regfile_alu_wdata_fw_i[22]), .A2(n811), .ZN(n697) );
  AOI22_X1 U929 ( .A1(n53), .A2(regfile_data_ra_id[22]), .B1(
        csr_hwlp_data_i[22]), .B2(n615), .ZN(n696) );
  OAI211_X1 U930 ( .C1(n814), .C2(n2333), .A(n697), .B(n696), .ZN(
        hwloop_cnt[22]) );
  NAND2_X1 U931 ( .A1(regfile_wdata_wb_i[4]), .A2(n2207), .ZN(n699) );
  NAND2_X1 U932 ( .A1(n2209), .A2(regfile_data_rb_id[4]), .ZN(n698) );
  NAND2_X1 U933 ( .A1(n699), .A2(n698), .ZN(n700) );
  AOI21_X1 U934 ( .B1(regfile_alu_wdata_fw_i[4]), .B2(n2205), .A(n700), .ZN(
        n1685) );
  INV_X1 U935 ( .A(n1685), .ZN(n701) );
  INV_X1 U939 ( .A(regfile_wdata_wb_i[18]), .ZN(n2294) );
  NAND2_X1 U940 ( .A1(regfile_alu_wdata_fw_i[18]), .A2(n811), .ZN(n705) );
  AOI22_X1 U941 ( .A1(n53), .A2(regfile_data_ra_id[18]), .B1(
        csr_hwlp_data_i[18]), .B2(n615), .ZN(n704) );
  OAI211_X1 U942 ( .C1(n814), .C2(n2294), .A(n705), .B(n704), .ZN(
        hwloop_cnt[18]) );
  INV_X1 U943 ( .A(regfile_wdata_wb_i[24]), .ZN(n2351) );
  NAND2_X1 U944 ( .A1(regfile_alu_wdata_fw_i[24]), .A2(n788), .ZN(n707) );
  AOI22_X1 U945 ( .A1(n53), .A2(regfile_data_ra_id[24]), .B1(
        csr_hwlp_data_i[24]), .B2(n615), .ZN(n706) );
  OAI211_X1 U946 ( .C1(n814), .C2(n2351), .A(n707), .B(n706), .ZN(
        hwloop_cnt[24]) );
  INV_X1 U947 ( .A(regfile_wdata_wb_i[21]), .ZN(n2324) );
  NAND2_X1 U948 ( .A1(regfile_alu_wdata_fw_i[21]), .A2(n788), .ZN(n709) );
  AOI22_X1 U949 ( .A1(n53), .A2(n2644), .B1(csr_hwlp_data_i[21]), .B2(n615), 
        .ZN(n708) );
  OAI211_X1 U950 ( .C1(n814), .C2(n2324), .A(n709), .B(n708), .ZN(
        hwloop_cnt[21]) );
  NAND2_X1 U951 ( .A1(regfile_wdata_wb_i[2]), .A2(n2207), .ZN(n711) );
  NAND2_X1 U952 ( .A1(n2209), .A2(regfile_data_rb_id[2]), .ZN(n710) );
  NAND2_X1 U953 ( .A1(n711), .A2(n710), .ZN(n712) );
  AOI21_X1 U954 ( .B1(regfile_alu_wdata_fw_i[2]), .B2(n2205), .A(n712), .ZN(
        n2148) );
  INV_X1 U955 ( .A(n2148), .ZN(n713) );
  NAND2_X1 U959 ( .A1(regfile_alu_wdata_fw_i[5]), .A2(n1879), .ZN(n718) );
  AOI22_X1 U960 ( .A1(regfile_wdata_wb_i[5]), .A2(n2179), .B1(n1649), .B2(
        regfile_data_ra_id[5]), .ZN(n717) );
  NAND2_X1 U961 ( .A1(n718), .A2(n717), .ZN(n1688) );
  INV_X1 U962 ( .A(n719), .ZN(n725) );
  NAND2_X1 U963 ( .A1(n1688), .A2(n725), .ZN(n721) );
  AOI22_X1 U964 ( .A1(n784), .A2(instr_rdata_i[25]), .B1(n615), .B2(
        csr_hwlp_data_i[5]), .ZN(n720) );
  NAND2_X1 U965 ( .A1(n721), .A2(n720), .ZN(hwloop_cnt[5]) );
  INV_X1 U966 ( .A(n185), .ZN(n722) );
  NAND3_X1 U967 ( .A1(n2577), .A2(n55), .A3(n722), .ZN(clear_instr_valid_o) );
  AND3_X1 U968 ( .A1(clear_instr_valid_o), .A2(instr_valid_i), .A3(is_hwlp_i), 
        .ZN(hwloop_valid) );
  NAND2_X1 U969 ( .A1(regfile_alu_wdata_fw_i[1]), .A2(n1879), .ZN(n724) );
  AOI22_X1 U970 ( .A1(regfile_wdata_wb_i[1]), .A2(n2179), .B1(n1649), .B2(
        regfile_data_ra_id[1]), .ZN(n723) );
  NAND2_X1 U971 ( .A1(n724), .A2(n723), .ZN(n1230) );
  NAND2_X1 U972 ( .A1(n2658), .A2(n725), .ZN(n727) );
  AOI22_X1 U973 ( .A1(n784), .A2(instr_rdata_i[21]), .B1(n615), .B2(
        csr_hwlp_data_i[1]), .ZN(n726) );
  NAND2_X1 U974 ( .A1(n727), .A2(n726), .ZN(hwloop_cnt[1]) );
  INV_X1 U975 ( .A(regc_mux[0]), .ZN(n728) );
  NOR2_X1 U976 ( .A1(regc_mux[1]), .A2(n728), .ZN(n739) );
  NAND2_X1 U977 ( .A1(n739), .A2(instr_rdata_i[9]), .ZN(n730) );
  AND2_X1 U978 ( .A1(regc_mux[1]), .A2(n728), .ZN(n740) );
  NAND2_X1 U979 ( .A1(n740), .A2(n110), .ZN(n729) );
  NAND2_X1 U980 ( .A1(n739), .A2(instr_rdata_i[8]), .ZN(n732) );
  NAND2_X1 U981 ( .A1(n740), .A2(n80), .ZN(n731) );
  NAND2_X1 U982 ( .A1(n739), .A2(instr_rdata_i[10]), .ZN(n734) );
  NAND2_X1 U983 ( .A1(n740), .A2(n33), .ZN(n733) );
  NAND2_X1 U984 ( .A1(n739), .A2(instr_rdata_i[11]), .ZN(n737) );
  NAND2_X1 U985 ( .A1(n740), .A2(n116), .ZN(n736) );
  OAI211_X1 U986 ( .C1(n743), .C2(n738), .A(n737), .B(n736), .ZN(n1638) );
  NAND2_X1 U987 ( .A1(n739), .A2(instr_rdata_i[7]), .ZN(n742) );
  NAND2_X1 U988 ( .A1(n740), .A2(n113), .ZN(n741) );
  OAI211_X1 U989 ( .C1(n743), .C2(n2429), .A(n742), .B(n741), .ZN(n1634) );
  NOR3_X1 U990 ( .A1(n1636), .A2(n1635), .A3(n1637), .ZN(n746) );
  INV_X1 U991 ( .A(n1638), .ZN(n745) );
  INV_X1 U992 ( .A(n1634), .ZN(n744) );
  NAND3_X1 U993 ( .A1(n746), .A2(n745), .A3(n744), .ZN(n747) );
  NAND2_X1 U994 ( .A1(n747), .A2(regc_used_dec), .ZN(n1023) );
  XNOR2_X1 U995 ( .A(n1636), .B(regfile_alu_waddr_ex_o[2]), .ZN(n750) );
  XNOR2_X1 U996 ( .A(n1638), .B(regfile_alu_waddr_ex_o[4]), .ZN(n749) );
  XNOR2_X1 U997 ( .A(n1635), .B(regfile_alu_waddr_ex_o[1]), .ZN(n748) );
  NAND3_X1 U998 ( .A1(n750), .A2(n749), .A3(n748), .ZN(n753) );
  XOR2_X1 U999 ( .A(regfile_alu_waddr_ex_o[0]), .B(n1634), .Z(n752) );
  XOR2_X1 U1000 ( .A(regfile_alu_waddr_ex_o[3]), .B(n1637), .Z(n751) );
  NOR4_X1 U1001 ( .A1(n1023), .A2(n753), .A3(n752), .A4(n751), .ZN(
        reg_d_alu_is_reg_c_id) );
  XNOR2_X1 U1002 ( .A(n1637), .B(regfile_waddr_ex_o[3]), .ZN(n756) );
  XNOR2_X1 U1003 ( .A(n1636), .B(regfile_waddr_ex_o[2]), .ZN(n755) );
  XNOR2_X1 U1004 ( .A(n1635), .B(regfile_waddr_ex_o[1]), .ZN(n754) );
  NAND3_X1 U1005 ( .A1(n756), .A2(n755), .A3(n754), .ZN(n759) );
  XOR2_X1 U1006 ( .A(regfile_waddr_ex_o[0]), .B(n1634), .Z(n758) );
  XOR2_X1 U1007 ( .A(regfile_waddr_ex_o[4]), .B(n1638), .Z(n757) );
  NOR4_X1 U1008 ( .A1(n1023), .A2(n759), .A3(n758), .A4(n757), .ZN(
        reg_d_ex_is_reg_c_id) );
  OR2_X1 U1009 ( .A1(n2604), .A2(instr_rdata_i[23]), .ZN(n1723) );
  NOR2_X1 U1010 ( .A1(n1723), .A2(instr_rdata_i[22]), .ZN(n1656) );
  NOR2_X1 U1011 ( .A1(instr_rdata_i[21]), .A2(instr_rdata_i[20]), .ZN(n1655)
         );
  AND2_X1 U1012 ( .A1(n1656), .A2(n1655), .ZN(n1207) );
  INV_X1 U1013 ( .A(n1207), .ZN(n760) );
  NAND2_X1 U1014 ( .A1(regb_used_dec), .A2(n760), .ZN(n1030) );
  XOR2_X1 U1015 ( .A(regfile_waddr_ex_o[4]), .B(n2604), .Z(n766) );
  XOR2_X1 U1016 ( .A(regfile_waddr_ex_o[3]), .B(instr_rdata_i[23]), .Z(n765)
         );
  XNOR2_X1 U1017 ( .A(instr_rdata_i[22]), .B(regfile_waddr_ex_o[2]), .ZN(n763)
         );
  XNOR2_X1 U1018 ( .A(instr_rdata_i[20]), .B(regfile_waddr_ex_o[0]), .ZN(n762)
         );
  XNOR2_X1 U1019 ( .A(instr_rdata_i[21]), .B(regfile_waddr_ex_o[1]), .ZN(n761)
         );
  NAND3_X1 U1020 ( .A1(n763), .A2(n762), .A3(n761), .ZN(n764) );
  NOR4_X1 U1021 ( .A1(n1030), .A2(n766), .A3(n765), .A4(n764), .ZN(
        reg_d_ex_is_reg_b_id) );
  NAND2_X1 U1022 ( .A1(regfile_alu_waddr_mux_sel), .A2(instr_rdata_i[7]), .ZN(
        n767) );
  OAI21_X1 U1023 ( .B1(regfile_alu_waddr_mux_sel), .B2(n768), .A(n767), .ZN(
        regfile_alu_waddr_id[0]) );
  NAND2_X1 U1024 ( .A1(regfile_alu_waddr_mux_sel), .A2(instr_rdata_i[9]), .ZN(
        n769) );
  OAI21_X1 U1025 ( .B1(regfile_alu_waddr_mux_sel), .B2(n770), .A(n769), .ZN(
        regfile_alu_waddr_id[2]) );
  INV_X1 U1040 ( .A(regfile_wdata_wb_i[7]), .ZN(n2182) );
  NAND2_X1 U1041 ( .A1(n53), .A2(n31), .ZN(n781) );
  AOI22_X1 U1042 ( .A1(n784), .A2(n2678), .B1(n615), .B2(csr_hwlp_data_i[7]), 
        .ZN(n780) );
  OAI211_X1 U1043 ( .C1(n814), .C2(n2182), .A(n781), .B(n780), .ZN(n782) );
  AOI21_X1 U1044 ( .B1(regfile_alu_wdata_fw_i[7]), .B2(n788), .A(n782), .ZN(
        n783) );
  INV_X1 U1045 ( .A(n783), .ZN(hwloop_cnt[7]) );
  INV_X1 U1046 ( .A(regfile_wdata_wb_i[10]), .ZN(n2215) );
  NAND2_X1 U1047 ( .A1(n53), .A2(n47), .ZN(n786) );
  AOI22_X1 U1048 ( .A1(n784), .A2(instr_rdata_i[30]), .B1(n615), .B2(
        csr_hwlp_data_i[10]), .ZN(n785) );
  OAI211_X1 U1049 ( .C1(n814), .C2(n2215), .A(n786), .B(n785), .ZN(n787) );
  AOI21_X1 U1050 ( .B1(regfile_alu_wdata_fw_i[10]), .B2(n788), .A(n787), .ZN(
        n789) );
  INV_X1 U1051 ( .A(n789), .ZN(hwloop_cnt[10]) );
  AOI22_X1 U1052 ( .A1(regfile_wdata_wb_i[7]), .A2(n2207), .B1(n2209), .B2(
        regfile_data_rb_id[7]), .ZN(n790) );
  INV_X1 U1053 ( .A(n790), .ZN(n791) );
  AOI21_X1 U1054 ( .B1(regfile_alu_wdata_fw_i[7]), .B2(n2205), .A(n791), .ZN(
        n2188) );
  XOR2_X1 U1057 ( .A(instr_rdata_i[17]), .B(regfile_waddr_wb_i[2]), .Z(n797)
         );
  XOR2_X1 U1058 ( .A(regfile_waddr_wb_i[1]), .B(n80), .Z(n796) );
  XOR2_X1 U1059 ( .A(regfile_waddr_wb_i[4]), .B(n116), .Z(n795) );
  NOR3_X1 U1060 ( .A1(n797), .A2(n796), .A3(n795), .ZN(n800) );
  XNOR2_X1 U1061 ( .A(regfile_waddr_wb_i[0]), .B(n113), .ZN(n799) );
  XNOR2_X1 U1062 ( .A(n33), .B(regfile_waddr_wb_i[3]), .ZN(n798) );
  NAND3_X1 U1063 ( .A1(n800), .A2(n799), .A3(n798), .ZN(n801) );
  NOR2_X1 U1064 ( .A1(n809), .A2(n801), .ZN(reg_d_wb_is_reg_a_id) );
  XOR2_X1 U1065 ( .A(n113), .B(regfile_alu_waddr_ex_o[0]), .Z(n804) );
  XOR2_X1 U1066 ( .A(regfile_alu_waddr_ex_o[3]), .B(n33), .Z(n803) );
  XOR2_X1 U1067 ( .A(regfile_alu_waddr_ex_o[1]), .B(n80), .Z(n802) );
  NOR3_X1 U1068 ( .A1(n804), .A2(n803), .A3(n802), .ZN(n807) );
  XNOR2_X1 U1069 ( .A(n110), .B(regfile_alu_waddr_ex_o[2]), .ZN(n806) );
  XNOR2_X1 U1070 ( .A(n116), .B(regfile_alu_waddr_ex_o[4]), .ZN(n805) );
  NAND3_X1 U1071 ( .A1(n807), .A2(n806), .A3(n805), .ZN(n808) );
  NOR2_X1 U1072 ( .A1(n809), .A2(n808), .ZN(reg_d_alu_is_reg_a_id) );
  INV_X1 U1073 ( .A(n810), .ZN(n2451) );
  NAND3_X1 U1074 ( .A1(n1032), .A2(jump_in_id[1]), .A3(jump_in_id[0]), .ZN(
        n2569) );
  INV_X1 U1076 ( .A(regfile_wdata_wb_i[16]), .ZN(n1849) );
  NAND2_X1 U1077 ( .A1(regfile_alu_wdata_fw_i[16]), .A2(n811), .ZN(n813) );
  AOI22_X1 U1078 ( .A1(n53), .A2(n38), .B1(csr_hwlp_data_i[16]), .B2(n615), 
        .ZN(n812) );
  OAI211_X1 U1079 ( .C1(n1849), .C2(n814), .A(n813), .B(n812), .ZN(
        hwloop_cnt[16]) );
  OAI22_X1 U1080 ( .A1(n860), .A2(csr_hwlp_data_i[0]), .B1(n854), .B2(
        pc_id_i[0]), .ZN(n815) );
  INV_X1 U1081 ( .A(n815), .ZN(hwloop_end[0]) );
  INV_X1 U1082 ( .A(n854), .ZN(n897) );
  XOR2_X1 U1083 ( .A(n816), .B(pc_id_i[1]), .Z(n902) );
  OAI22_X1 U1084 ( .A1(csr_hwlp_data_i[1]), .A2(n897), .B1(n854), .B2(n902), 
        .ZN(n817) );
  INV_X1 U1085 ( .A(n817), .ZN(hwloop_end[1]) );
  FA_X1 U1086 ( .A(pc_id_i[2]), .B(n819), .CI(n818), .CO(n823), .S(n906) );
  OAI22_X1 U1087 ( .A1(n897), .A2(csr_hwlp_data_i[2]), .B1(n854), .B2(n906), 
        .ZN(n820) );
  INV_X1 U1088 ( .A(n820), .ZN(hwloop_end[2]) );
  XNOR2_X1 U1089 ( .A(n823), .B(n822), .ZN(n908) );
  OAI22_X1 U1090 ( .A1(n860), .A2(csr_hwlp_data_i[3]), .B1(n854), .B2(n908), 
        .ZN(n824) );
  INV_X1 U1091 ( .A(n824), .ZN(hwloop_end[3]) );
  FA_X1 U1092 ( .A(pc_id_i[4]), .B(n826), .CI(n825), .CO(n828), .S(n912) );
  OAI22_X1 U1093 ( .A1(n897), .A2(csr_hwlp_data_i[4]), .B1(n854), .B2(n912), 
        .ZN(n827) );
  INV_X1 U1094 ( .A(n827), .ZN(hwloop_end[4]) );
  FA_X1 U1095 ( .A(pc_id_i[5]), .B(n829), .CI(n828), .CO(n833), .S(n916) );
  OAI22_X1 U1096 ( .A1(n860), .A2(csr_hwlp_data_i[5]), .B1(n854), .B2(n916), 
        .ZN(n830) );
  INV_X1 U1097 ( .A(n830), .ZN(hwloop_end[5]) );
  XNOR2_X1 U1098 ( .A(n831), .B(pc_id_i[6]), .ZN(n832) );
  XNOR2_X1 U1099 ( .A(n833), .B(n832), .ZN(n920) );
  OAI22_X1 U1100 ( .A1(n860), .A2(csr_hwlp_data_i[6]), .B1(n854), .B2(n920), 
        .ZN(n834) );
  INV_X1 U1101 ( .A(n834), .ZN(hwloop_end[6]) );
  XNOR2_X1 U1102 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U1103 ( .A(n838), .B(n837), .ZN(n922) );
  OAI22_X1 U1104 ( .A1(n860), .A2(csr_hwlp_data_i[7]), .B1(n854), .B2(n922), 
        .ZN(n839) );
  INV_X1 U1105 ( .A(n839), .ZN(hwloop_end[7]) );
  FA_X1 U1106 ( .A(pc_id_i[8]), .B(n841), .CI(n840), .CO(n843), .S(n924) );
  OAI22_X1 U1107 ( .A1(n860), .A2(csr_hwlp_data_i[8]), .B1(n854), .B2(n924), 
        .ZN(n842) );
  INV_X1 U1108 ( .A(n842), .ZN(hwloop_end[8]) );
  FA_X1 U1109 ( .A(pc_id_i[9]), .B(n844), .CI(n843), .CO(n846), .S(n928) );
  OAI22_X1 U1110 ( .A1(n860), .A2(csr_hwlp_data_i[9]), .B1(n854), .B2(n928), 
        .ZN(n845) );
  INV_X1 U1111 ( .A(n845), .ZN(hwloop_end[9]) );
  FA_X1 U1112 ( .A(pc_id_i[10]), .B(n847), .CI(n846), .CO(n849), .S(n932) );
  OAI22_X1 U1113 ( .A1(n860), .A2(csr_hwlp_data_i[10]), .B1(n854), .B2(n932), 
        .ZN(n848) );
  INV_X1 U1114 ( .A(n848), .ZN(hwloop_end[10]) );
  FA_X1 U1115 ( .A(pc_id_i[11]), .B(n850), .CI(n849), .CO(n852), .S(n934) );
  OAI22_X1 U1116 ( .A1(n934), .A2(n854), .B1(csr_hwlp_data_i[11]), .B2(n860), 
        .ZN(n851) );
  INV_X1 U1117 ( .A(n851), .ZN(hwloop_end[11]) );
  FA_X1 U1118 ( .A(pc_id_i[12]), .B(n853), .CI(n852), .CO(n856), .S(n936) );
  OAI22_X1 U1119 ( .A1(n936), .A2(n854), .B1(csr_hwlp_data_i[12]), .B2(n860), 
        .ZN(n855) );
  INV_X1 U1120 ( .A(n855), .ZN(hwloop_end[12]) );
  HA_X1 U1121 ( .A(n856), .B(pc_id_i[13]), .CO(n859), .S(n938) );
  OAI22_X1 U1122 ( .A1(n938), .A2(n854), .B1(csr_hwlp_data_i[13]), .B2(n860), 
        .ZN(n857) );
  INV_X1 U1123 ( .A(n857), .ZN(hwloop_end[13]) );
  INV_X1 U1124 ( .A(pc_id_i[14]), .ZN(n858) );
  OAI22_X1 U1125 ( .A1(n940), .A2(n854), .B1(csr_hwlp_data_i[14]), .B2(n860), 
        .ZN(n861) );
  INV_X1 U1126 ( .A(n861), .ZN(hwloop_end[14]) );
  XNOR2_X1 U1127 ( .A(n862), .B(pc_id_i[15]), .ZN(n942) );
  OAI22_X1 U1128 ( .A1(n942), .A2(n854), .B1(csr_hwlp_data_i[15]), .B2(n860), 
        .ZN(n863) );
  INV_X1 U1129 ( .A(n863), .ZN(hwloop_end[15]) );
  HA_X1 U1130 ( .A(n864), .B(pc_id_i[16]), .CO(n866), .S(n944) );
  OAI22_X1 U1131 ( .A1(n944), .A2(n854), .B1(csr_hwlp_data_i[16]), .B2(n860), 
        .ZN(n865) );
  INV_X1 U1132 ( .A(n865), .ZN(hwloop_end[16]) );
  HA_X1 U1133 ( .A(n866), .B(pc_id_i[17]), .CO(n868), .S(n947) );
  OAI22_X1 U1134 ( .A1(n947), .A2(n854), .B1(csr_hwlp_data_i[17]), .B2(n860), 
        .ZN(n867) );
  INV_X1 U1135 ( .A(n867), .ZN(hwloop_end[17]) );
  HA_X1 U1136 ( .A(n868), .B(pc_id_i[18]), .CO(n871), .S(n951) );
  OAI22_X1 U1137 ( .A1(n951), .A2(n854), .B1(n860), .B2(csr_hwlp_data_i[18]), 
        .ZN(n869) );
  INV_X1 U1138 ( .A(n869), .ZN(hwloop_end[18]) );
  INV_X1 U1139 ( .A(pc_id_i[19]), .ZN(n870) );
  XNOR2_X1 U1140 ( .A(n871), .B(n870), .ZN(n955) );
  OAI22_X1 U1141 ( .A1(n955), .A2(n854), .B1(csr_hwlp_data_i[19]), .B2(n860), 
        .ZN(n872) );
  INV_X1 U1142 ( .A(n872), .ZN(hwloop_end[19]) );
  XNOR2_X1 U1143 ( .A(n873), .B(pc_id_i[20]), .ZN(n959) );
  OAI22_X1 U1144 ( .A1(n959), .A2(n854), .B1(csr_hwlp_data_i[20]), .B2(n860), 
        .ZN(n874) );
  INV_X1 U1145 ( .A(n874), .ZN(hwloop_end[20]) );
  HA_X1 U1146 ( .A(n875), .B(pc_id_i[21]), .CO(n877), .S(n963) );
  OAI22_X1 U1147 ( .A1(n963), .A2(n854), .B1(csr_hwlp_data_i[21]), .B2(n860), 
        .ZN(n876) );
  INV_X1 U1148 ( .A(n876), .ZN(hwloop_end[21]) );
  HA_X1 U1149 ( .A(n877), .B(pc_id_i[22]), .CO(n880), .S(n967) );
  OAI22_X1 U1150 ( .A1(n967), .A2(n854), .B1(csr_hwlp_data_i[22]), .B2(n860), 
        .ZN(n878) );
  INV_X1 U1151 ( .A(n878), .ZN(hwloop_end[22]) );
  INV_X1 U1152 ( .A(pc_id_i[23]), .ZN(n879) );
  OAI22_X1 U1153 ( .A1(n971), .A2(n854), .B1(csr_hwlp_data_i[23]), .B2(n860), 
        .ZN(n881) );
  INV_X1 U1154 ( .A(n881), .ZN(hwloop_end[23]) );
  XNOR2_X1 U1155 ( .A(n882), .B(pc_id_i[24]), .ZN(n975) );
  OAI22_X1 U1156 ( .A1(n975), .A2(n854), .B1(csr_hwlp_data_i[24]), .B2(n897), 
        .ZN(n883) );
  INV_X1 U1157 ( .A(n883), .ZN(hwloop_end[24]) );
  HA_X1 U1158 ( .A(n884), .B(pc_id_i[25]), .CO(n886), .S(n979) );
  OAI22_X1 U1159 ( .A1(n979), .A2(n854), .B1(csr_hwlp_data_i[25]), .B2(n897), 
        .ZN(n885) );
  INV_X1 U1160 ( .A(n885), .ZN(hwloop_end[25]) );
  HA_X1 U1161 ( .A(n886), .B(pc_id_i[26]), .CO(n889), .S(n983) );
  OAI22_X1 U1162 ( .A1(n983), .A2(n854), .B1(csr_hwlp_data_i[26]), .B2(n897), 
        .ZN(n887) );
  INV_X1 U1163 ( .A(n887), .ZN(hwloop_end[26]) );
  XNOR2_X1 U1164 ( .A(n889), .B(n888), .ZN(n987) );
  OAI22_X1 U1165 ( .A1(n987), .A2(n854), .B1(csr_hwlp_data_i[27]), .B2(n897), 
        .ZN(n890) );
  INV_X1 U1166 ( .A(n890), .ZN(hwloop_end[27]) );
  OAI22_X1 U1167 ( .A1(n991), .A2(n854), .B1(csr_hwlp_data_i[28]), .B2(n897), 
        .ZN(n892) );
  INV_X1 U1168 ( .A(n892), .ZN(hwloop_end[28]) );
  HA_X1 U1169 ( .A(n893), .B(pc_id_i[29]), .CO(n895), .S(n996) );
  OAI22_X1 U1170 ( .A1(n996), .A2(n854), .B1(csr_hwlp_data_i[29]), .B2(n897), 
        .ZN(n894) );
  INV_X1 U1171 ( .A(n894), .ZN(hwloop_end[29]) );
  HA_X1 U1172 ( .A(n895), .B(pc_id_i[30]), .CO(n210), .S(n1001) );
  OAI22_X1 U1173 ( .A1(n1001), .A2(n854), .B1(csr_hwlp_data_i[30]), .B2(n897), 
        .ZN(n896) );
  INV_X1 U1174 ( .A(n896), .ZN(hwloop_end[30]) );
  OAI22_X1 U1175 ( .A1(n898), .A2(n854), .B1(csr_hwlp_data_i[31]), .B2(n897), 
        .ZN(n899) );
  INV_X1 U1176 ( .A(n899), .ZN(hwloop_end[31]) );
  AOI222_X1 U1177 ( .A1(n211), .A2(csr_hwlp_data_i[0]), .B1(n900), .B2(
        pc_if_i[0]), .C1(n1000), .C2(pc_id_i[0]), .ZN(n901) );
  INV_X1 U1178 ( .A(n901), .ZN(hwloop_start[0]) );
  INV_X1 U1179 ( .A(csr_hwlp_data_i[1]), .ZN(n905) );
  NAND2_X1 U1180 ( .A1(n1000), .A2(n902), .ZN(n904) );
  NAND2_X1 U1181 ( .A1(n900), .A2(pc_if_i[1]), .ZN(n903) );
  OAI211_X1 U1182 ( .C1(n1005), .C2(n905), .A(n904), .B(n903), .ZN(
        hwloop_start[1]) );
  AOI222_X1 U1184 ( .A1(n211), .A2(csr_hwlp_data_i[2]), .B1(n900), .B2(
        pc_if_i[2]), .C1(n1000), .C2(n906), .ZN(n907) );
  INV_X1 U1185 ( .A(n907), .ZN(hwloop_start[2]) );
  INV_X1 U1186 ( .A(csr_hwlp_data_i[3]), .ZN(n911) );
  NAND2_X1 U1187 ( .A1(n1000), .A2(n908), .ZN(n910) );
  NAND2_X1 U1188 ( .A1(n900), .A2(pc_if_i[3]), .ZN(n909) );
  OAI211_X1 U1189 ( .C1(n1005), .C2(n911), .A(n910), .B(n909), .ZN(
        hwloop_start[3]) );
  INV_X1 U1190 ( .A(csr_hwlp_data_i[4]), .ZN(n915) );
  NAND2_X1 U1191 ( .A1(n1000), .A2(n912), .ZN(n914) );
  NAND2_X1 U1192 ( .A1(n900), .A2(pc_if_i[4]), .ZN(n913) );
  OAI211_X1 U1193 ( .C1(n1005), .C2(n915), .A(n914), .B(n913), .ZN(
        hwloop_start[4]) );
  INV_X1 U1194 ( .A(csr_hwlp_data_i[5]), .ZN(n919) );
  NAND2_X1 U1195 ( .A1(n1000), .A2(n916), .ZN(n918) );
  NAND2_X1 U1196 ( .A1(n900), .A2(pc_if_i[5]), .ZN(n917) );
  OAI211_X1 U1197 ( .C1(n1005), .C2(n919), .A(n918), .B(n917), .ZN(
        hwloop_start[5]) );
  AOI222_X1 U1198 ( .A1(n211), .A2(csr_hwlp_data_i[6]), .B1(n900), .B2(
        pc_if_i[6]), .C1(n1000), .C2(n920), .ZN(n921) );
  INV_X1 U1199 ( .A(n921), .ZN(hwloop_start[6]) );
  AOI222_X1 U1200 ( .A1(n211), .A2(csr_hwlp_data_i[7]), .B1(n900), .B2(
        pc_if_i[7]), .C1(n1000), .C2(n922), .ZN(n923) );
  INV_X1 U1201 ( .A(n923), .ZN(hwloop_start[7]) );
  INV_X1 U1202 ( .A(csr_hwlp_data_i[8]), .ZN(n927) );
  NAND2_X1 U1203 ( .A1(n1000), .A2(n924), .ZN(n926) );
  NAND2_X1 U1204 ( .A1(n900), .A2(pc_if_i[8]), .ZN(n925) );
  OAI211_X1 U1205 ( .C1(n1005), .C2(n927), .A(n926), .B(n925), .ZN(
        hwloop_start[8]) );
  INV_X1 U1206 ( .A(csr_hwlp_data_i[9]), .ZN(n931) );
  NAND2_X1 U1207 ( .A1(n1000), .A2(n928), .ZN(n930) );
  NAND2_X1 U1208 ( .A1(n900), .A2(pc_if_i[9]), .ZN(n929) );
  OAI211_X1 U1209 ( .C1(n1005), .C2(n931), .A(n930), .B(n929), .ZN(
        hwloop_start[9]) );
  AOI222_X1 U1210 ( .A1(n211), .A2(csr_hwlp_data_i[10]), .B1(n900), .B2(
        pc_if_i[10]), .C1(n1000), .C2(n932), .ZN(n933) );
  INV_X1 U1211 ( .A(n933), .ZN(hwloop_start[10]) );
  AOI222_X1 U1212 ( .A1(n211), .A2(csr_hwlp_data_i[11]), .B1(n900), .B2(
        pc_if_i[11]), .C1(n1000), .C2(n934), .ZN(n935) );
  INV_X1 U1213 ( .A(n935), .ZN(hwloop_start[11]) );
  AOI222_X1 U1214 ( .A1(n211), .A2(csr_hwlp_data_i[12]), .B1(n900), .B2(
        pc_if_i[12]), .C1(n1000), .C2(n936), .ZN(n937) );
  INV_X1 U1215 ( .A(n937), .ZN(hwloop_start[12]) );
  AOI222_X1 U1216 ( .A1(n211), .A2(csr_hwlp_data_i[13]), .B1(n900), .B2(
        pc_if_i[13]), .C1(n1000), .C2(n938), .ZN(n939) );
  INV_X1 U1217 ( .A(n939), .ZN(hwloop_start[13]) );
  AOI222_X1 U1218 ( .A1(n211), .A2(csr_hwlp_data_i[14]), .B1(n900), .B2(
        pc_if_i[14]), .C1(n1000), .C2(n940), .ZN(n941) );
  INV_X1 U1219 ( .A(n941), .ZN(hwloop_start[14]) );
  AOI222_X1 U1220 ( .A1(n211), .A2(csr_hwlp_data_i[15]), .B1(n900), .B2(
        pc_if_i[15]), .C1(n1000), .C2(n942), .ZN(n943) );
  INV_X1 U1221 ( .A(n943), .ZN(hwloop_start[15]) );
  AOI222_X1 U1222 ( .A1(n211), .A2(csr_hwlp_data_i[16]), .B1(n900), .B2(
        pc_if_i[16]), .C1(n1000), .C2(n944), .ZN(n946) );
  INV_X1 U1223 ( .A(n946), .ZN(hwloop_start[16]) );
  INV_X1 U1224 ( .A(csr_hwlp_data_i[17]), .ZN(n950) );
  NAND2_X1 U1225 ( .A1(n947), .A2(n1000), .ZN(n949) );
  NAND2_X1 U1226 ( .A1(n900), .A2(pc_if_i[17]), .ZN(n948) );
  OAI211_X1 U1227 ( .C1(n1005), .C2(n950), .A(n949), .B(n948), .ZN(
        hwloop_start[17]) );
  INV_X1 U1228 ( .A(csr_hwlp_data_i[18]), .ZN(n954) );
  NAND2_X1 U1229 ( .A1(n951), .A2(n1000), .ZN(n953) );
  NAND2_X1 U1230 ( .A1(n900), .A2(pc_if_i[18]), .ZN(n952) );
  OAI211_X1 U1231 ( .C1(n1005), .C2(n954), .A(n953), .B(n952), .ZN(
        hwloop_start[18]) );
  INV_X1 U1232 ( .A(csr_hwlp_data_i[19]), .ZN(n958) );
  NAND2_X1 U1233 ( .A1(n955), .A2(n1000), .ZN(n957) );
  NAND2_X1 U1234 ( .A1(n900), .A2(pc_if_i[19]), .ZN(n956) );
  OAI211_X1 U1235 ( .C1(n1005), .C2(n958), .A(n957), .B(n956), .ZN(
        hwloop_start[19]) );
  INV_X1 U1236 ( .A(csr_hwlp_data_i[20]), .ZN(n962) );
  NAND2_X1 U1237 ( .A1(n959), .A2(n995), .ZN(n961) );
  NAND2_X1 U1238 ( .A1(n900), .A2(pc_if_i[20]), .ZN(n960) );
  OAI211_X1 U1239 ( .C1(n1005), .C2(n962), .A(n961), .B(n960), .ZN(
        hwloop_start[20]) );
  INV_X1 U1240 ( .A(csr_hwlp_data_i[21]), .ZN(n966) );
  NAND2_X1 U1241 ( .A1(n963), .A2(n995), .ZN(n965) );
  NAND2_X1 U1242 ( .A1(n900), .A2(pc_if_i[21]), .ZN(n964) );
  OAI211_X1 U1243 ( .C1(n1005), .C2(n966), .A(n965), .B(n964), .ZN(
        hwloop_start[21]) );
  INV_X1 U1244 ( .A(csr_hwlp_data_i[22]), .ZN(n970) );
  NAND2_X1 U1245 ( .A1(n967), .A2(n995), .ZN(n969) );
  NAND2_X1 U1246 ( .A1(n900), .A2(pc_if_i[22]), .ZN(n968) );
  OAI211_X1 U1247 ( .C1(n1005), .C2(n970), .A(n969), .B(n968), .ZN(
        hwloop_start[22]) );
  NAND2_X1 U1248 ( .A1(n971), .A2(n995), .ZN(n973) );
  NAND2_X1 U1249 ( .A1(n900), .A2(pc_if_i[23]), .ZN(n972) );
  OAI211_X1 U1250 ( .C1(n1005), .C2(n974), .A(n973), .B(n972), .ZN(
        hwloop_start[23]) );
  INV_X1 U1251 ( .A(csr_hwlp_data_i[24]), .ZN(n978) );
  NAND2_X1 U1252 ( .A1(n975), .A2(n995), .ZN(n977) );
  NAND2_X1 U1253 ( .A1(n900), .A2(pc_if_i[24]), .ZN(n976) );
  OAI211_X1 U1254 ( .C1(n1005), .C2(n978), .A(n977), .B(n976), .ZN(
        hwloop_start[24]) );
  INV_X1 U1255 ( .A(csr_hwlp_data_i[25]), .ZN(n982) );
  NAND2_X1 U1256 ( .A1(n979), .A2(n995), .ZN(n981) );
  NAND2_X1 U1257 ( .A1(n900), .A2(pc_if_i[25]), .ZN(n980) );
  OAI211_X1 U1258 ( .C1(n1005), .C2(n982), .A(n981), .B(n980), .ZN(
        hwloop_start[25]) );
  INV_X1 U1259 ( .A(csr_hwlp_data_i[26]), .ZN(n986) );
  NAND2_X1 U1260 ( .A1(n983), .A2(n995), .ZN(n985) );
  NAND2_X1 U1261 ( .A1(n900), .A2(pc_if_i[26]), .ZN(n984) );
  OAI211_X1 U1262 ( .C1(n1005), .C2(n986), .A(n985), .B(n984), .ZN(
        hwloop_start[26]) );
  INV_X1 U1263 ( .A(csr_hwlp_data_i[27]), .ZN(n990) );
  NAND2_X1 U1264 ( .A1(n987), .A2(n995), .ZN(n989) );
  NAND2_X1 U1265 ( .A1(n900), .A2(pc_if_i[27]), .ZN(n988) );
  OAI211_X1 U1266 ( .C1(n1005), .C2(n990), .A(n989), .B(n988), .ZN(
        hwloop_start[27]) );
  INV_X1 U1267 ( .A(csr_hwlp_data_i[28]), .ZN(n994) );
  NAND2_X1 U1268 ( .A1(n991), .A2(n995), .ZN(n993) );
  NAND2_X1 U1269 ( .A1(n900), .A2(pc_if_i[28]), .ZN(n992) );
  OAI211_X1 U1270 ( .C1(n1005), .C2(n994), .A(n993), .B(n992), .ZN(
        hwloop_start[28]) );
  INV_X1 U1271 ( .A(csr_hwlp_data_i[29]), .ZN(n999) );
  NAND2_X1 U1272 ( .A1(n996), .A2(n995), .ZN(n998) );
  NAND2_X1 U1273 ( .A1(n900), .A2(pc_if_i[29]), .ZN(n997) );
  OAI211_X1 U1274 ( .C1(n1005), .C2(n999), .A(n998), .B(n997), .ZN(
        hwloop_start[29]) );
  INV_X1 U1275 ( .A(csr_hwlp_data_i[30]), .ZN(n1004) );
  NAND2_X1 U1276 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  NAND2_X1 U1277 ( .A1(n900), .A2(pc_if_i[30]), .ZN(n1002) );
  OAI211_X1 U1278 ( .C1(n1005), .C2(n1004), .A(n1003), .B(n1002), .ZN(
        hwloop_start[30]) );
  NAND2_X1 U1279 ( .A1(n1032), .A2(regfile_alu_we_id), .ZN(n2452) );
  NAND2_X1 U1281 ( .A1(regfile_alu_waddr_mux_sel), .A2(instr_rdata_i[10]), 
        .ZN(n1006) );
  OAI21_X1 U1282 ( .B1(regfile_alu_waddr_mux_sel), .B2(n1914), .A(n1006), .ZN(
        regfile_alu_waddr_id[3]) );
  NAND2_X1 U1285 ( .A1(regfile_alu_waddr_mux_sel), .A2(instr_rdata_i[8]), .ZN(
        n1007) );
  OAI21_X1 U1286 ( .B1(regfile_alu_waddr_mux_sel), .B2(n1008), .A(n1007), .ZN(
        regfile_alu_waddr_id[1]) );
  NAND2_X1 U1288 ( .A1(regfile_alu_waddr_mux_sel), .A2(instr_rdata_i[11]), 
        .ZN(n1009) );
  OAI21_X1 U1289 ( .B1(regfile_alu_waddr_mux_sel), .B2(n1010), .A(n1009), .ZN(
        regfile_alu_waddr_id[4]) );
  XOR2_X1 U1291 ( .A(regfile_alu_waddr_ex_o[2]), .B(instr_rdata_i[22]), .Z(
        n1016) );
  XOR2_X1 U1292 ( .A(regfile_alu_waddr_ex_o[3]), .B(instr_rdata_i[23]), .Z(
        n1015) );
  XNOR2_X1 U1293 ( .A(n2604), .B(regfile_alu_waddr_ex_o[4]), .ZN(n1013) );
  XNOR2_X1 U1294 ( .A(instr_rdata_i[20]), .B(regfile_alu_waddr_ex_o[0]), .ZN(
        n1012) );
  XNOR2_X1 U1295 ( .A(instr_rdata_i[21]), .B(regfile_alu_waddr_ex_o[1]), .ZN(
        n1011) );
  NAND3_X1 U1296 ( .A1(n1013), .A2(n1012), .A3(n1011), .ZN(n1014) );
  NOR4_X1 U1297 ( .A1(n1030), .A2(n1016), .A3(n1015), .A4(n1014), .ZN(
        reg_d_alu_is_reg_b_id) );
  XNOR2_X1 U1298 ( .A(n1637), .B(regfile_waddr_wb_i[3]), .ZN(n1019) );
  XNOR2_X1 U1299 ( .A(n1634), .B(regfile_waddr_wb_i[0]), .ZN(n1018) );
  XNOR2_X1 U1300 ( .A(n1635), .B(regfile_waddr_wb_i[1]), .ZN(n1017) );
  NAND3_X1 U1301 ( .A1(n1019), .A2(n1018), .A3(n1017), .ZN(n1022) );
  XOR2_X1 U1302 ( .A(regfile_waddr_wb_i[4]), .B(n1638), .Z(n1021) );
  XOR2_X1 U1303 ( .A(n1636), .B(regfile_waddr_wb_i[2]), .Z(n1020) );
  NOR4_X1 U1304 ( .A1(n1023), .A2(n1022), .A3(n1021), .A4(n1020), .ZN(
        reg_d_wb_is_reg_c_id) );
  AOI22_X1 U1305 ( .A1(n1991), .A2(regfile_waddr_wb_i[3]), .B1(
        regfile_waddr_wb_i[0]), .B2(n2467), .ZN(n1024) );
  OAI221_X1 U1306 ( .B1(n1991), .B2(regfile_waddr_wb_i[3]), .C1(n2467), .C2(
        regfile_waddr_wb_i[0]), .A(n1024), .ZN(n1029) );
  XOR2_X1 U1307 ( .A(regfile_waddr_wb_i[4]), .B(n2604), .Z(n1028) );
  OAI22_X1 U1308 ( .A1(n1984), .A2(regfile_waddr_wb_i[2]), .B1(n1738), .B2(
        regfile_waddr_wb_i[1]), .ZN(n1025) );
  AOI221_X1 U1309 ( .B1(n1984), .B2(regfile_waddr_wb_i[2]), .C1(
        regfile_waddr_wb_i[1]), .C2(n1738), .A(n1025), .ZN(n1026) );
  INV_X1 U1310 ( .A(n1026), .ZN(n1027) );
  NOR4_X1 U1311 ( .A1(n1030), .A2(n1029), .A3(n1028), .A4(n1027), .ZN(
        reg_d_wb_is_reg_b_id) );
  NAND2_X1 U1319 ( .A1(n1032), .A2(data_req_id), .ZN(n2570) );
  NAND2_X1 U1322 ( .A1(n2671), .A2(data_misaligned_i), .ZN(n2503) );
  NAND2_X1 U1323 ( .A1(n2427), .A2(n2503), .ZN(n1033) );
  MUX2_X1 U1324 ( .A(prepost_useincr_ex_o), .B(prepost_useincr), .S(n1033), 
        .Z(n1353) );
  OAI21_X1 U1325 ( .B1(n2451), .B2(n2597), .A(n2503), .ZN(n1276) );
  INV_X1 U1326 ( .A(data_load_event_id), .ZN(n1034) );
  MUX2_X1 U1331 ( .A(csr_access), .B(csr_access_ex_o), .S(n2427), .Z(n1626) );
  INV_X1 U1332 ( .A(mult_dot_en), .ZN(n1035) );
  AOI22_X1 U1339 ( .A1(regfile_wdata_wb_i[0]), .A2(n2207), .B1(n2209), .B2(
        regfile_data_rb_id[0]), .ZN(n1036) );
  INV_X1 U1340 ( .A(n1205), .ZN(n1046) );
  INV_X1 U1341 ( .A(alu_op_c_mux_sel[1]), .ZN(n1037) );
  NAND2_X1 U1342 ( .A1(n1037), .A2(alu_op_c_mux_sel[0]), .ZN(n1101) );
  OR2_X1 U1343 ( .A1(operand_c_fw_mux_sel[1]), .A2(operand_c_fw_mux_sel[0]), 
        .ZN(n2185) );
  INV_X1 U1344 ( .A(n2185), .ZN(n1228) );
  NAND2_X1 U1345 ( .A1(operand_c_fw_mux_sel[0]), .A2(operand_c_fw_mux_sel[1]), 
        .ZN(n2178) );
  NAND2_X1 U1346 ( .A1(n2185), .A2(n2178), .ZN(n2140) );
  INV_X1 U1347 ( .A(n2140), .ZN(n1125) );
  INV_X1 U1348 ( .A(n2178), .ZN(n1227) );
  AOI22_X1 U1349 ( .A1(regfile_data_rc_id[0]), .A2(n1125), .B1(
        regfile_wdata_wb_i[0]), .B2(n1227), .ZN(n1038) );
  INV_X1 U1350 ( .A(alu_op_c_mux_sel[0]), .ZN(n1039) );
  NAND2_X1 U1351 ( .A1(n1039), .A2(alu_op_c_mux_sel[1]), .ZN(n1103) );
  OR2_X1 U1352 ( .A1(n1041), .A2(n1040), .ZN(n1043) );
  AND2_X1 U1353 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  AOI22_X1 U1354 ( .A1(n1206), .A2(n1073), .B1(n1044), .B2(n1194), .ZN(n1045)
         );
  INV_X1 U1357 ( .A(n1229), .ZN(n1051) );
  INV_X1 U1358 ( .A(n1073), .ZN(n1132) );
  NOR2_X1 U1359 ( .A1(n2185), .A2(n1132), .ZN(n1089) );
  INV_X1 U1360 ( .A(regfile_data_rc_id[1]), .ZN(n1048) );
  NOR2_X1 U1361 ( .A1(n2178), .A2(n1132), .ZN(n1091) );
  AOI22_X1 U1362 ( .A1(regfile_wdata_wb_i[1]), .A2(n1091), .B1(n1194), .B2(
        jump_target_o[1]), .ZN(n1047) );
  OAI21_X1 U1363 ( .B1(n1048), .B2(n1160), .A(n1047), .ZN(n1049) );
  AOI21_X1 U1364 ( .B1(regfile_alu_wdata_fw_i[1]), .B2(n1089), .A(n1049), .ZN(
        n1050) );
  OAI21_X1 U1365 ( .B1(n1051), .B2(n1101), .A(n1050), .ZN(n2470) );
  INV_X1 U1367 ( .A(jump_target_o[2]), .ZN(n1055) );
  INV_X1 U1368 ( .A(regfile_data_rc_id[2]), .ZN(n1052) );
  OAI22_X1 U1369 ( .A1(n1053), .A2(n2178), .B1(n1052), .B2(n2140), .ZN(n1054)
         );
  OAI222_X1 U1370 ( .A1(n1103), .A2(n1055), .B1(n1132), .B2(n2147), .C1(n1101), 
        .C2(n2148), .ZN(n2471) );
  AOI22_X1 U1372 ( .A1(regfile_data_rc_id[3]), .A2(n1125), .B1(
        regfile_wdata_wb_i[3]), .B2(n1227), .ZN(n1056) );
  INV_X1 U1373 ( .A(n1056), .ZN(n1057) );
  AOI21_X1 U1374 ( .B1(regfile_alu_wdata_fw_i[3]), .B2(n1228), .A(n1057), .ZN(
        n1663) );
  INV_X1 U1375 ( .A(n1663), .ZN(n1058) );
  NAND2_X1 U1376 ( .A1(n1058), .A2(n1073), .ZN(n1060) );
  NAND2_X1 U1377 ( .A1(jump_target_o[3]), .A2(n1194), .ZN(n1059) );
  OAI211_X1 U1378 ( .C1(n2161), .C2(n1101), .A(n1060), .B(n1059), .ZN(n2472)
         );
  AOI22_X1 U1380 ( .A1(regfile_data_rc_id[4]), .A2(n1125), .B1(
        regfile_wdata_wb_i[4]), .B2(n1227), .ZN(n1061) );
  INV_X1 U1381 ( .A(n1061), .ZN(n1062) );
  AOI21_X1 U1382 ( .B1(regfile_alu_wdata_fw_i[4]), .B2(n1228), .A(n1062), .ZN(
        n1680) );
  INV_X1 U1383 ( .A(n1680), .ZN(n1064) );
  NAND2_X1 U1384 ( .A1(n1064), .A2(n1073), .ZN(n1066) );
  NAND2_X1 U1385 ( .A1(jump_target_o[4]), .A2(n1194), .ZN(n1065) );
  OAI211_X1 U1386 ( .C1(n1685), .C2(n1101), .A(n1066), .B(n1065), .ZN(n2473)
         );
  NAND2_X1 U1388 ( .A1(regfile_alu_wdata_fw_i[5]), .A2(n1228), .ZN(n1068) );
  AOI22_X1 U1389 ( .A1(n1125), .A2(regfile_data_rc_id[5]), .B1(
        regfile_wdata_wb_i[5]), .B2(n1227), .ZN(n1067) );
  NAND2_X1 U1390 ( .A1(n1068), .A2(n1067), .ZN(n1693) );
  AOI22_X1 U1391 ( .A1(n1693), .A2(n1073), .B1(jump_target_o[5]), .B2(n1194), 
        .ZN(n1070) );
  INV_X1 U1392 ( .A(n1101), .ZN(n1130) );
  NAND2_X1 U1393 ( .A1(n1692), .A2(n1130), .ZN(n1069) );
  NAND2_X1 U1394 ( .A1(n1070), .A2(n1069), .ZN(n2474) );
  AOI22_X1 U1396 ( .A1(regfile_data_rc_id[6]), .A2(n1125), .B1(n1227), .B2(
        regfile_wdata_wb_i[6]), .ZN(n1071) );
  INV_X1 U1397 ( .A(n1071), .ZN(n1072) );
  INV_X1 U1398 ( .A(n2176), .ZN(n1074) );
  NAND2_X1 U1399 ( .A1(n1074), .A2(n1073), .ZN(n1076) );
  NAND2_X1 U1400 ( .A1(jump_target_o[6]), .A2(n1194), .ZN(n1075) );
  OAI211_X1 U1401 ( .C1(n2173), .C2(n1101), .A(n1076), .B(n1075), .ZN(n2475)
         );
  INV_X1 U1403 ( .A(n1091), .ZN(n1085) );
  INV_X1 U1404 ( .A(n1160), .ZN(n1083) );
  AOI22_X1 U1405 ( .A1(n1083), .A2(regfile_data_rc_id[7]), .B1(n1194), .B2(
        jump_target_o[7]), .ZN(n1077) );
  OAI21_X1 U1406 ( .B1(n2182), .B2(n1085), .A(n1077), .ZN(n1078) );
  AOI21_X1 U1407 ( .B1(regfile_alu_wdata_fw_i[7]), .B2(n1089), .A(n1078), .ZN(
        n1079) );
  OAI21_X1 U1408 ( .B1(n2188), .B2(n1101), .A(n1079), .ZN(n2476) );
  AOI22_X1 U1410 ( .A1(n1083), .A2(regfile_data_rc_id[8]), .B1(n1194), .B2(
        jump_target_o[8]), .ZN(n1080) );
  OAI21_X1 U1411 ( .B1(n2195), .B2(n1085), .A(n1080), .ZN(n1081) );
  AOI21_X1 U1412 ( .B1(regfile_alu_wdata_fw_i[8]), .B2(n1089), .A(n1081), .ZN(
        n1082) );
  OAI21_X1 U1413 ( .B1(n2198), .B2(n1101), .A(n1082), .ZN(n2477) );
  AOI22_X1 U1415 ( .A1(n1083), .A2(regfile_data_rc_id[9]), .B1(n1194), .B2(
        jump_target_o[9]), .ZN(n1084) );
  OAI21_X1 U1416 ( .B1(n2201), .B2(n1085), .A(n1084), .ZN(n1086) );
  AOI21_X1 U1417 ( .B1(regfile_alu_wdata_fw_i[9]), .B2(n1089), .A(n1086), .ZN(
        n1087) );
  OAI21_X1 U1418 ( .B1(n2204), .B2(n1101), .A(n1087), .ZN(n2478) );
  NOR2_X1 U1420 ( .A1(n1882), .A2(n1101), .ZN(n1088) );
  OR2_X1 U1421 ( .A1(n1089), .A2(n1088), .ZN(n1193) );
  NAND2_X1 U1422 ( .A1(regfile_alu_wdata_fw_i[10]), .A2(n1193), .ZN(n1096) );
  AND2_X1 U1423 ( .A1(n2207), .A2(n1130), .ZN(n1090) );
  OR2_X1 U1424 ( .A1(n1091), .A2(n1090), .ZN(n1198) );
  INV_X1 U1425 ( .A(regfile_data_rc_id[10]), .ZN(n1093) );
  AOI22_X1 U1426 ( .A1(n1195), .A2(regfile_data_rb_id[10]), .B1(n1194), .B2(
        jump_target_o[10]), .ZN(n1092) );
  OAI21_X1 U1427 ( .B1(n1160), .B2(n1093), .A(n1092), .ZN(n1094) );
  AOI21_X1 U1428 ( .B1(regfile_wdata_wb_i[10]), .B2(n1198), .A(n1094), .ZN(
        n1095) );
  NAND2_X1 U1429 ( .A1(n1096), .A2(n1095), .ZN(n2480) );
  INV_X1 U1431 ( .A(jump_target_o[11]), .ZN(n1102) );
  AOI22_X1 U1432 ( .A1(regfile_wdata_wb_i[11]), .A2(n2207), .B1(n2209), .B2(
        regfile_data_rb_id[11]), .ZN(n1097) );
  INV_X1 U1433 ( .A(n1097), .ZN(n1098) );
  AOI21_X1 U1434 ( .B1(regfile_alu_wdata_fw_i[11]), .B2(n2205), .A(n1098), 
        .ZN(n1778) );
  AOI22_X1 U1435 ( .A1(regfile_wdata_wb_i[11]), .A2(n1227), .B1(n1125), .B2(
        regfile_data_rc_id[11]), .ZN(n1099) );
  INV_X1 U1436 ( .A(n1099), .ZN(n1100) );
  AOI21_X1 U1437 ( .B1(regfile_alu_wdata_fw_i[11]), .B2(n1228), .A(n1100), 
        .ZN(n1780) );
  OAI222_X1 U1438 ( .A1(n1103), .A2(n1102), .B1(n1101), .B2(n1778), .C1(n1132), 
        .C2(n1780), .ZN(n2482) );
  NAND2_X1 U1440 ( .A1(regfile_alu_wdata_fw_i[12]), .A2(n1193), .ZN(n1108) );
  INV_X1 U1441 ( .A(regfile_data_rc_id[12]), .ZN(n1105) );
  AOI22_X1 U1442 ( .A1(n1195), .A2(regfile_data_rb_id[12]), .B1(n1194), .B2(
        jump_target_o[12]), .ZN(n1104) );
  OAI21_X1 U1443 ( .B1(n1160), .B2(n1105), .A(n1104), .ZN(n1106) );
  AOI21_X1 U1444 ( .B1(regfile_wdata_wb_i[12]), .B2(n1198), .A(n1106), .ZN(
        n1107) );
  NAND2_X1 U1445 ( .A1(n1108), .A2(n1107), .ZN(n2483) );
  NAND2_X1 U1447 ( .A1(regfile_alu_wdata_fw_i[13]), .A2(n1193), .ZN(n1114) );
  INV_X1 U1448 ( .A(regfile_data_rc_id[13]), .ZN(n1111) );
  AOI22_X1 U1449 ( .A1(n1195), .A2(regfile_data_rb_id[13]), .B1(n1194), .B2(
        jump_target_o[13]), .ZN(n1110) );
  OAI21_X1 U1450 ( .B1(n1160), .B2(n1111), .A(n1110), .ZN(n1112) );
  AOI21_X1 U1451 ( .B1(regfile_wdata_wb_i[13]), .B2(n1198), .A(n1112), .ZN(
        n1113) );
  NAND2_X1 U1452 ( .A1(n1114), .A2(n1113), .ZN(n2484) );
  NAND2_X1 U1454 ( .A1(regfile_alu_wdata_fw_i[14]), .A2(n1193), .ZN(n1119) );
  INV_X1 U1455 ( .A(regfile_data_rc_id[14]), .ZN(n1116) );
  AOI22_X1 U1456 ( .A1(n1195), .A2(regfile_data_rb_id[14]), .B1(n1194), .B2(
        jump_target_o[14]), .ZN(n1115) );
  OAI21_X1 U1457 ( .B1(n1160), .B2(n1116), .A(n1115), .ZN(n1117) );
  AOI21_X1 U1458 ( .B1(regfile_wdata_wb_i[14]), .B2(n1198), .A(n1117), .ZN(
        n1118) );
  NAND2_X1 U1459 ( .A1(n1119), .A2(n1118), .ZN(n2485) );
  NAND2_X1 U1461 ( .A1(n2663), .A2(n1193), .ZN(n1124) );
  INV_X1 U1462 ( .A(regfile_data_rc_id[15]), .ZN(n1121) );
  AOI22_X1 U1463 ( .A1(n1195), .A2(regfile_data_rb_id[15]), .B1(n1194), .B2(
        jump_target_o[15]), .ZN(n1120) );
  OAI21_X1 U1464 ( .B1(n1160), .B2(n1121), .A(n1120), .ZN(n1122) );
  AOI21_X1 U1465 ( .B1(regfile_wdata_wb_i[15]), .B2(n1198), .A(n1122), .ZN(
        n1123) );
  NAND2_X1 U1466 ( .A1(n1124), .A2(n1123), .ZN(n2486) );
  NAND2_X1 U1468 ( .A1(regfile_alu_wdata_fw_i[16]), .A2(n1228), .ZN(n1127) );
  AOI22_X1 U1469 ( .A1(regfile_wdata_wb_i[16]), .A2(n1227), .B1(n1125), .B2(
        regfile_data_rc_id[16]), .ZN(n1126) );
  NAND2_X1 U1470 ( .A1(n1127), .A2(n1126), .ZN(n1867) );
  INV_X1 U1471 ( .A(n1867), .ZN(n1133) );
  NAND2_X1 U1472 ( .A1(regfile_alu_wdata_fw_i[16]), .A2(n2205), .ZN(n1129) );
  AOI22_X1 U1473 ( .A1(regfile_wdata_wb_i[16]), .A2(n2207), .B1(n2209), .B2(
        regfile_data_rb_id[16]), .ZN(n1128) );
  NAND2_X1 U1474 ( .A1(n1129), .A2(n1128), .ZN(n1866) );
  AOI22_X1 U1475 ( .A1(n1866), .A2(n1130), .B1(jump_target_o[16]), .B2(n1194), 
        .ZN(n1131) );
  OAI21_X1 U1476 ( .B1(n1133), .B2(n1132), .A(n1131), .ZN(n2487) );
  NAND2_X1 U1478 ( .A1(regfile_alu_wdata_fw_i[17]), .A2(n1193), .ZN(n1138) );
  INV_X1 U1479 ( .A(regfile_data_rc_id[17]), .ZN(n1135) );
  AOI22_X1 U1480 ( .A1(n1195), .A2(regfile_data_rb_id[17]), .B1(n1194), .B2(
        jump_target_o[17]), .ZN(n1134) );
  OAI21_X1 U1481 ( .B1(n1160), .B2(n1135), .A(n1134), .ZN(n1136) );
  AOI21_X1 U1482 ( .B1(regfile_wdata_wb_i[17]), .B2(n1198), .A(n1136), .ZN(
        n1137) );
  NAND2_X1 U1483 ( .A1(n1138), .A2(n1137), .ZN(n2488) );
  NAND2_X1 U1485 ( .A1(regfile_alu_wdata_fw_i[18]), .A2(n1193), .ZN(n1143) );
  INV_X1 U1486 ( .A(regfile_data_rc_id[18]), .ZN(n1140) );
  AOI22_X1 U1487 ( .A1(n1195), .A2(regfile_data_rb_id[18]), .B1(n1194), .B2(
        jump_target_o[18]), .ZN(n1139) );
  OAI21_X1 U1488 ( .B1(n1160), .B2(n1140), .A(n1139), .ZN(n1141) );
  AOI21_X1 U1489 ( .B1(regfile_wdata_wb_i[18]), .B2(n1198), .A(n1141), .ZN(
        n1142) );
  NAND2_X1 U1490 ( .A1(n1143), .A2(n1142), .ZN(n2489) );
  NAND2_X1 U1492 ( .A1(regfile_alu_wdata_fw_i[19]), .A2(n1193), .ZN(n1147) );
  INV_X1 U1493 ( .A(regfile_data_rc_id[19]), .ZN(n2303) );
  AOI22_X1 U1494 ( .A1(n1195), .A2(regfile_data_rb_id[19]), .B1(n1194), .B2(
        jump_target_o[19]), .ZN(n1144) );
  OAI21_X1 U1495 ( .B1(n1160), .B2(n2303), .A(n1144), .ZN(n1145) );
  AOI21_X1 U1496 ( .B1(regfile_wdata_wb_i[19]), .B2(n1198), .A(n1145), .ZN(
        n1146) );
  NAND2_X1 U1497 ( .A1(n1147), .A2(n1146), .ZN(n2490) );
  NAND2_X1 U1499 ( .A1(regfile_alu_wdata_fw_i[20]), .A2(n1193), .ZN(n1151) );
  INV_X1 U1500 ( .A(regfile_data_rc_id[20]), .ZN(n2312) );
  AOI22_X1 U1501 ( .A1(n1195), .A2(regfile_data_rb_id[20]), .B1(n1194), .B2(
        jump_target_o[20]), .ZN(n1148) );
  OAI21_X1 U1502 ( .B1(n1160), .B2(n2312), .A(n1148), .ZN(n1149) );
  AOI21_X1 U1503 ( .B1(regfile_wdata_wb_i[20]), .B2(n1198), .A(n1149), .ZN(
        n1150) );
  NAND2_X1 U1504 ( .A1(n1151), .A2(n1150), .ZN(n2491) );
  NAND2_X1 U1506 ( .A1(regfile_alu_wdata_fw_i[21]), .A2(n1193), .ZN(n1155) );
  INV_X1 U1507 ( .A(regfile_data_rc_id[21]), .ZN(n2321) );
  AOI22_X1 U1508 ( .A1(n1195), .A2(regfile_data_rb_id[21]), .B1(n1194), .B2(
        jump_target_o[21]), .ZN(n1152) );
  OAI21_X1 U1509 ( .B1(n1160), .B2(n2321), .A(n1152), .ZN(n1153) );
  AOI21_X1 U1510 ( .B1(regfile_wdata_wb_i[21]), .B2(n1198), .A(n1153), .ZN(
        n1154) );
  NAND2_X1 U1511 ( .A1(n1155), .A2(n1154), .ZN(n2492) );
  NAND2_X1 U1513 ( .A1(regfile_alu_wdata_fw_i[22]), .A2(n1193), .ZN(n1159) );
  INV_X1 U1514 ( .A(regfile_data_rc_id[22]), .ZN(n2330) );
  AOI22_X1 U1515 ( .A1(n1195), .A2(regfile_data_rb_id[22]), .B1(n1194), .B2(
        jump_target_o[22]), .ZN(n1156) );
  OAI21_X1 U1516 ( .B1(n1160), .B2(n2330), .A(n1156), .ZN(n1157) );
  AOI21_X1 U1517 ( .B1(regfile_wdata_wb_i[22]), .B2(n1198), .A(n1157), .ZN(
        n1158) );
  NAND2_X1 U1518 ( .A1(n1159), .A2(n1158), .ZN(n2493) );
  NAND2_X1 U1520 ( .A1(regfile_alu_wdata_fw_i[23]), .A2(n1193), .ZN(n1164) );
  INV_X1 U1521 ( .A(regfile_data_rc_id[23]), .ZN(n2339) );
  AOI22_X1 U1522 ( .A1(n1195), .A2(regfile_data_rb_id[23]), .B1(n1194), .B2(
        jump_target_o[23]), .ZN(n1161) );
  OAI21_X1 U1523 ( .B1(n1160), .B2(n2339), .A(n1161), .ZN(n1162) );
  AOI21_X1 U1524 ( .B1(regfile_wdata_wb_i[23]), .B2(n1198), .A(n1162), .ZN(
        n1163) );
  NAND2_X1 U1525 ( .A1(n1164), .A2(n1163), .ZN(n2494) );
  NAND2_X1 U1527 ( .A1(regfile_alu_wdata_fw_i[24]), .A2(n1193), .ZN(n1168) );
  INV_X1 U1528 ( .A(regfile_data_rc_id[24]), .ZN(n2348) );
  AOI22_X1 U1529 ( .A1(n1195), .A2(regfile_data_rb_id[24]), .B1(n1194), .B2(
        jump_target_o[24]), .ZN(n1165) );
  OAI21_X1 U1530 ( .B1(n1160), .B2(n2348), .A(n1165), .ZN(n1166) );
  AOI21_X1 U1531 ( .B1(regfile_wdata_wb_i[24]), .B2(n1198), .A(n1166), .ZN(
        n1167) );
  NAND2_X1 U1532 ( .A1(n1168), .A2(n1167), .ZN(n2495) );
  NAND2_X1 U1534 ( .A1(regfile_alu_wdata_fw_i[25]), .A2(n1193), .ZN(n1172) );
  INV_X1 U1535 ( .A(regfile_data_rc_id[25]), .ZN(n2357) );
  AOI22_X1 U1536 ( .A1(n1195), .A2(regfile_data_rb_id[25]), .B1(n1194), .B2(
        jump_target_o[25]), .ZN(n1169) );
  OAI21_X1 U1537 ( .B1(n1160), .B2(n2357), .A(n1169), .ZN(n1170) );
  AOI21_X1 U1538 ( .B1(regfile_wdata_wb_i[25]), .B2(n1198), .A(n1170), .ZN(
        n1171) );
  NAND2_X1 U1539 ( .A1(n1172), .A2(n1171), .ZN(n2496) );
  INV_X1 U1541 ( .A(regfile_alu_wdata_fw_i[26]), .ZN(n2372) );
  INV_X1 U1542 ( .A(n1193), .ZN(n1176) );
  INV_X1 U1543 ( .A(regfile_data_rc_id[26]), .ZN(n2366) );
  AOI22_X1 U1544 ( .A1(n1195), .A2(regfile_data_rb_id[26]), .B1(n1194), .B2(
        jump_target_o[26]), .ZN(n1173) );
  OAI21_X1 U1545 ( .B1(n1160), .B2(n2366), .A(n1173), .ZN(n1174) );
  AOI21_X1 U1546 ( .B1(regfile_wdata_wb_i[26]), .B2(n1198), .A(n1174), .ZN(
        n1175) );
  OAI21_X1 U1547 ( .B1(n2372), .B2(n1176), .A(n1175), .ZN(n2497) );
  NAND2_X1 U1549 ( .A1(regfile_alu_wdata_fw_i[27]), .A2(n1193), .ZN(n1180) );
  INV_X1 U1550 ( .A(regfile_data_rc_id[27]), .ZN(n2375) );
  AOI22_X1 U1551 ( .A1(n1195), .A2(regfile_data_rb_id[27]), .B1(n1194), .B2(
        jump_target_o[27]), .ZN(n1177) );
  OAI21_X1 U1552 ( .B1(n1160), .B2(n2375), .A(n1177), .ZN(n1178) );
  AOI21_X1 U1553 ( .B1(regfile_wdata_wb_i[27]), .B2(n1198), .A(n1178), .ZN(
        n1179) );
  NAND2_X1 U1554 ( .A1(n1180), .A2(n1179), .ZN(n2498) );
  NAND2_X1 U1556 ( .A1(regfile_alu_wdata_fw_i[28]), .A2(n1193), .ZN(n1184) );
  INV_X1 U1557 ( .A(regfile_data_rc_id[28]), .ZN(n2384) );
  AOI22_X1 U1558 ( .A1(n1195), .A2(regfile_data_rb_id[28]), .B1(n1194), .B2(
        jump_target_o[28]), .ZN(n1181) );
  OAI21_X1 U1559 ( .B1(n1160), .B2(n2384), .A(n1181), .ZN(n1182) );
  AOI21_X1 U1560 ( .B1(regfile_wdata_wb_i[28]), .B2(n1198), .A(n1182), .ZN(
        n1183) );
  NAND2_X1 U1561 ( .A1(n1184), .A2(n1183), .ZN(n2499) );
  NAND2_X1 U1563 ( .A1(regfile_alu_wdata_fw_i[29]), .A2(n1193), .ZN(n1188) );
  INV_X1 U1564 ( .A(regfile_data_rc_id[29]), .ZN(n2393) );
  AOI22_X1 U1565 ( .A1(n1195), .A2(regfile_data_rb_id[29]), .B1(n1194), .B2(
        jump_target_o[29]), .ZN(n1185) );
  OAI21_X1 U1566 ( .B1(n1160), .B2(n2393), .A(n1185), .ZN(n1186) );
  AOI21_X1 U1567 ( .B1(regfile_wdata_wb_i[29]), .B2(n1198), .A(n1186), .ZN(
        n1187) );
  NAND2_X1 U1568 ( .A1(n1188), .A2(n1187), .ZN(n2500) );
  NAND2_X1 U1570 ( .A1(regfile_alu_wdata_fw_i[30]), .A2(n1193), .ZN(n1192) );
  INV_X1 U1571 ( .A(regfile_data_rc_id[30]), .ZN(n2403) );
  AOI22_X1 U1572 ( .A1(n1195), .A2(regfile_data_rb_id[30]), .B1(n1194), .B2(
        jump_target_o[30]), .ZN(n1189) );
  OAI21_X1 U1573 ( .B1(n1160), .B2(n2403), .A(n1189), .ZN(n1190) );
  AOI21_X1 U1574 ( .B1(regfile_wdata_wb_i[30]), .B2(n1198), .A(n1190), .ZN(
        n1191) );
  NAND2_X1 U1575 ( .A1(n1192), .A2(n1191), .ZN(n2501) );
  NAND2_X1 U1577 ( .A1(regfile_alu_wdata_fw_i[31]), .A2(n1193), .ZN(n1200) );
  INV_X1 U1578 ( .A(regfile_data_rc_id[31]), .ZN(n2415) );
  AOI22_X1 U1579 ( .A1(n1195), .A2(regfile_data_rb_id[31]), .B1(n1194), .B2(
        jump_target_o[31]), .ZN(n1196) );
  OAI21_X1 U1580 ( .B1(n1160), .B2(n2415), .A(n1196), .ZN(n1197) );
  AOI21_X1 U1581 ( .B1(regfile_wdata_wb_i[31]), .B2(n1198), .A(n1197), .ZN(
        n1199) );
  NAND2_X1 U1582 ( .A1(n1200), .A2(n1199), .ZN(n2502) );
  NAND2_X1 U1584 ( .A1(regfile_alu_wdata_fw_i[0]), .A2(n1879), .ZN(n1203) );
  NAND2_X1 U1585 ( .A1(n1203), .A2(n175), .ZN(n2136) );
  NAND2_X1 U1586 ( .A1(alu_op_b_mux_sel[1]), .A2(alu_op_b_mux_sel[0]), .ZN(
        n1876) );
  NOR2_X1 U1587 ( .A1(n1876), .A2(alu_op_b_mux_sel[2]), .ZN(n1865) );
  NAND2_X1 U1588 ( .A1(n2136), .A2(n1865), .ZN(n1226) );
  INV_X1 U1589 ( .A(alu_op_b_mux_sel[1]), .ZN(n1204) );
  INV_X1 U1590 ( .A(alu_op_b_mux_sel[0]), .ZN(n1689) );
  AOI21_X1 U1591 ( .B1(n1204), .B2(n1689), .A(alu_op_b_mux_sel[2]), .ZN(n1684)
         );
  INV_X1 U1592 ( .A(n1684), .ZN(n1690) );
  OR2_X1 U1593 ( .A1(alu_op_b_mux_sel[1]), .A2(n1689), .ZN(n1679) );
  INV_X1 U1594 ( .A(n1679), .ZN(n1875) );
  NAND2_X1 U1595 ( .A1(n1875), .A2(n1853), .ZN(n1779) );
  INV_X1 U1596 ( .A(n1865), .ZN(n1798) );
  OR2_X1 U1597 ( .A1(n2130), .A2(n1798), .ZN(n1863) );
  INV_X1 U1598 ( .A(n1863), .ZN(n1734) );
  NAND2_X1 U1599 ( .A1(alu_op_b_mux_sel[1]), .A2(n1689), .ZN(n1901) );
  NOR2_X1 U1600 ( .A1(n1901), .A2(alu_op_b_mux_sel[2]), .ZN(n1714) );
  NOR2_X1 U1601 ( .A1(imm_b_mux_sel[1]), .A2(imm_b_mux_sel[2]), .ZN(n1212) );
  AND2_X1 U1602 ( .A1(imm_b_mux_sel[3]), .A2(n1212), .ZN(n1209) );
  AND2_X1 U1603 ( .A1(n1209), .A2(imm_b_mux_sel[0]), .ZN(n1898) );
  AND2_X1 U1604 ( .A1(n1714), .A2(n1898), .ZN(n1859) );
  INV_X1 U1605 ( .A(n1656), .ZN(n1633) );
  NAND2_X1 U1606 ( .A1(instr_rdata_i[20]), .A2(n1738), .ZN(n2064) );
  NOR2_X1 U1607 ( .A1(n1633), .A2(n2064), .ZN(n1208) );
  XNOR2_X1 U1608 ( .A(n1208), .B(n1207), .ZN(n1231) );
  NAND2_X1 U1609 ( .A1(n1859), .A2(n1231), .ZN(n1223) );
  INV_X1 U1610 ( .A(imm_b_mux_sel[0]), .ZN(n2109) );
  NAND2_X1 U1611 ( .A1(n2109), .A2(n1209), .ZN(n1210) );
  OR2_X1 U1612 ( .A1(n1901), .A2(n1210), .ZN(n1855) );
  NOR2_X1 U1613 ( .A1(alu_op_b_mux_sel[2]), .A2(n1855), .ZN(n1211) );
  NAND2_X1 U1614 ( .A1(instr_rdata_i[25]), .A2(n1211), .ZN(n1222) );
  NOR2_X1 U1615 ( .A1(imm_b_mux_sel[3]), .A2(imm_b_mux_sel[1]), .ZN(n1788) );
  INV_X1 U1616 ( .A(n1788), .ZN(n1214) );
  INV_X1 U1617 ( .A(n1212), .ZN(n1703) );
  NAND2_X1 U1618 ( .A1(imm_b_mux_sel[3]), .A2(n1703), .ZN(n1213) );
  OAI21_X1 U1619 ( .B1(imm_b_mux_sel[0]), .B2(n1214), .A(n1213), .ZN(n1671) );
  AND2_X1 U1620 ( .A1(n1671), .A2(instr_rdata_i[20]), .ZN(n1220) );
  INV_X1 U1621 ( .A(imm_b_mux_sel[2]), .ZN(n1890) );
  INV_X1 U1622 ( .A(imm_b_mux_sel[3]), .ZN(n2108) );
  OAI211_X1 U1623 ( .C1(imm_b_mux_sel[0]), .C2(imm_b_mux_sel[1]), .A(
        instr_rdata_i[25]), .B(n2108), .ZN(n1218) );
  NOR2_X1 U1624 ( .A1(imm_b_mux_sel[3]), .A2(n1703), .ZN(n1215) );
  AND2_X1 U1625 ( .A1(imm_b_mux_sel[0]), .A2(n1215), .ZN(n1670) );
  INV_X1 U1626 ( .A(n1670), .ZN(n1217) );
  OAI22_X1 U1627 ( .A1(n1890), .A2(n1218), .B1(n1217), .B2(n1216), .ZN(n1219)
         );
  OAI21_X1 U1628 ( .B1(n1220), .B2(n1219), .A(n1714), .ZN(n1221) );
  NAND3_X1 U1629 ( .A1(n1223), .A2(n1222), .A3(n1221), .ZN(n1224) );
  AOI21_X1 U1630 ( .B1(n1734), .B2(n114), .A(n1224), .ZN(n1225) );
  AOI22_X1 U1632 ( .A1(regfile_alu_wdata_fw_i[1]), .A2(n1228), .B1(n1227), 
        .B2(regfile_wdata_wb_i[1]), .ZN(n2143) );
  OR2_X1 U1633 ( .A1(n2143), .A2(n1779), .ZN(n1632) );
  NAND2_X1 U1634 ( .A1(n1229), .A2(n1690), .ZN(n1396) );
  NAND2_X1 U1635 ( .A1(n1230), .A2(n1865), .ZN(n1328) );
  NOR2_X1 U1636 ( .A1(n2140), .A2(n1779), .ZN(n1842) );
  AND2_X1 U1637 ( .A1(alu_vec_mode[1]), .A2(alu_vec_mode[0]), .ZN(n1732) );
  INV_X1 U1638 ( .A(n1732), .ZN(n2002) );
  NOR2_X1 U1639 ( .A1(n1855), .A2(n2002), .ZN(n1889) );
  NAND2_X1 U1640 ( .A1(n1889), .A2(n1853), .ZN(n1751) );
  NAND2_X1 U1641 ( .A1(instr_rdata_i[21]), .A2(n2467), .ZN(n2021) );
  NOR2_X1 U1642 ( .A1(n1633), .A2(n2021), .ZN(n1232) );
  XOR2_X1 U1643 ( .A(n1232), .B(n1231), .Z(n1240) );
  NAND2_X1 U1644 ( .A1(imm_b_mux_sel[1]), .A2(n2108), .ZN(n1713) );
  INV_X1 U1645 ( .A(n1713), .ZN(n1233) );
  AND2_X1 U1646 ( .A1(imm_b_mux_sel[2]), .A2(n1233), .ZN(n1705) );
  NAND2_X1 U1647 ( .A1(n1705), .A2(instr_rdata_i[20]), .ZN(n1238) );
  NAND2_X1 U1648 ( .A1(is_compressed_i), .A2(n2455), .ZN(n1640) );
  INV_X1 U1649 ( .A(n1640), .ZN(n1234) );
  NOR3_X1 U1650 ( .A1(imm_b_mux_sel[2]), .A2(n2109), .A3(n1713), .ZN(n1639) );
  NOR4_X1 U1651 ( .A1(imm_b_mux_sel[1]), .A2(imm_b_mux_sel[3]), .A3(n2109), 
        .A4(n1890), .ZN(n1669) );
  AOI22_X1 U1652 ( .A1(n1234), .A2(n1639), .B1(n1669), .B2(n2683), .ZN(n1237)
         );
  NAND2_X1 U1653 ( .A1(n1671), .A2(instr_rdata_i[21]), .ZN(n1236) );
  NAND2_X1 U1654 ( .A1(n1670), .A2(instr_rdata_i[8]), .ZN(n1235) );
  NAND4_X1 U1655 ( .A1(n1238), .A2(n1237), .A3(n1236), .A4(n1235), .ZN(n1239)
         );
  AOI22_X1 U1656 ( .A1(n1859), .A2(n1240), .B1(n1714), .B2(n1239), .ZN(n1241)
         );
  OAI21_X1 U1657 ( .B1(n2467), .B2(n1751), .A(n1241), .ZN(n1242) );
  AOI21_X1 U1658 ( .B1(n1842), .B2(regfile_data_rc_id[1]), .A(n1242), .ZN(
        n1243) );
  NAND4_X1 U1659 ( .A1(n1632), .A2(n1396), .A3(n1328), .A4(n1243), .ZN(n1874)
         );
  NAND2_X1 U1661 ( .A1(n1898), .A2(n1633), .ZN(n1644) );
  NAND2_X1 U1662 ( .A1(n1670), .A2(instr_rdata_i[9]), .ZN(n1643) );
  NAND2_X1 U1663 ( .A1(n1671), .A2(instr_rdata_i[22]), .ZN(n1642) );
  AOI22_X1 U1664 ( .A1(n1640), .A2(n1639), .B1(n1669), .B2(n2678), .ZN(n1641)
         );
  NAND4_X1 U1665 ( .A1(n1644), .A2(n1643), .A3(n1642), .A4(n1641), .ZN(n1645)
         );
  AOI21_X1 U1666 ( .B1(n1705), .B2(instr_rdata_i[21]), .A(n1645), .ZN(n1646)
         );
  OAI22_X1 U1667 ( .A1(n1647), .A2(n1679), .B1(n1646), .B2(n1901), .ZN(n1652)
         );
  AND2_X1 U1668 ( .A1(regfile_wdata_wb_i[2]), .A2(n2179), .ZN(n1648) );
  AOI21_X1 U1669 ( .B1(regfile_alu_wdata_fw_i[2]), .B2(n1879), .A(n1648), .ZN(
        n2150) );
  NAND2_X1 U1670 ( .A1(n1649), .A2(n2627), .ZN(n1650) );
  AOI21_X1 U1671 ( .B1(n2150), .B2(n1650), .A(n1876), .ZN(n1651) );
  OAI21_X1 U1672 ( .B1(n1652), .B2(n1651), .A(n1853), .ZN(n1653) );
  INV_X1 U1674 ( .A(n1901), .ZN(n1677) );
  NAND2_X1 U1675 ( .A1(n1705), .A2(instr_rdata_i[22]), .ZN(n1660) );
  AOI22_X1 U1676 ( .A1(n1670), .A2(instr_rdata_i[10]), .B1(n1669), .B2(n2668), 
        .ZN(n1659) );
  INV_X1 U1677 ( .A(n1655), .ZN(n2050) );
  NAND3_X1 U1678 ( .A1(instr_rdata_i[22]), .A2(n1904), .A3(n1991), .ZN(n1694)
         );
  NOR2_X1 U1679 ( .A1(n2050), .A2(n1694), .ZN(n1657) );
  NOR2_X1 U1680 ( .A1(n1657), .A2(n1656), .ZN(n1696) );
  AOI22_X1 U1681 ( .A1(n1696), .A2(n1898), .B1(n1671), .B2(instr_rdata_i[23]), 
        .ZN(n1658) );
  NAND3_X1 U1682 ( .A1(n1660), .A2(n1659), .A3(n1658), .ZN(n1661) );
  NAND2_X1 U1683 ( .A1(n1677), .A2(n1661), .ZN(n1662) );
  OAI21_X1 U1684 ( .B1(n1663), .B2(n1679), .A(n1662), .ZN(n1666) );
  NOR2_X1 U1685 ( .A1(n1664), .A2(n1876), .ZN(n1665) );
  OAI21_X1 U1686 ( .B1(n1666), .B2(n1665), .A(n1853), .ZN(n1668) );
  NAND2_X1 U1687 ( .A1(n1668), .A2(n1667), .ZN(n1925) );
  NAND2_X1 U1689 ( .A1(n1705), .A2(instr_rdata_i[23]), .ZN(n1675) );
  AOI22_X1 U1690 ( .A1(n1670), .A2(instr_rdata_i[11]), .B1(n1669), .B2(
        instr_rdata_i[29]), .ZN(n1674) );
  OR2_X1 U1691 ( .A1(n2064), .A2(n1694), .ZN(n1695) );
  XNOR2_X1 U1692 ( .A(n1696), .B(n1695), .ZN(n1672) );
  AOI22_X1 U1693 ( .A1(n1672), .A2(n1898), .B1(n1671), .B2(n2604), .ZN(n1673)
         );
  NAND3_X1 U1694 ( .A1(n1675), .A2(n1674), .A3(n1673), .ZN(n1676) );
  NAND2_X1 U1695 ( .A1(n1677), .A2(n1676), .ZN(n1678) );
  OAI21_X1 U1696 ( .B1(n1680), .B2(n1679), .A(n1678), .ZN(n1683) );
  NOR2_X1 U1697 ( .A1(n1681), .A2(n1876), .ZN(n1682) );
  OAI21_X1 U1698 ( .B1(n1683), .B2(n1682), .A(n1853), .ZN(n1687) );
  NAND2_X1 U1699 ( .A1(n1687), .A2(n1686), .ZN(n1940) );
  NAND2_X1 U1701 ( .A1(n1688), .A2(n1865), .ZN(n1712) );
  NAND2_X1 U1702 ( .A1(alu_op_b_mux_sel[2]), .A2(n1689), .ZN(n1691) );
  OAI21_X1 U1703 ( .B1(alu_op_b_mux_sel[1]), .B2(n1691), .A(n1690), .ZN(n1881)
         );
  NAND2_X1 U1704 ( .A1(n1692), .A2(n134), .ZN(n1711) );
  NAND2_X1 U1705 ( .A1(n1693), .A2(n131), .ZN(n1710) );
  NOR2_X1 U1706 ( .A1(n2021), .A2(n1694), .ZN(n1698) );
  NAND2_X1 U1707 ( .A1(n1696), .A2(n1695), .ZN(n1697) );
  XNOR2_X1 U1708 ( .A(n1698), .B(n1697), .ZN(n1699) );
  NAND2_X1 U1709 ( .A1(n1859), .A2(n1699), .ZN(n1708) );
  NAND2_X1 U1710 ( .A1(imm_b_mux_sel[3]), .A2(imm_b_mux_sel[1]), .ZN(n1700) );
  NOR2_X1 U1711 ( .A1(imm_b_mux_sel[0]), .A2(n1700), .ZN(n1787) );
  INV_X1 U1712 ( .A(n1787), .ZN(n1702) );
  NAND2_X1 U1713 ( .A1(imm_b_mux_sel[2]), .A2(imm_b_mux_sel[3]), .ZN(n1701) );
  OAI211_X1 U1714 ( .C1(imm_b_mux_sel[3]), .C2(n1703), .A(n1702), .B(n1701), 
        .ZN(n1704) );
  AND2_X1 U1715 ( .A1(n1714), .A2(n1704), .ZN(n1770) );
  NAND2_X1 U1716 ( .A1(n1770), .A2(instr_rdata_i[25]), .ZN(n1707) );
  NAND2_X1 U1717 ( .A1(n1714), .A2(n1890), .ZN(n1803) );
  NAND4_X1 U1718 ( .A1(imm_b_mux_sel[0]), .A2(imm_b_mux_sel[3]), .A3(
        imm_b_mux_sel[1]), .A4(n2604), .ZN(n1789) );
  OR2_X1 U1719 ( .A1(n1803), .A2(n1789), .ZN(n1716) );
  NAND3_X1 U1720 ( .A1(n1714), .A2(n1705), .A3(n2604), .ZN(n1706) );
  AND4_X1 U1721 ( .A1(n1708), .A2(n1707), .A3(n1716), .A4(n1706), .ZN(n1709)
         );
  NOR2_X1 U1724 ( .A1(imm_b_mux_sel[0]), .A2(n1713), .ZN(n1892) );
  AND2_X1 U1725 ( .A1(n2604), .A2(n1892), .ZN(n1791) );
  NAND3_X1 U1726 ( .A1(n1714), .A2(imm_b_mux_sel[2]), .A3(n1791), .ZN(n1715)
         );
  AND2_X1 U1727 ( .A1(n1716), .A2(n1715), .ZN(n1772) );
  AOI22_X1 U1728 ( .A1(n1770), .A2(n2683), .B1(n1859), .B2(n1723), .ZN(n1717)
         );
  OAI211_X1 U1729 ( .C1(n1863), .C2(n1718), .A(n1772), .B(n1717), .ZN(n1719)
         );
  NAND2_X1 U1732 ( .A1(n1879), .A2(n1865), .ZN(n1721) );
  OAI21_X1 U1733 ( .B1(n2185), .B2(n1779), .A(n1721), .ZN(n1763) );
  NAND2_X1 U1734 ( .A1(n2179), .A2(n1865), .ZN(n1722) );
  OAI21_X1 U1735 ( .B1(n2178), .B2(n1779), .A(n1722), .ZN(n1766) );
  INV_X1 U1736 ( .A(n1766), .ZN(n1741) );
  NAND3_X1 U1737 ( .A1(instr_rdata_i[23]), .A2(n1984), .A3(n1904), .ZN(n1768)
         );
  NOR2_X1 U1738 ( .A1(n2050), .A2(n1768), .ZN(n1725) );
  INV_X1 U1739 ( .A(n1723), .ZN(n1724) );
  XNOR2_X1 U1740 ( .A(n1725), .B(n1724), .ZN(n1746) );
  AOI22_X1 U1741 ( .A1(n2678), .A2(n1770), .B1(n1859), .B2(n1746), .ZN(n1726)
         );
  OAI211_X1 U1742 ( .C1(n1863), .C2(n1727), .A(n1772), .B(n1726), .ZN(n1728)
         );
  AOI21_X1 U1743 ( .B1(n1842), .B2(regfile_data_rc_id[7]), .A(n1728), .ZN(
        n1729) );
  OAI21_X1 U1744 ( .B1(n2182), .B2(n1741), .A(n1729), .ZN(n1730) );
  AOI21_X1 U1745 ( .B1(regfile_alu_wdata_fw_i[7]), .B2(n1763), .A(n1730), .ZN(
        n1731) );
  NAND2_X1 U1747 ( .A1(n1872), .A2(n1848), .ZN(n2013) );
  INV_X1 U1748 ( .A(n1772), .ZN(n1733) );
  AOI21_X1 U1749 ( .B1(n1734), .B2(n24), .A(n1733), .ZN(n1737) );
  OR2_X1 U1750 ( .A1(n2064), .A2(n1768), .ZN(n1745) );
  XNOR2_X1 U1751 ( .A(n1746), .B(n1745), .ZN(n1735) );
  AOI22_X1 U1752 ( .A1(n1770), .A2(n2668), .B1(n1859), .B2(n1735), .ZN(n1736)
         );
  OAI211_X1 U1753 ( .C1(n1738), .C2(n1751), .A(n1737), .B(n1736), .ZN(n1739)
         );
  AOI21_X1 U1754 ( .B1(n1842), .B2(regfile_data_rc_id[8]), .A(n1739), .ZN(
        n1740) );
  OAI21_X1 U1755 ( .B1(n2195), .B2(n1741), .A(n1740), .ZN(n1742) );
  AOI21_X1 U1756 ( .B1(regfile_alu_wdata_fw_i[8]), .B2(n1763), .A(n1742), .ZN(
        n1743) );
  OAI21_X1 U1757 ( .B1(n2198), .B2(n1881), .A(n1743), .ZN(n2012) );
  INV_X1 U1758 ( .A(n1848), .ZN(n2035) );
  NAND2_X1 U1759 ( .A1(n2012), .A2(n2035), .ZN(n1744) );
  NAND2_X1 U1760 ( .A1(n2013), .A2(n1744), .ZN(n2507) );
  NAND2_X1 U1762 ( .A1(regfile_wdata_wb_i[9]), .A2(n1766), .ZN(n1757) );
  NOR2_X1 U1763 ( .A1(n2021), .A2(n1768), .ZN(n1748) );
  NAND2_X1 U1764 ( .A1(n1746), .A2(n1745), .ZN(n1747) );
  XNOR2_X1 U1765 ( .A(n1748), .B(n1747), .ZN(n1784) );
  NAND2_X1 U1766 ( .A1(n1859), .A2(n1784), .ZN(n1750) );
  NAND2_X1 U1767 ( .A1(n1770), .A2(instr_rdata_i[29]), .ZN(n1749) );
  OAI211_X1 U1768 ( .C1(n1751), .C2(n1984), .A(n1750), .B(n1749), .ZN(n1752)
         );
  INV_X1 U1769 ( .A(n1752), .ZN(n1753) );
  OAI211_X1 U1770 ( .C1(n1863), .C2(n1754), .A(n1753), .B(n1772), .ZN(n1755)
         );
  AOI21_X1 U1771 ( .B1(n1842), .B2(regfile_data_rc_id[9]), .A(n1755), .ZN(
        n1756) );
  NAND2_X1 U1772 ( .A1(n1757), .A2(n1756), .ZN(n1758) );
  AOI21_X1 U1773 ( .B1(regfile_alu_wdata_fw_i[9]), .B2(n1763), .A(n1758), .ZN(
        n1759) );
  OAI21_X1 U1774 ( .B1(n2204), .B2(n1881), .A(n1759), .ZN(n2014) );
  OR2_X1 U1775 ( .A1(n2014), .A2(n1848), .ZN(n1760) );
  OAI21_X1 U1776 ( .B1(n1874), .B2(n2035), .A(n1760), .ZN(n2508) );
  NAND2_X1 U1779 ( .A1(n1912), .A2(n1848), .ZN(n2048) );
  NOR2_X1 U1780 ( .A1(n1882), .A2(n1881), .ZN(n1762) );
  OR2_X1 U1781 ( .A1(n1763), .A2(n1762), .ZN(n1847) );
  NOR2_X1 U1782 ( .A1(n1764), .A2(n1881), .ZN(n1765) );
  NOR2_X1 U1783 ( .A1(n1766), .A2(n1765), .ZN(n1845) );
  INV_X1 U1784 ( .A(n2209), .ZN(n1767) );
  NOR2_X1 U1785 ( .A1(n1767), .A2(n1881), .ZN(n1886) );
  NAND2_X1 U1786 ( .A1(instr_rdata_i[21]), .A2(instr_rdata_i[20]), .ZN(n2083)
         );
  OR2_X1 U1787 ( .A1(n2083), .A2(n1768), .ZN(n1783) );
  XNOR2_X1 U1788 ( .A(n1784), .B(n1783), .ZN(n1769) );
  AOI22_X1 U1789 ( .A1(n1770), .A2(instr_rdata_i[30]), .B1(n1859), .B2(n1769), 
        .ZN(n1771) );
  OAI211_X1 U1790 ( .C1(n1863), .C2(n1773), .A(n1772), .B(n1771), .ZN(n1774)
         );
  AOI21_X1 U1791 ( .B1(n1886), .B2(regfile_data_rb_id[10]), .A(n1774), .ZN(
        n1776) );
  NAND2_X1 U1792 ( .A1(regfile_data_rc_id[10]), .A2(n1842), .ZN(n1775) );
  OAI211_X1 U1793 ( .C1(n2215), .C2(n1845), .A(n1776), .B(n1775), .ZN(n1777)
         );
  AOI21_X1 U1794 ( .B1(regfile_alu_wdata_fw_i[10]), .B2(n1847), .A(n1777), 
        .ZN(n2045) );
  NAND2_X1 U1795 ( .A1(n2048), .A2(n182), .ZN(n2509) );
  OAI22_X1 U1797 ( .A1(n1780), .A2(n1779), .B1(n1778), .B2(n1881), .ZN(n1800)
         );
  NOR2_X1 U1798 ( .A1(n1781), .A2(n1884), .ZN(n1782) );
  AOI21_X1 U1799 ( .B1(regfile_alu_wdata_fw_i[11]), .B2(n1879), .A(n1782), 
        .ZN(n2224) );
  NAND3_X1 U1800 ( .A1(instr_rdata_i[22]), .A2(instr_rdata_i[23]), .A3(n1904), 
        .ZN(n1824) );
  NOR2_X1 U1801 ( .A1(n2050), .A2(n1824), .ZN(n1786) );
  NAND2_X1 U1802 ( .A1(n1784), .A2(n1783), .ZN(n1785) );
  XNOR2_X1 U1803 ( .A(n1786), .B(n1785), .ZN(n1813) );
  OAI21_X1 U1804 ( .B1(n1788), .B2(n1787), .A(instr_rdata_i[31]), .ZN(n1790)
         );
  NAND3_X1 U1805 ( .A1(n1890), .A2(n1790), .A3(n1789), .ZN(n1794) );
  AOI21_X1 U1806 ( .B1(imm_b_mux_sel[3]), .B2(instr_rdata_i[31]), .A(n1791), 
        .ZN(n1792) );
  NAND2_X1 U1807 ( .A1(imm_b_mux_sel[2]), .A2(n1792), .ZN(n1793) );
  NAND2_X1 U1808 ( .A1(n1794), .A2(n1793), .ZN(n1795) );
  NOR2_X1 U1809 ( .A1(n1901), .A2(n1795), .ZN(n1893) );
  AND2_X1 U1810 ( .A1(n1893), .A2(n1853), .ZN(n1856) );
  AOI211_X1 U1811 ( .C1(n1859), .C2(n1813), .A(n1856), .B(n1796), .ZN(n1797)
         );
  OAI21_X1 U1812 ( .B1(n2224), .B2(n1798), .A(n1797), .ZN(n1799) );
  NOR2_X1 U1813 ( .A1(n1800), .A2(n1799), .ZN(n2059) );
  NAND2_X1 U1815 ( .A1(n1940), .A2(n1848), .ZN(n2078) );
  INV_X1 U1816 ( .A(n1845), .ZN(n1823) );
  NAND2_X1 U1817 ( .A1(regfile_wdata_wb_i[12]), .A2(n1823), .ZN(n1810) );
  OR2_X1 U1818 ( .A1(n2064), .A2(n1824), .ZN(n1812) );
  XNOR2_X1 U1819 ( .A(n1813), .B(n1812), .ZN(n1801) );
  AOI21_X1 U1820 ( .B1(n1859), .B2(n1801), .A(n1856), .ZN(n1805) );
  INV_X1 U1821 ( .A(n1892), .ZN(n1802) );
  NOR2_X1 U1822 ( .A1(n1803), .A2(n1802), .ZN(n1860) );
  NAND2_X1 U1823 ( .A1(n1860), .A2(instr_rdata_i[12]), .ZN(n1804) );
  OAI211_X1 U1824 ( .C1(n1863), .C2(n1806), .A(n1805), .B(n1804), .ZN(n1807)
         );
  AOI21_X1 U1825 ( .B1(n1886), .B2(regfile_data_rb_id[12]), .A(n1807), .ZN(
        n1809) );
  NAND2_X1 U1826 ( .A1(regfile_data_rc_id[12]), .A2(n1842), .ZN(n1808) );
  NAND3_X1 U1827 ( .A1(n1810), .A2(n1809), .A3(n1808), .ZN(n1811) );
  AOI21_X1 U1828 ( .B1(regfile_alu_wdata_fw_i[12]), .B2(n1847), .A(n1811), 
        .ZN(n2063) );
  NAND2_X1 U1829 ( .A1(n2078), .A2(n181), .ZN(n2511) );
  NAND2_X1 U1831 ( .A1(regfile_wdata_wb_i[13]), .A2(n1823), .ZN(n1820) );
  NOR2_X1 U1832 ( .A1(n2021), .A2(n1824), .ZN(n1815) );
  NAND2_X1 U1833 ( .A1(n1813), .A2(n1812), .ZN(n1814) );
  XNOR2_X1 U1834 ( .A(n1815), .B(n1814), .ZN(n1835) );
  AOI21_X1 U1835 ( .B1(n1859), .B2(n1835), .A(n1856), .ZN(n1816) );
  AOI21_X1 U1836 ( .B1(n1886), .B2(regfile_data_rb_id[13]), .A(n1817), .ZN(
        n1819) );
  NAND2_X1 U1837 ( .A1(regfile_data_rc_id[13]), .A2(n1842), .ZN(n1818) );
  NAND3_X1 U1838 ( .A1(n1820), .A2(n1819), .A3(n1818), .ZN(n1821) );
  AOI21_X1 U1839 ( .B1(regfile_alu_wdata_fw_i[13]), .B2(n1847), .A(n1821), 
        .ZN(n2092) );
  OR2_X1 U1841 ( .A1(n1822), .A2(n2035), .ZN(n2107) );
  NAND2_X1 U1842 ( .A1(regfile_wdata_wb_i[14]), .A2(n1823), .ZN(n1832) );
  OR2_X1 U1843 ( .A1(n2083), .A2(n1824), .ZN(n1834) );
  XNOR2_X1 U1844 ( .A(n1835), .B(n1834), .ZN(n1825) );
  AOI21_X1 U1845 ( .B1(n1859), .B2(n1825), .A(n1856), .ZN(n1827) );
  NAND2_X1 U1846 ( .A1(n1860), .A2(instr_rdata_i[14]), .ZN(n1826) );
  OAI211_X1 U1847 ( .C1(n1863), .C2(n1828), .A(n1827), .B(n1826), .ZN(n1829)
         );
  AOI21_X1 U1848 ( .B1(n1886), .B2(regfile_data_rb_id[14]), .A(n1829), .ZN(
        n1831) );
  NAND2_X1 U1849 ( .A1(regfile_data_rc_id[14]), .A2(n1842), .ZN(n1830) );
  NAND3_X1 U1850 ( .A1(n1832), .A2(n1831), .A3(n1830), .ZN(n1833) );
  AOI21_X1 U1851 ( .B1(regfile_alu_wdata_fw_i[14]), .B2(n1847), .A(n1833), 
        .ZN(n2106) );
  NAND2_X1 U1852 ( .A1(n2107), .A2(n183), .ZN(n2513) );
  INV_X1 U1854 ( .A(regfile_wdata_wb_i[15]), .ZN(n2262) );
  NAND3_X1 U1855 ( .A1(n2604), .A2(n1984), .A3(n1991), .ZN(n1913) );
  NOR2_X1 U1856 ( .A1(n2050), .A2(n1913), .ZN(n1837) );
  NAND2_X1 U1857 ( .A1(n1835), .A2(n1834), .ZN(n1836) );
  XNOR2_X1 U1858 ( .A(n1837), .B(n1836), .ZN(n1895) );
  AOI21_X1 U1859 ( .B1(n1859), .B2(n1895), .A(n1856), .ZN(n1839) );
  NAND2_X1 U1860 ( .A1(n1860), .A2(n113), .ZN(n1838) );
  OAI211_X1 U1861 ( .C1(n1863), .C2(n1840), .A(n1839), .B(n1838), .ZN(n1841)
         );
  AOI21_X1 U1862 ( .B1(n1886), .B2(regfile_data_rb_id[15]), .A(n1841), .ZN(
        n1844) );
  NAND2_X1 U1863 ( .A1(regfile_data_rc_id[15]), .A2(n1842), .ZN(n1843) );
  OAI211_X1 U1864 ( .C1(n2262), .C2(n1845), .A(n1844), .B(n1843), .ZN(n1846)
         );
  AOI21_X1 U1865 ( .B1(n2663), .B2(n1847), .A(n1846), .ZN(n2126) );
  NAND2_X1 U1866 ( .A1(n2506), .A2(n1848), .ZN(n2124) );
  INV_X1 U1868 ( .A(scalar_replication), .ZN(n1983) );
  NAND2_X1 U1869 ( .A1(regfile_alu_wdata_fw_i[16]), .A2(n1879), .ZN(n1851) );
  NAND2_X1 U1870 ( .A1(n1851), .A2(n1850), .ZN(n2271) );
  OR2_X1 U1871 ( .A1(n2064), .A2(n1913), .ZN(n1894) );
  XNOR2_X1 U1872 ( .A(n1895), .B(n1894), .ZN(n1858) );
  NAND2_X1 U1873 ( .A1(n2002), .A2(n2467), .ZN(n1852) );
  OAI211_X1 U1874 ( .C1(instr_rdata_i[23]), .C2(n2002), .A(n1853), .B(n1852), 
        .ZN(n1854) );
  OAI21_X1 U1875 ( .B1(n1855), .B2(n1854), .A(n1983), .ZN(n1857) );
  AOI211_X1 U1876 ( .C1(n1859), .C2(n1858), .A(n1857), .B(n1856), .ZN(n1862)
         );
  NAND2_X1 U1877 ( .A1(n1860), .A2(n80), .ZN(n1861) );
  OAI211_X1 U1878 ( .C1(n2274), .C2(n1863), .A(n1862), .B(n1861), .ZN(n1864)
         );
  AOI21_X1 U1879 ( .B1(n2271), .B2(n1865), .A(n1864), .ZN(n1870) );
  NAND2_X1 U1880 ( .A1(n1866), .A2(n134), .ZN(n1869) );
  NAND2_X1 U1881 ( .A1(n1867), .A2(n131), .ZN(n1868) );
  NAND3_X1 U1882 ( .A1(n1870), .A2(n1869), .A3(n1868), .ZN(n1871) );
  OAI21_X1 U1883 ( .B1(n1872), .B2(n1983), .A(n1871), .ZN(n2515) );
  NOR2_X1 U1887 ( .A1(scalar_replication), .A2(alu_op_b_mux_sel[2]), .ZN(n1899) );
  NAND2_X1 U1888 ( .A1(n1875), .A2(n1899), .ZN(n1907) );
  INV_X1 U1889 ( .A(n1876), .ZN(n1877) );
  NAND2_X1 U1890 ( .A1(n1877), .A2(n1899), .ZN(n1887) );
  INV_X1 U1891 ( .A(n1887), .ZN(n1878) );
  NAND2_X1 U1892 ( .A1(n1879), .A2(n1878), .ZN(n1880) );
  OAI21_X1 U1893 ( .B1(n2185), .B2(n1907), .A(n1880), .ZN(n1966) );
  NOR2_X1 U1894 ( .A1(n1881), .A2(scalar_replication), .ZN(n1885) );
  INV_X1 U1895 ( .A(n1885), .ZN(n1968) );
  NOR2_X1 U1896 ( .A1(n1882), .A2(n1968), .ZN(n1883) );
  OR2_X1 U1897 ( .A1(n1966), .A2(n1883), .ZN(n2122) );
  OR2_X1 U1898 ( .A1(n2178), .A2(n1907), .ZN(n1998) );
  NOR2_X1 U1899 ( .A1(n1884), .A2(n1887), .ZN(n1951) );
  AOI21_X1 U1900 ( .B1(n2207), .B2(n1885), .A(n1951), .ZN(n1926) );
  AND2_X1 U1901 ( .A1(n1998), .A2(n1926), .ZN(n2120) );
  AND2_X1 U1902 ( .A1(n1886), .A2(n1983), .ZN(n2116) );
  OR2_X1 U1903 ( .A1(n2130), .A2(n1887), .ZN(n2114) );
  NOR2_X1 U1904 ( .A1(n2114), .A2(n1888), .ZN(n1906) );
  NAND2_X1 U1905 ( .A1(n1889), .A2(n1899), .ZN(n2018) );
  NAND2_X1 U1906 ( .A1(n1890), .A2(n1899), .ZN(n1891) );
  NOR2_X1 U1907 ( .A1(n1901), .A2(n1891), .ZN(n2110) );
  AND2_X1 U1908 ( .A1(n2110), .A2(n1892), .ZN(n2096) );
  AND2_X1 U1909 ( .A1(n1893), .A2(n1899), .ZN(n2095) );
  AOI21_X1 U1910 ( .B1(n2096), .B2(n110), .A(n2095), .ZN(n1903) );
  NOR2_X1 U1911 ( .A1(n2021), .A2(n1913), .ZN(n1897) );
  NAND2_X1 U1912 ( .A1(n1895), .A2(n1894), .ZN(n1896) );
  XNOR2_X1 U1913 ( .A(n1897), .B(n1896), .ZN(n1928) );
  NAND2_X1 U1914 ( .A1(n1899), .A2(n1898), .ZN(n1900) );
  NAND2_X1 U1915 ( .A1(n1928), .A2(n2084), .ZN(n1902) );
  OAI211_X1 U1916 ( .C1(n2018), .C2(n1904), .A(n1903), .B(n1902), .ZN(n1905)
         );
  AOI211_X1 U1917 ( .C1(n2116), .C2(regfile_data_rb_id[17]), .A(n1906), .B(
        n1905), .ZN(n1909) );
  NOR2_X1 U1918 ( .A1(n2140), .A2(n1907), .ZN(n2117) );
  NAND2_X1 U1919 ( .A1(n2117), .A2(regfile_data_rc_id[17]), .ZN(n1908) );
  OAI211_X1 U1920 ( .C1(n2285), .C2(n2120), .A(n1909), .B(n1908), .ZN(n1910)
         );
  AOI21_X1 U1921 ( .B1(regfile_alu_wdata_fw_i[17]), .B2(n2122), .A(n1910), 
        .ZN(n1911) );
  OAI21_X1 U1922 ( .B1(n2665), .B2(n1983), .A(n1911), .ZN(n2517) );
  NAND2_X1 U1924 ( .A1(n2116), .A2(regfile_data_rb_id[18]), .ZN(n1918) );
  OR2_X1 U1925 ( .A1(n2083), .A2(n1913), .ZN(n1927) );
  XNOR2_X1 U1926 ( .A(n1928), .B(n1927), .ZN(n1916) );
  INV_X1 U1927 ( .A(n2096), .ZN(n1990) );
  NOR2_X1 U1928 ( .A1(n1990), .A2(n1914), .ZN(n1915) );
  AOI211_X1 U1929 ( .C1(n2084), .C2(n1916), .A(n2095), .B(n1915), .ZN(n1917)
         );
  OAI211_X1 U1930 ( .C1(n2114), .C2(n1919), .A(n1918), .B(n1917), .ZN(n1921)
         );
  NOR2_X1 U1931 ( .A1(n2294), .A2(n1926), .ZN(n1920) );
  AOI211_X1 U1932 ( .C1(n2117), .C2(regfile_data_rc_id[18]), .A(n1921), .B(
        n1920), .ZN(n1924) );
  NAND2_X1 U1933 ( .A1(regfile_alu_wdata_fw_i[18]), .A2(n2122), .ZN(n1923) );
  INV_X1 U1934 ( .A(n1998), .ZN(n1952) );
  NAND2_X1 U1935 ( .A1(regfile_wdata_wb_i[18]), .A2(n1952), .ZN(n1922) );
  INV_X1 U1937 ( .A(n1926), .ZN(n1996) );
  INV_X1 U1938 ( .A(n2117), .ZN(n2029) );
  NAND3_X1 U1939 ( .A1(n2604), .A2(instr_rdata_i[22]), .A3(n1991), .ZN(n1973)
         );
  NOR2_X1 U1940 ( .A1(n2050), .A2(n1973), .ZN(n1930) );
  NAND2_X1 U1941 ( .A1(n1928), .A2(n1927), .ZN(n1929) );
  XNOR2_X1 U1942 ( .A(n1930), .B(n1929), .ZN(n1954) );
  NAND2_X1 U1943 ( .A1(n1954), .A2(n2084), .ZN(n1932) );
  AOI21_X1 U1944 ( .B1(n2096), .B2(n116), .A(n2095), .ZN(n1931) );
  OAI211_X1 U1945 ( .C1(n2114), .C2(n1933), .A(n1932), .B(n1931), .ZN(n1934)
         );
  AOI21_X1 U1946 ( .B1(n2116), .B2(regfile_data_rb_id[19]), .A(n1934), .ZN(
        n1935) );
  OAI21_X1 U1947 ( .B1(n2029), .B2(n2303), .A(n1935), .ZN(n1936) );
  AOI21_X1 U1948 ( .B1(regfile_wdata_wb_i[19]), .B2(n1996), .A(n1936), .ZN(
        n1939) );
  NAND2_X1 U1949 ( .A1(regfile_alu_wdata_fw_i[19]), .A2(n2122), .ZN(n1938) );
  NAND2_X1 U1950 ( .A1(regfile_wdata_wb_i[19]), .A2(n1952), .ZN(n1937) );
  NAND2_X1 U1952 ( .A1(n1940), .A2(scalar_replication), .ZN(n1950) );
  NAND2_X1 U1953 ( .A1(regfile_alu_wdata_fw_i[20]), .A2(n2122), .ZN(n1949) );
  OR2_X1 U1954 ( .A1(n2064), .A2(n1973), .ZN(n1953) );
  XNOR2_X1 U1955 ( .A(n1954), .B(n1953), .ZN(n1943) );
  INV_X1 U1956 ( .A(n2114), .ZN(n2015) );
  NAND2_X1 U1957 ( .A1(n2015), .A2(regfile_data_ra_id[20]), .ZN(n1941) );
  INV_X1 U1958 ( .A(n2095), .ZN(n2112) );
  OAI211_X1 U1959 ( .C1(n1990), .C2(n2467), .A(n1941), .B(n2112), .ZN(n1942)
         );
  AOI21_X1 U1960 ( .B1(n2084), .B2(n1943), .A(n1942), .ZN(n1945) );
  NAND2_X1 U1961 ( .A1(n2116), .A2(regfile_data_rb_id[20]), .ZN(n1944) );
  OAI211_X1 U1962 ( .C1(n2029), .C2(n2312), .A(n1945), .B(n1944), .ZN(n1946)
         );
  AOI21_X1 U1963 ( .B1(regfile_wdata_wb_i[20]), .B2(n1996), .A(n1946), .ZN(
        n1948) );
  NAND2_X1 U1964 ( .A1(regfile_wdata_wb_i[20]), .A2(n1952), .ZN(n1947) );
  NAND3_X1 U1965 ( .A1(n1950), .A2(n1949), .A3(n180), .ZN(n2520) );
  AOI22_X1 U1967 ( .A1(regfile_alu_wdata_fw_i[21]), .A2(n2205), .B1(n2207), 
        .B2(regfile_wdata_wb_i[21]), .ZN(n1969) );
  OAI21_X1 U1968 ( .B1(n1952), .B2(n1951), .A(regfile_wdata_wb_i[21]), .ZN(
        n1964) );
  NAND2_X1 U1969 ( .A1(n2116), .A2(regfile_data_rb_id[21]), .ZN(n1961) );
  NOR2_X1 U1970 ( .A1(n2021), .A2(n1973), .ZN(n1956) );
  NAND2_X1 U1971 ( .A1(n1954), .A2(n1953), .ZN(n1955) );
  XNOR2_X1 U1972 ( .A(n1956), .B(n1955), .ZN(n1986) );
  AOI21_X1 U1973 ( .B1(instr_rdata_i[21]), .B2(n2096), .A(n2095), .ZN(n1957)
         );
  OAI21_X1 U1974 ( .B1(n2114), .B2(n1958), .A(n1957), .ZN(n1959) );
  AOI21_X1 U1975 ( .B1(n1986), .B2(n2084), .A(n1959), .ZN(n1960) );
  NAND2_X1 U1976 ( .A1(n1961), .A2(n1960), .ZN(n1962) );
  AOI21_X1 U1977 ( .B1(n2117), .B2(regfile_data_rc_id[21]), .A(n1962), .ZN(
        n1963) );
  NAND2_X1 U1978 ( .A1(n1964), .A2(n1963), .ZN(n1965) );
  AOI21_X1 U1979 ( .B1(regfile_alu_wdata_fw_i[21]), .B2(n1966), .A(n1965), 
        .ZN(n1967) );
  OAI21_X1 U1980 ( .B1(n1969), .B2(n1968), .A(n1967), .ZN(n1970) );
  AOI21_X1 U1981 ( .B1(n2662), .B2(scalar_replication), .A(n1970), .ZN(n2521)
         );
  OR2_X1 U1983 ( .A1(n2083), .A2(n1973), .ZN(n1985) );
  XNOR2_X1 U1984 ( .A(n1986), .B(n1985), .ZN(n1976) );
  NAND2_X1 U1985 ( .A1(n2015), .A2(regfile_data_ra_id[22]), .ZN(n1974) );
  OAI211_X1 U1986 ( .C1(n1984), .C2(n1990), .A(n1974), .B(n2112), .ZN(n1975)
         );
  AOI21_X1 U1987 ( .B1(n1976), .B2(n2084), .A(n1975), .ZN(n1978) );
  NAND2_X1 U1988 ( .A1(n2116), .A2(regfile_data_rb_id[22]), .ZN(n1977) );
  OAI211_X1 U1989 ( .C1(n2029), .C2(n2330), .A(n1978), .B(n1977), .ZN(n1979)
         );
  AOI21_X1 U1990 ( .B1(regfile_wdata_wb_i[22]), .B2(n1996), .A(n1979), .ZN(
        n1980) );
  OAI21_X1 U1991 ( .B1(n2333), .B2(n1998), .A(n1980), .ZN(n1981) );
  AOI21_X1 U1992 ( .B1(regfile_alu_wdata_fw_i[22]), .B2(n2122), .A(n1981), 
        .ZN(n1982) );
  OAI21_X1 U1993 ( .B1(n1822), .B2(n1983), .A(n1982), .ZN(n2523) );
  NAND2_X1 U1995 ( .A1(n2506), .A2(scalar_replication), .ZN(n2001) );
  NAND3_X1 U1996 ( .A1(n2604), .A2(instr_rdata_i[23]), .A3(n1984), .ZN(n2020)
         );
  NOR2_X1 U1997 ( .A1(n2050), .A2(n2020), .ZN(n1988) );
  NAND2_X1 U1998 ( .A1(n1986), .A2(n1985), .ZN(n1987) );
  XNOR2_X1 U1999 ( .A(n1988), .B(n1987), .ZN(n2023) );
  NAND2_X1 U2000 ( .A1(n2015), .A2(regfile_data_ra_id[23]), .ZN(n1989) );
  OAI211_X1 U2001 ( .C1(n1991), .C2(n1990), .A(n1989), .B(n2112), .ZN(n1992)
         );
  AOI21_X1 U2002 ( .B1(n2023), .B2(n2084), .A(n1992), .ZN(n1994) );
  NAND2_X1 U2003 ( .A1(n2116), .A2(regfile_data_rb_id[23]), .ZN(n1993) );
  OAI211_X1 U2004 ( .C1(n2029), .C2(n2339), .A(n1994), .B(n1993), .ZN(n1995)
         );
  AOI21_X1 U2005 ( .B1(regfile_wdata_wb_i[23]), .B2(n1996), .A(n1995), .ZN(
        n1997) );
  OAI21_X1 U2006 ( .B1(n1998), .B2(n2342), .A(n1997), .ZN(n1999) );
  AOI21_X1 U2007 ( .B1(regfile_alu_wdata_fw_i[23]), .B2(n2122), .A(n1999), 
        .ZN(n2000) );
  NAND2_X1 U2008 ( .A1(n2001), .A2(n2000), .ZN(n2524) );
  NAND2_X1 U2010 ( .A1(scalar_replication), .A2(n2002), .ZN(n2125) );
  INV_X1 U2011 ( .A(n2125), .ZN(n2033) );
  NAND2_X1 U2012 ( .A1(regfile_alu_wdata_fw_i[24]), .A2(n2122), .ZN(n2011) );
  INV_X1 U2013 ( .A(n2120), .ZN(n2100) );
  NAND2_X1 U2014 ( .A1(n2015), .A2(regfile_data_ra_id[24]), .ZN(n2004) );
  AOI21_X1 U2015 ( .B1(n2604), .B2(n2096), .A(n2095), .ZN(n2003) );
  OAI211_X1 U2016 ( .C1(n2018), .C2(n2429), .A(n2004), .B(n2003), .ZN(n2005)
         );
  AOI21_X1 U2017 ( .B1(n2116), .B2(regfile_data_rb_id[24]), .A(n2005), .ZN(
        n2008) );
  OR2_X1 U2018 ( .A1(n2064), .A2(n2020), .ZN(n2022) );
  XNOR2_X1 U2019 ( .A(n2023), .B(n2022), .ZN(n2006) );
  NAND2_X1 U2020 ( .A1(n2006), .A2(n2084), .ZN(n2007) );
  OAI211_X1 U2021 ( .C1(n2029), .C2(n2348), .A(n2008), .B(n2007), .ZN(n2009)
         );
  AOI21_X1 U2022 ( .B1(regfile_wdata_wb_i[24]), .B2(n2100), .A(n2009), .ZN(
        n2010) );
  NAND2_X1 U2024 ( .A1(regfile_alu_wdata_fw_i[25]), .A2(n2122), .ZN(n2032) );
  NAND2_X1 U2025 ( .A1(n2015), .A2(regfile_data_ra_id[25]), .ZN(n2017) );
  AOI21_X1 U2026 ( .B1(n2096), .B2(instr_rdata_i[25]), .A(n2095), .ZN(n2016)
         );
  OAI211_X1 U2027 ( .C1(n2018), .C2(n2430), .A(n2017), .B(n2016), .ZN(n2019)
         );
  AOI21_X1 U2028 ( .B1(n2116), .B2(regfile_data_rb_id[25]), .A(n2019), .ZN(
        n2028) );
  NOR2_X1 U2029 ( .A1(n2021), .A2(n2020), .ZN(n2025) );
  NAND2_X1 U2030 ( .A1(n2023), .A2(n2022), .ZN(n2024) );
  XNOR2_X1 U2031 ( .A(n2025), .B(n2024), .ZN(n2026) );
  NAND2_X1 U2032 ( .A1(n2026), .A2(n2084), .ZN(n2027) );
  OAI211_X1 U2033 ( .C1(n2029), .C2(n2357), .A(n2028), .B(n2027), .ZN(n2030)
         );
  AOI21_X1 U2034 ( .B1(regfile_wdata_wb_i[25]), .B2(n2100), .A(n2030), .ZN(
        n2031) );
  OAI21_X1 U2035 ( .B1(n2665), .B2(n2035), .A(n2034), .ZN(n2526) );
  NAND3_X1 U2037 ( .A1(instr_rdata_i[22]), .A2(n2604), .A3(instr_rdata_i[23]), 
        .ZN(n2082) );
  INV_X1 U2038 ( .A(n2082), .ZN(n2041) );
  NAND2_X1 U2039 ( .A1(n2116), .A2(regfile_data_rb_id[26]), .ZN(n2038) );
  AOI21_X1 U2040 ( .B1(n2096), .B2(n2683), .A(n2095), .ZN(n2037) );
  OAI211_X1 U2041 ( .C1(n2114), .C2(n2039), .A(n2038), .B(n2037), .ZN(n2040)
         );
  AOI21_X1 U2042 ( .B1(n2041), .B2(n2084), .A(n2040), .ZN(n2043) );
  NAND2_X1 U2043 ( .A1(regfile_data_rc_id[26]), .A2(n2117), .ZN(n2042) );
  OAI211_X1 U2044 ( .C1(n2369), .C2(n2120), .A(n2043), .B(n2042), .ZN(n2044)
         );
  AOI21_X1 U2045 ( .B1(regfile_alu_wdata_fw_i[26]), .B2(n2122), .A(n2044), 
        .ZN(n2047) );
  OR2_X1 U2046 ( .A1(n2045), .A2(n2125), .ZN(n2046) );
  NOR2_X1 U2047 ( .A1(n2050), .A2(n2082), .ZN(n2051) );
  XNOR2_X1 U2048 ( .A(n2051), .B(n2082), .ZN(n2066) );
  NAND2_X1 U2049 ( .A1(n2116), .A2(regfile_data_rb_id[27]), .ZN(n2053) );
  AOI21_X1 U2050 ( .B1(n2678), .B2(n2096), .A(n2095), .ZN(n2052) );
  OAI211_X1 U2051 ( .C1(n2114), .C2(n2054), .A(n2053), .B(n2052), .ZN(n2055)
         );
  AOI21_X1 U2052 ( .B1(n2066), .B2(n2084), .A(n2055), .ZN(n2057) );
  NAND2_X1 U2053 ( .A1(regfile_data_rc_id[27]), .A2(n2117), .ZN(n2056) );
  OAI211_X1 U2054 ( .C1(n2378), .C2(n2120), .A(n2057), .B(n2056), .ZN(n2058)
         );
  AOI21_X1 U2055 ( .B1(regfile_alu_wdata_fw_i[27]), .B2(n2122), .A(n2058), 
        .ZN(n2061) );
  OR2_X1 U2056 ( .A1(n2059), .A2(n2125), .ZN(n2060) );
  NAND2_X1 U2058 ( .A1(regfile_alu_wdata_fw_i[28]), .A2(n2122), .ZN(n2076) );
  OR2_X1 U2059 ( .A1(n2064), .A2(n2082), .ZN(n2065) );
  XNOR2_X1 U2060 ( .A(n2066), .B(n2065), .ZN(n2067) );
  NAND2_X1 U2061 ( .A1(n2067), .A2(n2084), .ZN(n2073) );
  NAND2_X1 U2062 ( .A1(regfile_data_rc_id[28]), .A2(n2117), .ZN(n2072) );
  AOI21_X1 U2063 ( .B1(n2668), .B2(n2096), .A(n2095), .ZN(n2068) );
  OAI21_X1 U2064 ( .B1(n2114), .B2(n2069), .A(n2068), .ZN(n2070) );
  AOI21_X1 U2065 ( .B1(n2116), .B2(regfile_data_rb_id[28]), .A(n2070), .ZN(
        n2071) );
  NAND3_X1 U2066 ( .A1(n2073), .A2(n2072), .A3(n2071), .ZN(n2074) );
  AOI21_X1 U2067 ( .B1(regfile_wdata_wb_i[28]), .B2(n2100), .A(n2074), .ZN(
        n2075) );
  NAND2_X1 U2068 ( .A1(n2078), .A2(n2077), .ZN(n2528) );
  NAND2_X1 U2070 ( .A1(regfile_wdata_wb_i[29]), .A2(n2100), .ZN(n2089) );
  AOI21_X1 U2071 ( .B1(instr_rdata_i[29]), .B2(n2096), .A(n2095), .ZN(n2079)
         );
  OAI21_X1 U2072 ( .B1(n2114), .B2(n2080), .A(n2079), .ZN(n2081) );
  AOI21_X1 U2073 ( .B1(n2116), .B2(regfile_data_rb_id[29]), .A(n2081), .ZN(
        n2088) );
  NOR2_X1 U2074 ( .A1(n2083), .A2(n2082), .ZN(n2085) );
  NAND2_X1 U2075 ( .A1(n2085), .A2(n2084), .ZN(n2087) );
  NAND2_X1 U2076 ( .A1(regfile_data_rc_id[29]), .A2(n2117), .ZN(n2086) );
  NAND4_X1 U2077 ( .A1(n2089), .A2(n2088), .A3(n2087), .A4(n2086), .ZN(n2090)
         );
  AOI21_X1 U2078 ( .B1(regfile_alu_wdata_fw_i[29]), .B2(n2122), .A(n2090), 
        .ZN(n2091) );
  OAI21_X1 U2079 ( .B1(n2092), .B2(n2125), .A(n2091), .ZN(n2093) );
  INV_X1 U2080 ( .A(n2093), .ZN(n2094) );
  INV_X1 U2082 ( .A(regfile_data_ra_id[30]), .ZN(n2098) );
  AOI21_X1 U2083 ( .B1(instr_rdata_i[30]), .B2(n2096), .A(n2095), .ZN(n2097)
         );
  OAI21_X1 U2084 ( .B1(n2114), .B2(n2098), .A(n2097), .ZN(n2099) );
  AOI21_X1 U2085 ( .B1(n2116), .B2(regfile_data_rb_id[30]), .A(n2099), .ZN(
        n2103) );
  NAND2_X1 U2086 ( .A1(regfile_data_rc_id[30]), .A2(n2117), .ZN(n2102) );
  NAND2_X1 U2087 ( .A1(regfile_wdata_wb_i[30]), .A2(n2100), .ZN(n2101) );
  NAND3_X1 U2088 ( .A1(n2103), .A2(n2102), .A3(n2101), .ZN(n2104) );
  AOI21_X1 U2089 ( .B1(regfile_alu_wdata_fw_i[30]), .B2(n2122), .A(n2104), 
        .ZN(n2105) );
  INV_X1 U2091 ( .A(regfile_data_ra_id[31]), .ZN(n2113) );
  NAND4_X1 U2092 ( .A1(n2110), .A2(instr_rdata_i[31]), .A3(n2109), .A4(n2108), 
        .ZN(n2111) );
  OAI211_X1 U2093 ( .C1(n2114), .C2(n2113), .A(n2112), .B(n2111), .ZN(n2115)
         );
  AOI21_X1 U2094 ( .B1(n2116), .B2(regfile_data_rb_id[31]), .A(n2115), .ZN(
        n2119) );
  NAND2_X1 U2095 ( .A1(regfile_data_rc_id[31]), .A2(n2117), .ZN(n2118) );
  OAI211_X1 U2096 ( .C1(n2420), .C2(n2120), .A(n2119), .B(n2118), .ZN(n2121)
         );
  AOI21_X1 U2097 ( .B1(regfile_alu_wdata_fw_i[31]), .B2(n2122), .A(n2121), 
        .ZN(n2123) );
  INV_X1 U2098 ( .A(alu_op_a_mux_sel[2]), .ZN(n2127) );
  NAND2_X1 U2099 ( .A1(alu_op_a_mux_sel[1]), .A2(n2127), .ZN(n2132) );
  INV_X1 U2100 ( .A(n2132), .ZN(n2128) );
  NAND2_X1 U2101 ( .A1(n2128), .A2(alu_op_a_mux_sel[0]), .ZN(n2220) );
  INV_X1 U2102 ( .A(n2220), .ZN(n2269) );
  NOR2_X1 U2103 ( .A1(alu_op_a_mux_sel[0]), .A2(alu_op_a_mux_sel[1]), .ZN(
        n2129) );
  NAND2_X1 U2104 ( .A1(n2129), .A2(alu_op_a_mux_sel[2]), .ZN(n2219) );
  INV_X1 U2105 ( .A(n2219), .ZN(n2270) );
  AOI22_X1 U2106 ( .A1(n2269), .A2(n1205), .B1(n1206), .B2(n2270), .ZN(n2138)
         );
  OAI21_X1 U2107 ( .B1(alu_op_a_mux_sel[2]), .B2(n2129), .A(n2219), .ZN(n2223)
         );
  INV_X1 U2108 ( .A(n2223), .ZN(n2277) );
  NOR2_X1 U2109 ( .A1(n2130), .A2(n2223), .ZN(n2400) );
  INV_X1 U2110 ( .A(n2400), .ZN(n2275) );
  INV_X1 U2111 ( .A(alu_op_a_mux_sel[0]), .ZN(n2131) );
  OR3_X1 U2112 ( .A1(n2131), .A2(alu_op_a_mux_sel[2]), .A3(alu_op_a_mux_sel[1]), .ZN(n2273) );
  NOR3_X1 U2113 ( .A1(n2132), .A2(alu_op_a_mux_sel[0]), .A3(imm_a_mux_sel_0_), 
        .ZN(n2162) );
  AOI22_X1 U2114 ( .A1(n2410), .A2(pc_id_i[0]), .B1(n2162), .B2(n113), .ZN(
        n2133) );
  OAI21_X1 U2115 ( .B1(n2275), .B2(n2134), .A(n2133), .ZN(n2135) );
  AOI21_X1 U2116 ( .B1(n2136), .B2(n2277), .A(n2135), .ZN(n2137) );
  NAND2_X1 U2117 ( .A1(n2138), .A2(n2137), .ZN(n2534) );
  AOI22_X1 U2119 ( .A1(n2269), .A2(n1229), .B1(n2658), .B2(n2277), .ZN(n2146)
         );
  AOI22_X1 U2120 ( .A1(n2410), .A2(pc_id_i[1]), .B1(n2162), .B2(n80), .ZN(
        n2142) );
  NAND2_X1 U2121 ( .A1(regfile_data_rc_id[1]), .A2(n107), .ZN(n2141) );
  OAI211_X1 U2122 ( .C1(n2143), .C2(n2219), .A(n2142), .B(n2141), .ZN(n2144)
         );
  INV_X1 U2123 ( .A(n2144), .ZN(n2145) );
  NAND2_X1 U2124 ( .A1(n2146), .A2(n2145), .ZN(n2535) );
  OAI22_X1 U2126 ( .A1(n2148), .A2(n2220), .B1(n2147), .B2(n2219), .ZN(n2149)
         );
  INV_X1 U2127 ( .A(n2149), .ZN(n2156) );
  NOR2_X1 U2128 ( .A1(n2150), .A2(n2223), .ZN(n2154) );
  AOI22_X1 U2129 ( .A1(n2410), .A2(pc_id_i[2]), .B1(n2162), .B2(n110), .ZN(
        n2151) );
  OAI21_X1 U2130 ( .B1(n2275), .B2(n2152), .A(n2151), .ZN(n2153) );
  NOR2_X1 U2131 ( .A1(n2154), .A2(n2153), .ZN(n2155) );
  NAND2_X1 U2132 ( .A1(n2156), .A2(n2155), .ZN(n2536) );
  AOI22_X1 U2134 ( .A1(n2410), .A2(pc_id_i[3]), .B1(n2162), .B2(n33), .ZN(
        n2157) );
  OAI21_X1 U2135 ( .B1(n1664), .B2(n2223), .A(n2157), .ZN(n2158) );
  INV_X1 U2136 ( .A(n2158), .ZN(n2160) );
  OR2_X1 U2137 ( .A1(n1663), .A2(n2219), .ZN(n2159) );
  OAI211_X1 U2138 ( .C1(n2161), .C2(n2220), .A(n2160), .B(n2159), .ZN(n2538)
         );
  AOI22_X1 U2140 ( .A1(n2410), .A2(pc_id_i[4]), .B1(n2162), .B2(n116), .ZN(
        n2163) );
  OAI21_X1 U2141 ( .B1(n1681), .B2(n2223), .A(n2163), .ZN(n2165) );
  INV_X1 U2142 ( .A(n2165), .ZN(n2167) );
  OR2_X1 U2143 ( .A1(n1680), .A2(n2219), .ZN(n2166) );
  OAI211_X1 U2144 ( .C1(n1685), .C2(n2220), .A(n2167), .B(n2166), .ZN(n2539)
         );
  AOI22_X1 U2146 ( .A1(n2269), .A2(n2660), .B1(n1693), .B2(n2270), .ZN(n2169)
         );
  AOI22_X1 U2147 ( .A1(n1688), .A2(n2277), .B1(pc_id_i[5]), .B2(n2410), .ZN(
        n2168) );
  NAND2_X1 U2148 ( .A1(n2169), .A2(n2168), .ZN(n2540) );
  INV_X1 U2150 ( .A(n2275), .ZN(n2411) );
  AOI22_X1 U2151 ( .A1(n2411), .A2(n32), .B1(n2410), .B2(pc_id_i[6]), .ZN(
        n2170) );
  OAI21_X1 U2152 ( .B1(n2171), .B2(n2223), .A(n2170), .ZN(n2172) );
  INV_X1 U2153 ( .A(n2172), .ZN(n2175) );
  OR2_X1 U2154 ( .A1(n2173), .A2(n2220), .ZN(n2174) );
  OAI211_X1 U2155 ( .C1(n2176), .C2(n2219), .A(n2175), .B(n2174), .ZN(n2541)
         );
  NOR2_X1 U2157 ( .A1(n2177), .A2(n2223), .ZN(n2190) );
  OR2_X1 U2158 ( .A1(n2178), .A2(n2219), .ZN(n2261) );
  NOR2_X1 U2159 ( .A1(n2182), .A2(n2261), .ZN(n2184) );
  NAND2_X1 U2160 ( .A1(n2179), .A2(n2277), .ZN(n2208) );
  AOI22_X1 U2161 ( .A1(n2411), .A2(n31), .B1(n2410), .B2(pc_id_i[7]), .ZN(
        n2181) );
  NAND2_X1 U2162 ( .A1(regfile_data_rc_id[7]), .A2(n107), .ZN(n2180) );
  OAI211_X1 U2163 ( .C1(n2182), .C2(n2208), .A(n2181), .B(n2180), .ZN(n2183)
         );
  AOI211_X1 U2164 ( .C1(regfile_alu_wdata_fw_i[7]), .C2(n2190), .A(n2184), .B(
        n2183), .ZN(n2187) );
  NOR2_X1 U2165 ( .A1(n2185), .A2(n2219), .ZN(n2189) );
  NAND2_X1 U2166 ( .A1(regfile_alu_wdata_fw_i[7]), .A2(n2189), .ZN(n2186) );
  OAI211_X1 U2167 ( .C1(n2188), .C2(n2220), .A(n2187), .B(n2186), .ZN(n2542)
         );
  INV_X1 U2169 ( .A(n2189), .ZN(n2266) );
  INV_X1 U2170 ( .A(n2190), .ZN(n2206) );
  NAND2_X1 U2171 ( .A1(n2266), .A2(n2206), .ZN(n2422) );
  INV_X1 U2172 ( .A(n2261), .ZN(n2192) );
  INV_X1 U2173 ( .A(n2208), .ZN(n2191) );
  NOR2_X1 U2174 ( .A1(n2192), .A2(n2191), .ZN(n2298) );
  AOI22_X1 U2175 ( .A1(n2411), .A2(n24), .B1(n2410), .B2(pc_id_i[8]), .ZN(
        n2194) );
  NAND2_X1 U2176 ( .A1(regfile_data_rc_id[8]), .A2(n107), .ZN(n2193) );
  OAI211_X1 U2177 ( .C1(n2195), .C2(n2298), .A(n2194), .B(n2193), .ZN(n2196)
         );
  AOI21_X1 U2178 ( .B1(regfile_alu_wdata_fw_i[8]), .B2(n2422), .A(n2196), .ZN(
        n2197) );
  OAI21_X1 U2179 ( .B1(n2198), .B2(n2220), .A(n2197), .ZN(n2543) );
  AOI22_X1 U2181 ( .A1(n2411), .A2(regfile_data_ra_id[9]), .B1(n2410), .B2(
        pc_id_i[9]), .ZN(n2200) );
  NAND2_X1 U2182 ( .A1(regfile_data_rc_id[9]), .A2(n107), .ZN(n2199) );
  OAI211_X1 U2183 ( .C1(n2201), .C2(n2298), .A(n2200), .B(n2199), .ZN(n2202)
         );
  AOI21_X1 U2184 ( .B1(regfile_alu_wdata_fw_i[9]), .B2(n2422), .A(n2202), .ZN(
        n2203) );
  OAI21_X1 U2185 ( .B1(n2204), .B2(n2220), .A(n2203), .ZN(n2544) );
  INV_X1 U2187 ( .A(regfile_alu_wdata_fw_i[10]), .ZN(n2218) );
  NAND2_X1 U2188 ( .A1(n2424), .A2(n2206), .ZN(n2264) );
  NAND2_X1 U2189 ( .A1(n2207), .A2(n2269), .ZN(n2419) );
  NAND2_X1 U2190 ( .A1(n2419), .A2(n2208), .ZN(n2259) );
  INV_X1 U2191 ( .A(regfile_data_rb_id[10]), .ZN(n2212) );
  NAND2_X1 U2192 ( .A1(n2209), .A2(n2269), .ZN(n2300) );
  NAND2_X1 U2193 ( .A1(n107), .A2(regfile_data_rc_id[10]), .ZN(n2211) );
  AOI22_X1 U2194 ( .A1(n2411), .A2(n47), .B1(n2410), .B2(pc_id_i[10]), .ZN(
        n2210) );
  OAI211_X1 U2195 ( .C1(n2212), .C2(n2300), .A(n2211), .B(n2210), .ZN(n2213)
         );
  AOI21_X1 U2196 ( .B1(regfile_wdata_wb_i[10]), .B2(n2259), .A(n2213), .ZN(
        n2214) );
  OAI21_X1 U2197 ( .B1(n2215), .B2(n2261), .A(n2214), .ZN(n2216) );
  AOI21_X1 U2198 ( .B1(regfile_alu_wdata_fw_i[10]), .B2(n2264), .A(n2216), 
        .ZN(n2217) );
  OAI21_X1 U2199 ( .B1(n2218), .B2(n2266), .A(n2217), .ZN(n2545) );
  OAI22_X1 U2201 ( .A1(n1778), .A2(n2220), .B1(n1780), .B2(n2219), .ZN(n2221)
         );
  INV_X1 U2202 ( .A(n2221), .ZN(n2227) );
  AOI22_X1 U2203 ( .A1(n2411), .A2(n25), .B1(n2410), .B2(pc_id_i[11]), .ZN(
        n2222) );
  OAI21_X1 U2204 ( .B1(n2224), .B2(n2223), .A(n2222), .ZN(n2225) );
  INV_X1 U2205 ( .A(n2225), .ZN(n2226) );
  NAND2_X1 U2206 ( .A1(n2227), .A2(n2226), .ZN(n2546) );
  INV_X1 U2208 ( .A(regfile_alu_wdata_fw_i[12]), .ZN(n2236) );
  INV_X1 U2209 ( .A(regfile_wdata_wb_i[12]), .ZN(n2233) );
  INV_X1 U2210 ( .A(regfile_data_rb_id[12]), .ZN(n2230) );
  NAND2_X1 U2211 ( .A1(n107), .A2(regfile_data_rc_id[12]), .ZN(n2229) );
  AOI22_X1 U2212 ( .A1(n2411), .A2(regfile_data_ra_id[12]), .B1(n2410), .B2(
        pc_id_i[12]), .ZN(n2228) );
  OAI211_X1 U2213 ( .C1(n2300), .C2(n2230), .A(n2229), .B(n2228), .ZN(n2231)
         );
  AOI21_X1 U2214 ( .B1(regfile_wdata_wb_i[12]), .B2(n2259), .A(n2231), .ZN(
        n2232) );
  OAI21_X1 U2215 ( .B1(n2233), .B2(n2261), .A(n2232), .ZN(n2234) );
  AOI21_X1 U2216 ( .B1(regfile_alu_wdata_fw_i[12]), .B2(n2264), .A(n2234), 
        .ZN(n2235) );
  OAI21_X1 U2217 ( .B1(n2236), .B2(n2266), .A(n2235), .ZN(n2547) );
  INV_X1 U2219 ( .A(regfile_alu_wdata_fw_i[13]), .ZN(n2245) );
  INV_X1 U2220 ( .A(regfile_wdata_wb_i[13]), .ZN(n2242) );
  INV_X1 U2221 ( .A(regfile_data_rb_id[13]), .ZN(n2239) );
  NAND2_X1 U2222 ( .A1(n107), .A2(regfile_data_rc_id[13]), .ZN(n2238) );
  AOI22_X1 U2223 ( .A1(n2411), .A2(regfile_data_ra_id[13]), .B1(n2410), .B2(
        pc_id_i[13]), .ZN(n2237) );
  OAI211_X1 U2224 ( .C1(n2300), .C2(n2239), .A(n2238), .B(n2237), .ZN(n2240)
         );
  AOI21_X1 U2225 ( .B1(regfile_wdata_wb_i[13]), .B2(n2259), .A(n2240), .ZN(
        n2241) );
  OAI21_X1 U2226 ( .B1(n2242), .B2(n2261), .A(n2241), .ZN(n2243) );
  AOI21_X1 U2227 ( .B1(regfile_alu_wdata_fw_i[13]), .B2(n2264), .A(n2243), 
        .ZN(n2244) );
  OAI21_X1 U2228 ( .B1(n2245), .B2(n2266), .A(n2244), .ZN(n2548) );
  INV_X1 U2230 ( .A(regfile_alu_wdata_fw_i[14]), .ZN(n2254) );
  INV_X1 U2231 ( .A(regfile_wdata_wb_i[14]), .ZN(n2251) );
  INV_X1 U2232 ( .A(regfile_data_rb_id[14]), .ZN(n2248) );
  NAND2_X1 U2233 ( .A1(n107), .A2(regfile_data_rc_id[14]), .ZN(n2247) );
  AOI22_X1 U2234 ( .A1(n2411), .A2(regfile_data_ra_id[14]), .B1(n2410), .B2(
        pc_id_i[14]), .ZN(n2246) );
  OAI211_X1 U2235 ( .C1(n2300), .C2(n2248), .A(n2247), .B(n2246), .ZN(n2249)
         );
  AOI21_X1 U2236 ( .B1(regfile_wdata_wb_i[14]), .B2(n2259), .A(n2249), .ZN(
        n2250) );
  OAI21_X1 U2237 ( .B1(n2251), .B2(n2261), .A(n2250), .ZN(n2252) );
  AOI21_X1 U2238 ( .B1(regfile_alu_wdata_fw_i[14]), .B2(n2264), .A(n2252), 
        .ZN(n2253) );
  OAI21_X1 U2239 ( .B1(n2254), .B2(n2266), .A(n2253), .ZN(n2549) );
  INV_X1 U2241 ( .A(n2663), .ZN(n2267) );
  INV_X1 U2242 ( .A(regfile_data_rb_id[15]), .ZN(n2257) );
  NAND2_X1 U2243 ( .A1(n107), .A2(regfile_data_rc_id[15]), .ZN(n2256) );
  AOI22_X1 U2244 ( .A1(n2411), .A2(regfile_data_ra_id[15]), .B1(n2410), .B2(
        pc_id_i[15]), .ZN(n2255) );
  OAI211_X1 U2245 ( .C1(n2300), .C2(n2257), .A(n2256), .B(n2255), .ZN(n2258)
         );
  AOI21_X1 U2246 ( .B1(regfile_wdata_wb_i[15]), .B2(n2259), .A(n2258), .ZN(
        n2260) );
  OAI21_X1 U2247 ( .B1(n2262), .B2(n2261), .A(n2260), .ZN(n2263) );
  AOI21_X1 U2248 ( .B1(n2663), .B2(n2264), .A(n2263), .ZN(n2265) );
  OAI21_X1 U2249 ( .B1(n2267), .B2(n2266), .A(n2265), .ZN(n2550) );
  AOI22_X1 U2251 ( .A1(n2270), .A2(n1867), .B1(n1866), .B2(n2269), .ZN(n2279)
         );
  INV_X1 U2252 ( .A(pc_id_i[16]), .ZN(n2272) );
  OAI22_X1 U2253 ( .A1(n2275), .A2(n2274), .B1(n2273), .B2(n2272), .ZN(n2276)
         );
  AOI21_X1 U2254 ( .B1(n2271), .B2(n2277), .A(n2276), .ZN(n2278) );
  NAND2_X1 U2255 ( .A1(n2279), .A2(n2278), .ZN(n2552) );
  INV_X1 U2257 ( .A(regfile_alu_wdata_fw_i[17]), .ZN(n2288) );
  INV_X1 U2258 ( .A(regfile_data_rb_id[17]), .ZN(n2281) );
  AOI22_X1 U2259 ( .A1(n2411), .A2(regfile_data_ra_id[17]), .B1(n2410), .B2(
        pc_id_i[17]), .ZN(n2280) );
  OAI21_X1 U2260 ( .B1(n2300), .B2(n2281), .A(n2280), .ZN(n2283) );
  NOR2_X1 U2261 ( .A1(n2285), .A2(n2298), .ZN(n2282) );
  AOI211_X1 U2262 ( .C1(n107), .C2(regfile_data_rc_id[17]), .A(n2283), .B(
        n2282), .ZN(n2284) );
  OAI21_X1 U2263 ( .B1(n2285), .B2(n2419), .A(n2284), .ZN(n2286) );
  AOI21_X1 U2264 ( .B1(regfile_alu_wdata_fw_i[17]), .B2(n2422), .A(n2286), 
        .ZN(n2287) );
  OAI21_X1 U2265 ( .B1(n2288), .B2(n2424), .A(n2287), .ZN(n2553) );
  INV_X1 U2267 ( .A(regfile_alu_wdata_fw_i[18]), .ZN(n2297) );
  INV_X1 U2268 ( .A(regfile_data_rb_id[18]), .ZN(n2290) );
  AOI22_X1 U2269 ( .A1(n2411), .A2(regfile_data_ra_id[18]), .B1(n2410), .B2(
        pc_id_i[18]), .ZN(n2289) );
  OAI21_X1 U2270 ( .B1(n2300), .B2(n2290), .A(n2289), .ZN(n2292) );
  NOR2_X1 U2271 ( .A1(n2294), .A2(n2298), .ZN(n2291) );
  AOI211_X1 U2272 ( .C1(n107), .C2(regfile_data_rc_id[18]), .A(n2292), .B(
        n2291), .ZN(n2293) );
  OAI21_X1 U2273 ( .B1(n2294), .B2(n2419), .A(n2293), .ZN(n2295) );
  AOI21_X1 U2274 ( .B1(regfile_alu_wdata_fw_i[18]), .B2(n2422), .A(n2295), 
        .ZN(n2296) );
  OAI21_X1 U2275 ( .B1(n2297), .B2(n2424), .A(n2296), .ZN(n2554) );
  INV_X1 U2277 ( .A(regfile_alu_wdata_fw_i[19]), .ZN(n2309) );
  INV_X1 U2278 ( .A(n2298), .ZN(n2417) );
  AOI22_X1 U2279 ( .A1(n2400), .A2(regfile_data_ra_id[19]), .B1(n2410), .B2(
        pc_id_i[19]), .ZN(n2302) );
  INV_X1 U2280 ( .A(n2300), .ZN(n2412) );
  NAND2_X1 U2281 ( .A1(n2412), .A2(regfile_data_rb_id[19]), .ZN(n2301) );
  OAI211_X1 U2282 ( .C1(n2299), .C2(n2303), .A(n2302), .B(n2301), .ZN(n2304)
         );
  AOI21_X1 U2283 ( .B1(regfile_wdata_wb_i[19]), .B2(n2417), .A(n2304), .ZN(
        n2305) );
  OAI21_X1 U2284 ( .B1(n2306), .B2(n2419), .A(n2305), .ZN(n2307) );
  AOI21_X1 U2285 ( .B1(regfile_alu_wdata_fw_i[19]), .B2(n2422), .A(n2307), 
        .ZN(n2308) );
  OAI21_X1 U2286 ( .B1(n2309), .B2(n2424), .A(n2308), .ZN(n2555) );
  INV_X1 U2288 ( .A(regfile_alu_wdata_fw_i[20]), .ZN(n2318) );
  AOI22_X1 U2289 ( .A1(n2400), .A2(regfile_data_ra_id[20]), .B1(n2410), .B2(
        pc_id_i[20]), .ZN(n2311) );
  NAND2_X1 U2290 ( .A1(n2412), .A2(regfile_data_rb_id[20]), .ZN(n2310) );
  OAI211_X1 U2291 ( .C1(n2299), .C2(n2312), .A(n2311), .B(n2310), .ZN(n2313)
         );
  AOI21_X1 U2292 ( .B1(regfile_wdata_wb_i[20]), .B2(n2417), .A(n2313), .ZN(
        n2314) );
  OAI21_X1 U2293 ( .B1(n2315), .B2(n2419), .A(n2314), .ZN(n2316) );
  AOI21_X1 U2294 ( .B1(regfile_alu_wdata_fw_i[20]), .B2(n2422), .A(n2316), 
        .ZN(n2317) );
  OAI21_X1 U2295 ( .B1(n2318), .B2(n2424), .A(n2317), .ZN(n2556) );
  INV_X1 U2297 ( .A(regfile_alu_wdata_fw_i[21]), .ZN(n2327) );
  AOI22_X1 U2298 ( .A1(n2411), .A2(n2644), .B1(n2410), .B2(pc_id_i[21]), .ZN(
        n2320) );
  NAND2_X1 U2299 ( .A1(n2412), .A2(regfile_data_rb_id[21]), .ZN(n2319) );
  OAI211_X1 U2300 ( .C1(n2299), .C2(n2321), .A(n2320), .B(n2319), .ZN(n2322)
         );
  AOI21_X1 U2301 ( .B1(regfile_wdata_wb_i[21]), .B2(n2417), .A(n2322), .ZN(
        n2323) );
  OAI21_X1 U2302 ( .B1(n2324), .B2(n2419), .A(n2323), .ZN(n2325) );
  AOI21_X1 U2303 ( .B1(regfile_alu_wdata_fw_i[21]), .B2(n2422), .A(n2325), 
        .ZN(n2326) );
  OAI21_X1 U2304 ( .B1(n2327), .B2(n2424), .A(n2326), .ZN(n2557) );
  INV_X1 U2306 ( .A(regfile_alu_wdata_fw_i[22]), .ZN(n2336) );
  AOI22_X1 U2307 ( .A1(n2400), .A2(regfile_data_ra_id[22]), .B1(n2410), .B2(
        pc_id_i[22]), .ZN(n2329) );
  NAND2_X1 U2308 ( .A1(n2412), .A2(regfile_data_rb_id[22]), .ZN(n2328) );
  OAI211_X1 U2309 ( .C1(n2299), .C2(n2330), .A(n2329), .B(n2328), .ZN(n2331)
         );
  AOI21_X1 U2310 ( .B1(regfile_wdata_wb_i[22]), .B2(n2417), .A(n2331), .ZN(
        n2332) );
  OAI21_X1 U2311 ( .B1(n2333), .B2(n2419), .A(n2332), .ZN(n2334) );
  AOI21_X1 U2312 ( .B1(regfile_alu_wdata_fw_i[22]), .B2(n2422), .A(n2334), 
        .ZN(n2335) );
  OAI21_X1 U2313 ( .B1(n2336), .B2(n2424), .A(n2335), .ZN(n2558) );
  INV_X1 U2315 ( .A(regfile_alu_wdata_fw_i[23]), .ZN(n2345) );
  AOI22_X1 U2316 ( .A1(n2411), .A2(regfile_data_ra_id[23]), .B1(n2410), .B2(
        pc_id_i[23]), .ZN(n2338) );
  NAND2_X1 U2317 ( .A1(n2412), .A2(regfile_data_rb_id[23]), .ZN(n2337) );
  OAI211_X1 U2318 ( .C1(n2299), .C2(n2339), .A(n2338), .B(n2337), .ZN(n2340)
         );
  AOI21_X1 U2319 ( .B1(regfile_wdata_wb_i[23]), .B2(n2417), .A(n2340), .ZN(
        n2341) );
  OAI21_X1 U2320 ( .B1(n2342), .B2(n2419), .A(n2341), .ZN(n2343) );
  AOI21_X1 U2321 ( .B1(regfile_alu_wdata_fw_i[23]), .B2(n2422), .A(n2343), 
        .ZN(n2344) );
  OAI21_X1 U2322 ( .B1(n2345), .B2(n2424), .A(n2344), .ZN(n2559) );
  INV_X1 U2324 ( .A(regfile_alu_wdata_fw_i[24]), .ZN(n2354) );
  AOI22_X1 U2325 ( .A1(n2400), .A2(regfile_data_ra_id[24]), .B1(n2410), .B2(
        pc_id_i[24]), .ZN(n2347) );
  NAND2_X1 U2326 ( .A1(n2412), .A2(regfile_data_rb_id[24]), .ZN(n2346) );
  OAI211_X1 U2327 ( .C1(n2299), .C2(n2348), .A(n2347), .B(n2346), .ZN(n2349)
         );
  AOI21_X1 U2328 ( .B1(regfile_wdata_wb_i[24]), .B2(n2417), .A(n2349), .ZN(
        n2350) );
  OAI21_X1 U2329 ( .B1(n2351), .B2(n2419), .A(n2350), .ZN(n2352) );
  AOI21_X1 U2330 ( .B1(regfile_alu_wdata_fw_i[24]), .B2(n2422), .A(n2352), 
        .ZN(n2353) );
  OAI21_X1 U2331 ( .B1(n2354), .B2(n2424), .A(n2353), .ZN(n2560) );
  INV_X1 U2333 ( .A(regfile_alu_wdata_fw_i[25]), .ZN(n2363) );
  AOI22_X1 U2334 ( .A1(n2411), .A2(regfile_data_ra_id[25]), .B1(n2410), .B2(
        pc_id_i[25]), .ZN(n2356) );
  NAND2_X1 U2335 ( .A1(n2412), .A2(regfile_data_rb_id[25]), .ZN(n2355) );
  OAI211_X1 U2336 ( .C1(n2299), .C2(n2357), .A(n2356), .B(n2355), .ZN(n2358)
         );
  AOI21_X1 U2337 ( .B1(regfile_wdata_wb_i[25]), .B2(n2417), .A(n2358), .ZN(
        n2359) );
  OAI21_X1 U2338 ( .B1(n2360), .B2(n2419), .A(n2359), .ZN(n2361) );
  AOI21_X1 U2339 ( .B1(regfile_alu_wdata_fw_i[25]), .B2(n2422), .A(n2361), 
        .ZN(n2362) );
  OAI21_X1 U2340 ( .B1(n2363), .B2(n2424), .A(n2362), .ZN(n2561) );
  AOI22_X1 U2342 ( .A1(n2400), .A2(regfile_data_ra_id[26]), .B1(n2410), .B2(
        pc_id_i[26]), .ZN(n2365) );
  NAND2_X1 U2343 ( .A1(n2412), .A2(regfile_data_rb_id[26]), .ZN(n2364) );
  OAI211_X1 U2344 ( .C1(n2299), .C2(n2366), .A(n2365), .B(n2364), .ZN(n2367)
         );
  AOI21_X1 U2345 ( .B1(regfile_wdata_wb_i[26]), .B2(n2417), .A(n2367), .ZN(
        n2368) );
  OAI21_X1 U2346 ( .B1(n2369), .B2(n2419), .A(n2368), .ZN(n2370) );
  AOI21_X1 U2347 ( .B1(regfile_alu_wdata_fw_i[26]), .B2(n2422), .A(n2370), 
        .ZN(n2371) );
  OAI21_X1 U2348 ( .B1(n2372), .B2(n2424), .A(n2371), .ZN(n2562) );
  INV_X1 U2350 ( .A(regfile_alu_wdata_fw_i[27]), .ZN(n2381) );
  AOI22_X1 U2351 ( .A1(n2400), .A2(regfile_data_ra_id[27]), .B1(n2410), .B2(
        pc_id_i[27]), .ZN(n2374) );
  NAND2_X1 U2352 ( .A1(n2412), .A2(regfile_data_rb_id[27]), .ZN(n2373) );
  OAI211_X1 U2353 ( .C1(n2299), .C2(n2375), .A(n2374), .B(n2373), .ZN(n2376)
         );
  AOI21_X1 U2354 ( .B1(regfile_wdata_wb_i[27]), .B2(n2417), .A(n2376), .ZN(
        n2377) );
  OAI21_X1 U2355 ( .B1(n2378), .B2(n2419), .A(n2377), .ZN(n2379) );
  AOI21_X1 U2356 ( .B1(regfile_alu_wdata_fw_i[27]), .B2(n2422), .A(n2379), 
        .ZN(n2380) );
  OAI21_X1 U2357 ( .B1(n2381), .B2(n2424), .A(n2380), .ZN(n2563) );
  INV_X1 U2359 ( .A(regfile_alu_wdata_fw_i[28]), .ZN(n2390) );
  AOI22_X1 U2360 ( .A1(n2400), .A2(regfile_data_ra_id[28]), .B1(n2410), .B2(
        pc_id_i[28]), .ZN(n2383) );
  NAND2_X1 U2361 ( .A1(n2412), .A2(regfile_data_rb_id[28]), .ZN(n2382) );
  OAI211_X1 U2362 ( .C1(n2299), .C2(n2384), .A(n2383), .B(n2382), .ZN(n2385)
         );
  AOI21_X1 U2363 ( .B1(regfile_wdata_wb_i[28]), .B2(n2417), .A(n2385), .ZN(
        n2386) );
  OAI21_X1 U2364 ( .B1(n2387), .B2(n2419), .A(n2386), .ZN(n2388) );
  AOI21_X1 U2365 ( .B1(regfile_alu_wdata_fw_i[28]), .B2(n2422), .A(n2388), 
        .ZN(n2389) );
  OAI21_X1 U2366 ( .B1(n2390), .B2(n2424), .A(n2389), .ZN(n2564) );
  INV_X1 U2368 ( .A(regfile_alu_wdata_fw_i[29]), .ZN(n2399) );
  AOI22_X1 U2369 ( .A1(n2400), .A2(regfile_data_ra_id[29]), .B1(n2410), .B2(
        pc_id_i[29]), .ZN(n2392) );
  NAND2_X1 U2370 ( .A1(n2412), .A2(regfile_data_rb_id[29]), .ZN(n2391) );
  OAI211_X1 U2371 ( .C1(n2299), .C2(n2393), .A(n2392), .B(n2391), .ZN(n2394)
         );
  AOI21_X1 U2372 ( .B1(regfile_wdata_wb_i[29]), .B2(n2417), .A(n2394), .ZN(
        n2395) );
  OAI21_X1 U2373 ( .B1(n2396), .B2(n2419), .A(n2395), .ZN(n2397) );
  AOI21_X1 U2374 ( .B1(regfile_alu_wdata_fw_i[29]), .B2(n2422), .A(n2397), 
        .ZN(n2398) );
  OAI21_X1 U2375 ( .B1(n2399), .B2(n2424), .A(n2398), .ZN(n2565) );
  INV_X1 U2377 ( .A(regfile_alu_wdata_fw_i[30]), .ZN(n2409) );
  AOI22_X1 U2378 ( .A1(n2400), .A2(regfile_data_ra_id[30]), .B1(n2410), .B2(
        pc_id_i[30]), .ZN(n2402) );
  NAND2_X1 U2379 ( .A1(n2412), .A2(regfile_data_rb_id[30]), .ZN(n2401) );
  OAI211_X1 U2380 ( .C1(n2299), .C2(n2403), .A(n2402), .B(n2401), .ZN(n2404)
         );
  AOI21_X1 U2381 ( .B1(regfile_wdata_wb_i[30]), .B2(n2417), .A(n2404), .ZN(
        n2405) );
  OAI21_X1 U2382 ( .B1(n2406), .B2(n2419), .A(n2405), .ZN(n2407) );
  AOI21_X1 U2383 ( .B1(regfile_alu_wdata_fw_i[30]), .B2(n2422), .A(n2407), 
        .ZN(n2408) );
  OAI21_X1 U2384 ( .B1(n2409), .B2(n2424), .A(n2408), .ZN(n2566) );
  INV_X1 U2386 ( .A(regfile_alu_wdata_fw_i[31]), .ZN(n2425) );
  AOI22_X1 U2387 ( .A1(n2411), .A2(regfile_data_ra_id[31]), .B1(n2410), .B2(
        pc_id_i[31]), .ZN(n2414) );
  NAND2_X1 U2388 ( .A1(n2412), .A2(regfile_data_rb_id[31]), .ZN(n2413) );
  OAI211_X1 U2389 ( .C1(n2299), .C2(n2415), .A(n2414), .B(n2413), .ZN(n2416)
         );
  AOI21_X1 U2390 ( .B1(regfile_wdata_wb_i[31]), .B2(n2417), .A(n2416), .ZN(
        n2418) );
  OAI21_X1 U2391 ( .B1(n2420), .B2(n2419), .A(n2418), .ZN(n2421) );
  AOI21_X1 U2392 ( .B1(regfile_alu_wdata_fw_i[31]), .B2(n2422), .A(n2421), 
        .ZN(n2423) );
  OAI21_X1 U2393 ( .B1(n2425), .B2(n2424), .A(n2423), .ZN(n2568) );
  INV_X1 U2395 ( .A(mult_int_en), .ZN(n2426) );
  NOR2_X1 U2408 ( .A1(data_misaligned_i), .A2(n2434), .ZN(n2456) );
  INV_X1 U2517 ( .A(regfile_alu_we_id), .ZN(n2453) );
  OAI21_X1 U2518 ( .B1(n2453), .B2(n2455), .A(n2452), .ZN(n2459) );
  AOI21_X1 U2519 ( .B1(csr_access_ex_o), .B2(n2455), .A(n2671), .ZN(n2457) );
  NOR2_X1 U2520 ( .A1(n2457), .A2(n2456), .ZN(n2458) );
  MUX2_X1 U2521 ( .A(regfile_alu_we_ex_o), .B(n2459), .S(n2458), .Z(n1352) );
  NAND2_X1 U2563 ( .A1(n638), .A2(n2503), .ZN(n2533) );
  NAND2_X1 U2596 ( .A1(n638), .A2(n2599), .ZN(n2532) );
  NAND2_X1 U2630 ( .A1(n2570), .A2(n2569), .ZN(n2571) );
  AOI21_X1 U2664 ( .B1(n2574), .B2(csr_hwlp_we_i[1]), .A(n897), .ZN(n2572) );
  INV_X1 U2665 ( .A(n2572), .ZN(hwloop_we[1]) );
  AOI21_X1 U2666 ( .B1(n2574), .B2(csr_hwlp_we_i[2]), .A(hwloop_we_int[2]), 
        .ZN(n2573) );
  INV_X1 U2667 ( .A(n2573), .ZN(hwloop_we[2]) );
  MUX2_X1 U2668 ( .A(instr_rdata_i[7]), .B(csr_hwlp_regid_i[0]), .S(n2574), 
        .Z(hwloop_regid_0_) );
  SDFFR_X1 data_req_ex_o_reg ( .D(n3483), .SI(1'b0), .SE(1'b0), .CK(n3504), 
        .RN(rst_n), .Q(data_req_ex_o) );
  SDFFR_X1 branch_in_ex_o_reg ( .D(n3499), .SI(1'b0), .SE(1'b0), .CK(n3504), 
        .RN(rst_n), .Q(branch_in_ex_o) );
  SDFFR_X1 prepost_useincr_ex_o_reg ( .D(n1353), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(rst_n), .Q(prepost_useincr_ex_o), .QN(n2599) );
  SDFFR_X1 data_we_ex_o_reg ( .D(data_we_id), .SI(1'b0), .SE(1'b0), .CK(n3481), 
        .RN(rst_n), .Q(data_we_ex_o) );
  SDFFR_X1 data_type_ex_o_reg_0_ ( .D(data_type_id[0]), .SI(1'b0), .SE(1'b0), 
        .CK(n3481), .RN(rst_n), .Q(data_type_ex_o[0]) );
  SDFFR_X1 data_type_ex_o_reg_1_ ( .D(data_type_id[1]), .SI(1'b0), .SE(1'b0), 
        .CK(n3481), .RN(rst_n), .Q(data_type_ex_o[1]) );
  SDFFR_X1 data_sign_ext_ex_o_reg_0_ ( .D(data_sign_ext_id_0_), .SI(1'b0), 
        .SE(1'b0), .CK(n3481), .RN(rst_n), .Q(data_sign_ext_ex_o[0]) );
  SDFFR_X1 csr_op_ex_o_reg_0_ ( .D(n3500), .SI(1'b0), .SE(1'b0), .CK(n3504), 
        .RN(rst_n), .Q(csr_op_ex_o[0]) );
  SDFFR_X1 csr_op_ex_o_reg_1_ ( .D(n3501), .SI(1'b0), .SE(1'b0), .CK(n3504), 
        .RN(rst_n), .Q(csr_op_ex_o[1]) );
  SDFFR_X1 regfile_alu_waddr_ex_o_reg_0_ ( .D(regfile_alu_waddr_id[0]), .SI(
        1'b0), .SE(1'b0), .CK(n3484), .RN(rst_n), .Q(regfile_alu_waddr_ex_o[0]) );
  SDFFR_X1 regfile_alu_waddr_ex_o_reg_1_ ( .D(regfile_alu_waddr_id[1]), .SI(
        1'b0), .SE(1'b0), .CK(n3484), .RN(rst_n), .Q(regfile_alu_waddr_ex_o[1]) );
  SDFFR_X1 regfile_alu_waddr_ex_o_reg_2_ ( .D(regfile_alu_waddr_id[2]), .SI(
        1'b0), .SE(1'b0), .CK(n3484), .RN(rst_n), .Q(regfile_alu_waddr_ex_o[2]) );
  SDFFR_X1 regfile_alu_waddr_ex_o_reg_3_ ( .D(regfile_alu_waddr_id[3]), .SI(
        1'b0), .SE(1'b0), .CK(n3484), .RN(rst_n), .Q(regfile_alu_waddr_ex_o[3]) );
  SDFFR_X1 regfile_alu_waddr_ex_o_reg_4_ ( .D(regfile_alu_waddr_id[4]), .SI(
        1'b0), .SE(1'b0), .CK(n3484), .RN(rst_n), .Q(regfile_alu_waddr_ex_o[4]) );
  SDFFR_X1 regfile_alu_we_ex_o_reg ( .D(n1352), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(rst_n), .Q(regfile_alu_we_ex_o) );
  SDFFR_X1 regfile_waddr_ex_o_reg_0_ ( .D(instr_rdata_i[7]), .SI(1'b0), .SE(
        1'b0), .CK(n3487), .RN(rst_n), .Q(regfile_waddr_ex_o[0]) );
  SDFFR_X1 regfile_waddr_ex_o_reg_1_ ( .D(instr_rdata_i[8]), .SI(1'b0), .SE(
        1'b0), .CK(n3487), .RN(rst_n), .Q(regfile_waddr_ex_o[1]) );
  SDFFR_X1 regfile_waddr_ex_o_reg_2_ ( .D(instr_rdata_i[9]), .SI(1'b0), .SE(
        1'b0), .CK(n3487), .RN(rst_n), .Q(regfile_waddr_ex_o[2]) );
  SDFFR_X1 regfile_waddr_ex_o_reg_3_ ( .D(instr_rdata_i[10]), .SI(1'b0), .SE(
        1'b0), .CK(n3487), .RN(rst_n), .Q(regfile_waddr_ex_o[3]) );
  SDFFR_X1 regfile_waddr_ex_o_reg_4_ ( .D(instr_rdata_i[11]), .SI(1'b0), .SE(
        1'b0), .CK(n3487), .RN(rst_n), .Q(regfile_waddr_ex_o[4]) );
  SDFFR_X1 regfile_we_ex_o_reg ( .D(n2693), .SI(1'b0), .SE(1'b0), .CK(n3504), 
        .RN(rst_n), .Q(regfile_we_ex_o) );
  SDFFR_X1 mult_dot_signed_ex_o_reg_1_ ( .D(mult_dot_signed[1]), .SI(1'b0), 
        .SE(1'b0), .CK(n3540), .RN(rst_n), .Q(mult_dot_signed_ex_o[1]) );
  SDFFR_X1 mult_clpx_img_ex_o_reg ( .D(instr_rdata_i[25]), .SI(1'b0), .SE(1'b0), .CK(n3540), .RN(rst_n), .Q(mult_clpx_img_ex_o) );
  SDFFR_X1 mult_clpx_shift_ex_o_reg_0_ ( .D(instr_rdata_i[13]), .SI(1'b0), 
        .SE(1'b0), .CK(n3540), .RN(rst_n), .Q(mult_clpx_shift_ex_o[0]) );
  SDFFR_X1 mult_dot_signed_ex_o_reg_0_ ( .D(mult_dot_signed[0]), .SI(1'b0), 
        .SE(1'b0), .CK(n3540), .RN(rst_n), .Q(mult_dot_signed_ex_o[0]) );
  SDFFR_X1 mult_sel_subword_ex_o_reg ( .D(mult_sel_subword), .SI(1'b0), .SE(
        1'b0), .CK(n3538), .RN(rst_n), .QN(mult_sel_subword_ex_o_BAR) );
  SDFFR_X1 mult_signed_mode_ex_o_reg_0_ ( .D(mult_signed_mode[0]), .SI(1'b0), 
        .SE(1'b0), .CK(n3538), .RN(rst_n), .Q(mult_signed_mode_ex_o[0]) );
  SDFFR_X1 mult_signed_mode_ex_o_reg_1_ ( .D(mult_signed_mode[1]), .SI(1'b0), 
        .SE(1'b0), .CK(n3538), .RN(rst_n), .Q(mult_signed_mode_ex_o[1]) );
  SDFFR_X1 mult_imm_ex_o_reg_0_ ( .D(n3532), .SI(1'b0), .SE(1'b0), .CK(n3538), 
        .RN(rst_n), .Q(mult_imm_ex_o[0]) );
  SDFFR_X1 mult_imm_ex_o_reg_1_ ( .D(n3533), .SI(1'b0), .SE(1'b0), .CK(n3538), 
        .RN(rst_n), .Q(mult_imm_ex_o[1]) );
  SDFFR_X1 mult_imm_ex_o_reg_2_ ( .D(n3534), .SI(1'b0), .SE(1'b0), .CK(n3538), 
        .RN(rst_n), .Q(mult_imm_ex_o[2]) );
  SDFFR_X1 mult_imm_ex_o_reg_3_ ( .D(n3535), .SI(1'b0), .SE(1'b0), .CK(n3538), 
        .RN(rst_n), .Q(mult_imm_ex_o[3]) );
  SDFFR_X1 mult_imm_ex_o_reg_4_ ( .D(n3536), .SI(1'b0), .SE(1'b0), .CK(n3538), 
        .RN(rst_n), .Q(mult_imm_ex_o[4]) );
  SDFFR_X1 mult_en_ex_o_reg ( .D(n2692), .SI(1'b0), .SE(1'b0), .CK(n3504), 
        .RN(rst_n), .Q(mult_en_ex_o) );
  SDFFR_X1 mult_operator_ex_o_reg_0_ ( .D(mult_operator[0]), .SI(1'b0), .SE(
        1'b0), .CK(n3479), .RN(rst_n), .Q(mult_operator_ex_o[0]) );
  SDFFR_X1 mult_operator_ex_o_reg_1_ ( .D(mult_operator[1]), .SI(1'b0), .SE(
        1'b0), .CK(n3479), .RN(rst_n), .Q(mult_operator_ex_o[1]) );
  SDFFR_X1 mult_operator_ex_o_reg_2_ ( .D(mult_operator[2]), .SI(1'b0), .SE(
        1'b0), .CK(n3479), .RN(rst_n), .Q(mult_operator_ex_o[2]) );
  SDFFR_X1 mult_is_clpx_ex_o_reg ( .D(is_clpx), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_is_clpx_ex_o) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_1_ ( .D(n2470), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[1]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_1_ ( .D(n2470), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[1]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_2_ ( .D(n2471), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[2]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_2_ ( .D(n2471), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[2]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_3_ ( .D(n2472), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[3]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_3_ ( .D(n2472), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[3]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_4_ ( .D(n2473), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[4]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_4_ ( .D(n2473), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[4]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_5_ ( .D(n2474), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[5]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_6_ ( .D(n2475), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[6]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_6_ ( .D(n2475), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[6]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_7_ ( .D(n2476), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[7]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_7_ ( .D(n2476), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[7]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_8_ ( .D(n2477), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[8]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_8_ ( .D(n2477), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[8]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_9_ ( .D(n2478), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[9]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_9_ ( .D(n2478), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[9]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_10_ ( .D(n2480), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[10]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_10_ ( .D(n2480), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[10]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_11_ ( .D(n2482), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[11]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_11_ ( .D(n2482), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[11]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_12_ ( .D(n2483), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[12]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_12_ ( .D(n2483), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[12]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_13_ ( .D(n2484), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[13]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_13_ ( .D(n2484), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[13]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_14_ ( .D(n2485), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[14]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_14_ ( .D(n2485), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[14]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_15_ ( .D(n2486), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[15]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_15_ ( .D(n2486), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[15]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_16_ ( .D(n2487), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[16]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_16_ ( .D(n2487), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[16]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_17_ ( .D(n2488), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[17]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_17_ ( .D(n2488), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[17]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_18_ ( .D(n2489), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[18]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_18_ ( .D(n2489), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[18]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_19_ ( .D(n2490), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[19]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_19_ ( .D(n2490), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[19]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_20_ ( .D(n2491), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[20]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_20_ ( .D(n2491), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[20]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_21_ ( .D(n2492), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[21]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_21_ ( .D(n2492), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[21]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_22_ ( .D(n2493), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[22]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_22_ ( .D(n2493), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[22]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_23_ ( .D(n2494), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[23]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_23_ ( .D(n2494), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[23]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_24_ ( .D(n2495), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[24]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_24_ ( .D(n2495), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[24]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_25_ ( .D(n2496), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[25]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_25_ ( .D(n2496), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[25]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_26_ ( .D(n2497), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[26]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_26_ ( .D(n2497), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[26]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_27_ ( .D(n2498), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[27]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_27_ ( .D(n2498), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[27]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_28_ ( .D(n2499), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[28]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_28_ ( .D(n2499), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[28]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_29_ ( .D(n2500), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[29]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_29_ ( .D(n2500), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[29]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_30_ ( .D(n2501), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[30]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_30_ ( .D(n2501), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[30]) );
  SDFFR_X1 mult_dot_op_c_ex_o_reg_31_ ( .D(n2502), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[31]) );
  SDFFR_X1 mult_operand_c_ex_o_reg_31_ ( .D(n2502), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[31]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_23_ ( .D(n2524), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[23]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_6_ ( .D(n3509), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[6]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_6_ ( .D(n3509), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[6]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_30_ ( .D(n2531), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[30]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_30_ ( .D(n2531), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[30]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_22_ ( .D(n2523), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[22]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_22_ ( .D(n2523), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[22]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_14_ ( .D(n2513), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[14]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_14_ ( .D(n2513), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[14]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_29_ ( .D(n2530), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[29]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_29_ ( .D(n2530), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[29]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_21_ ( .D(n3512), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[21]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_25_ ( .D(n2526), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[25]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_9_ ( .D(n3537), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[9]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_0_ ( .D(n1872), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[0]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_0_ ( .D(n1872), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[0]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_24_ ( .D(n2525), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[24]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_24_ ( .D(n2525), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[24]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_16_ ( .D(n3510), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[16]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_8_ ( .D(n2507), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[8]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_3_ ( .D(n1925), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[3]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_27_ ( .D(n2527), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[27]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_27_ ( .D(n2527), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[27]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_19_ ( .D(n2519), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[19]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_11_ ( .D(n2510), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[11]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_2_ ( .D(n1912), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[2]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_2_ ( .D(n1912), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[2]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_18_ ( .D(n2518), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[18]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_18_ ( .D(n2518), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[18]) );
  SDFFR_X1 mult_dot_op_b_ex_o_reg_10_ ( .D(n2509), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[10]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_10_ ( .D(n2509), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[10]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_0_ ( .D(n2534), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[0]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_0_ ( .D(n2534), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[0]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_31_ ( .D(n2568), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[31]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_31_ ( .D(n2568), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[31]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_30_ ( .D(n2566), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[30]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_30_ ( .D(n2566), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[30]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_28_ ( .D(n2564), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[28]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_28_ ( .D(n2564), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[28]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_27_ ( .D(n2563), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[27]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_27_ ( .D(n2563), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[27]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_26_ ( .D(n2562), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[26]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_26_ ( .D(n2562), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[26]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_25_ ( .D(n2561), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[25]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_25_ ( .D(n2561), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[25]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_24_ ( .D(n2560), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[24]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_24_ ( .D(n2560), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[24]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_23_ ( .D(n2559), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[23]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_23_ ( .D(n2559), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[23]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_22_ ( .D(n2558), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[22]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_22_ ( .D(n2558), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[22]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_21_ ( .D(n2557), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[21]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_21_ ( .D(n2557), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[21]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_20_ ( .D(n2556), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[20]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_20_ ( .D(n2556), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[20]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_19_ ( .D(n2555), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[19]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_19_ ( .D(n2555), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[19]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_18_ ( .D(n2554), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[18]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_18_ ( .D(n2554), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[18]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_17_ ( .D(n2553), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[17]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_17_ ( .D(n2553), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[17]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_16_ ( .D(n2552), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[16]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_16_ ( .D(n2552), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[16]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_15_ ( .D(n2550), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[15]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_15_ ( .D(n2550), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[15]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_1_ ( .D(n2535), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[1]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_14_ ( .D(n2549), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[14]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_14_ ( .D(n2549), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[14]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_13_ ( .D(n2548), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[13]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_13_ ( .D(n2548), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[13]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_12_ ( .D(n2547), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[12]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_11_ ( .D(n2546), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[11]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_11_ ( .D(n2546), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[11]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_10_ ( .D(n2545), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[10]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_10_ ( .D(n2545), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[10]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_9_ ( .D(n2544), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[9]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_9_ ( .D(n2544), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[9]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_8_ ( .D(n2543), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[8]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_7_ ( .D(n2542), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[7]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_7_ ( .D(n2542), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[7]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_6_ ( .D(n2541), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[6]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_5_ ( .D(n2540), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[5]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_5_ ( .D(n2540), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[5]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_4_ ( .D(n2539), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[4]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_4_ ( .D(n2539), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[4]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_3_ ( .D(n2538), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[3]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_3_ ( .D(n2538), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[3]) );
  SDFFR_X1 mult_operand_a_ex_o_reg_2_ ( .D(n2536), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[2]) );
  SDFFR_X1 alu_operator_ex_o_reg_2_ ( .D(n3489), .SI(1'b0), .SE(1'b0), .CK(
        n3496), .RN(rst_n), .Q(alu_operator_ex_o[2]) );
  SDFFR_X1 alu_operator_ex_o_reg_3_ ( .D(n3490), .SI(1'b0), .SE(1'b0), .CK(
        n3496), .RN(rst_n), .Q(alu_operator_ex_o[3]) );
  SDFFR_X1 alu_operator_ex_o_reg_4_ ( .D(n3491), .SI(1'b0), .SE(1'b0), .CK(
        n3496), .RN(rst_n), .Q(alu_operator_ex_o[4]) );
  SDFFR_X1 alu_operator_ex_o_reg_5_ ( .D(n3492), .SI(1'b0), .SE(1'b0), .CK(
        n3496), .RN(rst_n), .Q(alu_operator_ex_o[5]) );
  SDFFR_X1 alu_en_ex_o_reg ( .D(n3502), .SI(1'b0), .SE(1'b0), .CK(n3504), .RN(
        rst_n), .QN(alu_en_ex_o_BAR) );
  SDFFR_X1 alu_clpx_shift_ex_o_reg_0_ ( .D(instr_rdata_i[13]), .SI(1'b0), .SE(
        1'b0), .CK(n3530), .RN(rst_n), .Q(alu_clpx_shift_ex_o[0]) );
  SDFFR_X1 alu_is_subrot_ex_o_reg ( .D(is_subrot), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_is_subrot_ex_o) );
  SDFFR_X1 alu_is_clpx_ex_o_reg ( .D(is_clpx), .SI(1'b0), .SE(1'b0), .CK(n3530), .RN(rst_n), .Q(alu_is_clpx_ex_o) );
  SDFFR_X1 alu_vec_mode_ex_o_reg_0_ ( .D(alu_vec_mode[0]), .SI(1'b0), .SE(1'b0), .CK(n3530), .RN(rst_n), .Q(alu_vec_mode_ex_o[0]) );
  SDFFR_X1 imm_vec_ext_ex_o_reg_1_ ( .D(instr_rdata_i[20]), .SI(1'b0), .SE(
        1'b0), .CK(n3530), .RN(rst_n), .Q(imm_vec_ext_ex_o[1]) );
  SDFFR_X1 imm_vec_ext_ex_o_reg_0_ ( .D(instr_rdata_i[25]), .SI(1'b0), .SE(
        1'b0), .CK(n3530), .RN(rst_n), .Q(imm_vec_ext_ex_o[0]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_31_ ( .D(n2502), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[31]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_30_ ( .D(n2501), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[30]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_29_ ( .D(n2500), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[29]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_28_ ( .D(n2499), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[28]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_27_ ( .D(n2498), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[27]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_26_ ( .D(n2497), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[26]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_25_ ( .D(n2496), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[25]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_24_ ( .D(n2495), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[24]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_23_ ( .D(n2494), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[23]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_22_ ( .D(n2493), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[22]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_21_ ( .D(n2492), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[21]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_20_ ( .D(n2491), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[20]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_19_ ( .D(n2490), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[19]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_17_ ( .D(n2488), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[17]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_16_ ( .D(n2487), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[16]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_15_ ( .D(n2486), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[15]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_13_ ( .D(n2484), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[13]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_12_ ( .D(n2483), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[12]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_11_ ( .D(n2482), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[11]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_10_ ( .D(n2480), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[10]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_9_ ( .D(n2478), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[9]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_8_ ( .D(n2477), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[8]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_7_ ( .D(n2476), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[7]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_6_ ( .D(n2475), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[6]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_5_ ( .D(n2474), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[5]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_4_ ( .D(n2473), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[4]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_3_ ( .D(n2472), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[3]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_2_ ( .D(n2471), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[2]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_1_ ( .D(n2470), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[1]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_0_ ( .D(n1872), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[0]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_30_ ( .D(n2531), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[30]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_29_ ( .D(n2530), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[29]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_27_ ( .D(n2527), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[27]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_22_ ( .D(n2523), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[22]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_14_ ( .D(n2513), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[14]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_13_ ( .D(n2512), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[13]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_11_ ( .D(n2510), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[11]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_6_ ( .D(n3509), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[6]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_3_ ( .D(n1925), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[3]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_2_ ( .D(n1912), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[2]) );
  SDFFR_X1 alu_operand_a_ex_o_reg_0_ ( .D(n2534), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[0]) );
  SDFFR_X1 alu_operand_a_ex_o_reg_6_ ( .D(n2541), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[6]) );
  SDFFR_X1 bmask_b_ex_o_reg_0_ ( .D(n3520), .SI(1'b0), .SE(1'b0), .CK(n3530), 
        .RN(rst_n), .Q(bmask_b_ex_o[0]) );
  SDFFR_X1 bmask_b_ex_o_reg_1_ ( .D(n3521), .SI(1'b0), .SE(1'b0), .CK(n3530), 
        .RN(rst_n), .Q(bmask_b_ex_o[1]) );
  SDFFR_X1 bmask_b_ex_o_reg_2_ ( .D(n3522), .SI(1'b0), .SE(1'b0), .CK(n3530), 
        .RN(rst_n), .Q(bmask_b_ex_o[2]) );
  SDFFR_X1 bmask_b_ex_o_reg_3_ ( .D(n3523), .SI(1'b0), .SE(1'b0), .CK(n3530), 
        .RN(rst_n), .Q(bmask_b_ex_o[3]) );
  SDFFR_X1 bmask_b_ex_o_reg_4_ ( .D(n3524), .SI(1'b0), .SE(1'b0), .CK(n3530), 
        .RN(rst_n), .Q(bmask_b_ex_o[4]) );
  SDFFR_X1 bmask_a_ex_o_reg_0_ ( .D(n3525), .SI(1'b0), .SE(1'b0), .CK(n3530), 
        .RN(rst_n), .Q(bmask_a_ex_o[0]) );
  SDFFR_X1 bmask_a_ex_o_reg_1_ ( .D(n3526), .SI(1'b0), .SE(1'b0), .CK(n3530), 
        .RN(rst_n), .Q(bmask_a_ex_o[1]) );
  SDFFR_X1 bmask_a_ex_o_reg_2_ ( .D(n3527), .SI(1'b0), .SE(1'b0), .CK(n3530), 
        .RN(rst_n), .Q(bmask_a_ex_o[2]) );
  SDFFR_X1 bmask_a_ex_o_reg_3_ ( .D(n3528), .SI(1'b0), .SE(1'b0), .CK(n3530), 
        .RN(rst_n), .Q(bmask_a_ex_o[3]) );
  SDFFR_X1 bmask_a_ex_o_reg_4_ ( .D(n3529), .SI(1'b0), .SE(1'b0), .CK(n3530), 
        .RN(rst_n), .Q(bmask_a_ex_o[4]) );
  SDFFR_X1 data_load_event_ex_o_reg ( .D(n3503), .SI(1'b0), .SE(1'b0), .CK(
        n3504), .RN(rst_n), .Q(data_load_event_ex_o) );
  SDFFR_X1 data_misaligned_ex_o_reg ( .D(n1276), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(rst_n), .QN(n2597) );
  SDFFR_X1 pc_ex_o_reg_31_ ( .D(pc_id_i[31]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[31]) );
  SDFFR_X1 pc_ex_o_reg_30_ ( .D(pc_id_i[30]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[30]) );
  SDFFR_X1 pc_ex_o_reg_29_ ( .D(pc_id_i[29]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[29]) );
  SDFFR_X1 pc_ex_o_reg_28_ ( .D(pc_id_i[28]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[28]) );
  SDFFR_X1 pc_ex_o_reg_27_ ( .D(pc_id_i[27]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[27]) );
  SDFFR_X1 pc_ex_o_reg_26_ ( .D(pc_id_i[26]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[26]) );
  SDFFR_X1 pc_ex_o_reg_25_ ( .D(pc_id_i[25]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[25]) );
  SDFFR_X1 pc_ex_o_reg_24_ ( .D(pc_id_i[24]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[24]) );
  SDFFR_X1 pc_ex_o_reg_23_ ( .D(pc_id_i[23]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[23]) );
  SDFFR_X1 pc_ex_o_reg_22_ ( .D(pc_id_i[22]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[22]) );
  SDFFR_X1 pc_ex_o_reg_21_ ( .D(pc_id_i[21]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[21]) );
  SDFFR_X1 pc_ex_o_reg_20_ ( .D(pc_id_i[20]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[20]) );
  SDFFR_X1 pc_ex_o_reg_19_ ( .D(pc_id_i[19]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[19]) );
  SDFFR_X1 pc_ex_o_reg_18_ ( .D(pc_id_i[18]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[18]) );
  SDFFR_X1 pc_ex_o_reg_17_ ( .D(pc_id_i[17]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[17]) );
  SDFFR_X1 pc_ex_o_reg_16_ ( .D(pc_id_i[16]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[16]) );
  SDFFR_X1 pc_ex_o_reg_15_ ( .D(pc_id_i[15]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[15]) );
  SDFFR_X1 pc_ex_o_reg_14_ ( .D(pc_id_i[14]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[14]) );
  SDFFR_X1 pc_ex_o_reg_13_ ( .D(pc_id_i[13]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[13]) );
  SDFFR_X1 pc_ex_o_reg_12_ ( .D(pc_id_i[12]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[12]) );
  SDFFR_X1 pc_ex_o_reg_11_ ( .D(pc_id_i[11]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[11]) );
  SDFFR_X1 pc_ex_o_reg_10_ ( .D(pc_id_i[10]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[10]) );
  SDFFR_X1 pc_ex_o_reg_9_ ( .D(pc_id_i[9]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[9]) );
  SDFFR_X1 pc_ex_o_reg_8_ ( .D(pc_id_i[8]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[8]) );
  SDFFR_X1 pc_ex_o_reg_7_ ( .D(pc_id_i[7]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[7]) );
  SDFFR_X1 pc_ex_o_reg_6_ ( .D(pc_id_i[6]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[6]) );
  SDFFR_X1 pc_ex_o_reg_5_ ( .D(pc_id_i[5]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[5]) );
  SDFFR_X1 pc_ex_o_reg_4_ ( .D(pc_id_i[4]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[4]) );
  SDFFR_X1 pc_ex_o_reg_3_ ( .D(pc_id_i[3]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[3]) );
  SDFFR_X1 pc_ex_o_reg_2_ ( .D(pc_id_i[2]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[2]) );
  SDFFR_X1 pc_ex_o_reg_1_ ( .D(pc_id_i[1]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[1]) );
  SDFFR_X1 pc_ex_o_reg_0_ ( .D(pc_id_i[0]), .SI(1'b0), .SE(1'b0), .CK(n3518), 
        .RN(rst_n), .Q(pc_ex_o[0]) );
  SDFFR_X1 alu_operator_ex_o_reg_6_ ( .D(n3493), .SI(1'b0), .SE(1'b0), .CK(
        n3496), .RN(rst_n), .Q(alu_operator_ex_o[6]) );
  SDFFS_X1 alu_operator_ex_o_reg_0_ ( .D(n3494), .SI(1'b0), .SE(1'b0), .CK(
        n3496), .SN(rst_n), .Q(alu_operator_ex_o[0]) );
  SDFFR_X1 alu_operand_a_ex_o_reg_10_ ( .D(n2545), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[10]) );
  SDFFR_X1 alu_operand_a_ex_o_reg_18_ ( .D(n2554), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[18]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_31_ ( .D(n150), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[31]) );
  SDFFR_X1 alu_operand_a_ex_o_reg_13_ ( .D(n2548), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[13]) );
  SDFFS_X1 alu_operand_b_ex_o_reg_9_ ( .D(n2508), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .SN(rst_n), .QN(alu_operand_b_ex_o[9]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_18_ ( .D(n3511), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[18]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_8_ ( .D(n2507), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[8]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_2_ ( .D(n2536), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[2]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_1_ ( .D(n2535), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[1]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_12_ ( .D(n2547), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[12]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_21_ ( .D(n3512), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[21]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_15_ ( .D(n2514), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[15]) );
  SDFFR_X1 alu_operand_a_ex_o_reg_3_ ( .D(n2538), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[3]) );
  SDFFR_X1 alu_operand_a_ex_o_reg_14_ ( .D(n2549), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[14]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_24_ ( .D(n2525), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[24]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_26_ ( .D(n162), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[26]) );
  SDFFR_X1 alu_operand_a_ex_o_reg_12_ ( .D(n2547), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[12]) );
  SDFFR_X1 alu_operand_a_ex_o_reg_8_ ( .D(n2543), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[8]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_6_ ( .D(n2541), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[6]) );
  SDFFR_X1 mult_dot_op_a_ex_o_reg_8_ ( .D(n2543), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[8]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_18_ ( .D(n2489), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[18]) );
  SDFFR_X1 alu_operand_c_ex_o_reg_14_ ( .D(n2485), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[14]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_9_ ( .D(n2544), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[9]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_16_ ( .D(n2552), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[16]) );
  SDFFR_X2 alu_operand_b_ex_o_reg_16_ ( .D(n3510), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[16]) );
  SDFFR_X2 alu_operand_b_ex_o_reg_21_ ( .D(n3512), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[21]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_7_ ( .D(n2542), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[7]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_23_ ( .D(n2559), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[23]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_26_ ( .D(n2562), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[26]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_5_ ( .D(n2540), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[5]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_4_ ( .D(n2539), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[4]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_20_ ( .D(n2556), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[20]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_25_ ( .D(n2561), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[25]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_31_ ( .D(n2568), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[31]) );
  register_file_test_wrap_ADDR_WIDTH6_FPU0_Zfinx0 registers_i ( .clk(clk), 
        .rst_n(rst_n), .test_en_i(1'b0), .raddr_a_i({1'b0, 
        instr_rdata_i[19:15]}), .rdata_a_o({regfile_data_ra_id[31:22], n2644, 
        regfile_data_ra_id[20:11], n47, regfile_data_ra_id[9:0]}), .raddr_b_i(
        {1'b0, n2604, instr_rdata_i[23:20]}), .rdata_b_o(regfile_data_rb_id), 
        .raddr_c_i({1'b0, n1638, n1637, n1636, n1635, n1634}), .rdata_c_o(
        regfile_data_rc_id), .waddr_a_i({1'b0, regfile_waddr_wb_i[4:0]}), 
        .wdata_a_i(regfile_wdata_wb_i), .we_a_i(regfile_we_wb_i), .waddr_b_i({
        1'b0, regfile_alu_waddr_fw_i[4:0]}), .wdata_b_i({
        regfile_alu_wdata_fw_i[31:29], n2667, regfile_alu_wdata_fw_i[27:0]}), 
        .we_b_i(regfile_alu_we_fw_i), .BIST(1'b0), .CSN_T(1'b0), .WEN_T(1'b0), 
        .A_T({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D_T({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  riscv_decoder_FPU0_FP_DIVSQRT0_PULP_SECURE1_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_WOP_CPU6 decoder_i ( 
        .deassert_we_i(deassert_we), .data_misaligned_i(data_misaligned_i), 
        .mult_multicycle_i(mult_multicycle_i), .illegal_insn_o(
        illegal_insn_dec), .ebrk_insn_o(n2645), .mret_insn_o(mret_insn_dec), 
        .uret_insn_o(uret_insn_dec), .dret_insn_o(dret_insn_dec), .mret_dec_o(
        mret_dec), .dret_dec_o(dret_dec), .ecall_insn_o(ecall_insn_dec), 
        .pipe_flush_o(pipe_flush_dec), .fencei_insn_o(fencei_insn_dec), 
        .rega_used_o(rega_used_dec), .regb_used_o(regb_used_dec), 
        .regc_used_o(regc_used_dec), .bmask_a_mux_o(bmask_a_mux_0_), 
        .bmask_b_mux_o(bmask_b_mux), .alu_bmask_a_mux_sel_o(
        alu_bmask_a_mux_sel), .alu_bmask_b_mux_sel_o(alu_bmask_b_mux_sel), 
        .instr_rdata_i({instr_rdata_i[31:25], n2604, instr_rdata_i[23:20], 
        n116, n33, n110, n80, n113, instr_rdata_i[14:0]}), .illegal_c_insn_i(
        illegal_c_insn_i), .alu_en_o(alu_en), .alu_operator_o(alu_operator), 
        .alu_op_a_mux_sel_o(alu_op_a_mux_sel), .alu_op_b_mux_sel_o(
        alu_op_b_mux_sel), .alu_op_c_mux_sel_o(alu_op_c_mux_sel), 
        .alu_vec_mode_o(alu_vec_mode), .scalar_replication_o(
        scalar_replication), .imm_a_mux_sel_o(imm_a_mux_sel_0_), 
        .imm_b_mux_sel_o(imm_b_mux_sel), .regc_mux_o(regc_mux), .is_clpx_o(
        is_clpx), .is_subrot_o(is_subrot), .mult_operator_o(mult_operator), 
        .mult_int_en_o(mult_int_en), .mult_dot_en_o(mult_dot_en), 
        .mult_sel_subword_o(mult_sel_subword), .mult_signed_mode_o(
        mult_signed_mode), .mult_dot_signed_o(mult_dot_signed), .frm_i({1'b0, 
        1'b0, 1'b0}), .regfile_mem_we_o(regfile_we_id), .regfile_alu_we_o(
        regfile_alu_we_id), .regfile_alu_we_dec_o(regfile_alu_we_dec_id), 
        .regfile_alu_waddr_sel_o(regfile_alu_waddr_mux_sel), .csr_access_o(
        csr_access), .csr_status_o(csr_status), .csr_op_o(csr_op), 
        .current_priv_lvl_i(current_priv_lvl_i), .data_req_o(data_req_id), 
        .data_we_o(data_we_id), .prepost_useincr_o(prepost_useincr), 
        .data_type_o(data_type_id), .data_sign_extension_o({
        SYNOPSYS_UNCONNECTED__0, data_sign_ext_id_0_}), .data_load_event_o(
        data_load_event_id), .hwloop_we_o(hwloop_we_int), 
        .hwloop_target_mux_sel_o(n2631), .hwloop_start_mux_sel_o(
        hwloop_start_mux_sel), .hwloop_cnt_mux_sel_o(hwloop_cnt_mux_sel), 
        .jump_in_dec_o(jump_in_dec), .jump_in_id_o(jump_in_id), 
        .jump_target_mux_sel_o(jump_target_mux_sel), .\mult_imm_mux_o[0]_BAR (
        mult_imm_mux_0_) );
  riscv_controller_FPU0 controller_i ( .clk(clk), .rst_n(rst_n), 
        .fetch_enable_i(fetch_enable_i), .ctrl_busy_o(ctrl_busy_o), 
        .first_fetch_o(core_ctrl_firstfetch_o), .is_fetch_failed_i(1'b0), 
        .deassert_we_o(deassert_we), .illegal_insn_i(illegal_insn_dec), 
        .ecall_insn_i(ecall_insn_dec), .mret_insn_i(mret_insn_dec), 
        .uret_insn_i(uret_insn_dec), .dret_insn_i(dret_insn_dec), .mret_dec_i(
        mret_dec), .uret_dec_i(1'b0), .dret_dec_i(dret_dec), .pipe_flush_i(
        pipe_flush_dec), .ebrk_insn_i(n2645), .fencei_insn_i(fencei_insn_dec), 
        .csr_status_i(csr_status), .instr_multicycle_i(1'b0), .instr_valid_i(
        instr_valid_i), .instr_req_o(instr_req_o), .pc_set_o(pc_set_o), 
        .pc_mux_o(pc_mux_o), .exc_pc_mux_o({SYNOPSYS_UNCONNECTED__1, 
        exc_pc_mux_o[1:0]}), .trap_addr_mux_o(trap_addr_mux_o), 
        .data_req_ex_i(data_req_ex_o), .data_we_ex_i(data_we_ex_o), 
        .data_misaligned_i(data_misaligned_i), .data_load_event_i(
        data_load_event_id), .mult_multicycle_i(mult_multicycle_i), .apu_en_i(
        1'b0), .apu_read_dep_i(1'b0), .apu_write_dep_i(1'b0), 
        .branch_taken_ex_i(branch_taken_ex), .jump_in_id_i(jump_in_id), 
        .jump_in_dec_i(jump_in_dec), .irq_i(irq_i), .irq_req_ctrl_i(
        irq_req_ctrl), .irq_sec_ctrl_i(irq_sec_ctrl), .irq_id_ctrl_i(
        irq_id_ctrl), .m_IE_i(m_irq_enable_i), .u_IE_i(u_irq_enable_i), 
        .current_priv_lvl_i(current_priv_lvl_i), .irq_id_o(irq_id_o), 
        .exc_cause_o({SYNOPSYS_UNCONNECTED__2, exc_cause_o[4:0]}), 
        .exc_kill_o(exc_kill), .debug_cause_o({debug_cause_o[2:1], 
        SYNOPSYS_UNCONNECTED__3}), .debug_csr_save_o(debug_csr_save_o), 
        .debug_req_i(debug_req_i), .debug_single_step_i(debug_single_step_i), 
        .debug_ebreakm_i(debug_ebreakm_i), .debug_ebreaku_i(debug_ebreaku_i), 
        .csr_save_if_o(csr_save_if_o), .csr_save_id_o(csr_save_id_o), 
        .csr_irq_sec_o(csr_irq_sec_o), .csr_restore_mret_id_o(
        csr_restore_mret_id_o), .csr_restore_uret_id_o(csr_restore_uret_id_o), 
        .csr_restore_dret_id_o(csr_restore_dret_id_o), .csr_save_cause_o(
        csr_save_cause_o), .regfile_we_id_i(regfile_alu_we_dec_id), 
        .regfile_alu_waddr_id_i({1'b0, regfile_alu_waddr_id}), 
        .regfile_we_ex_i(regfile_we_ex_o), .regfile_waddr_ex_i({1'b0, 
        regfile_waddr_ex_o[4:0]}), .regfile_we_wb_i(regfile_we_wb_i), 
        .regfile_alu_we_fw_i(regfile_alu_we_fw_i), .operand_a_fw_mux_sel_o(
        operand_a_fw_mux_sel), .operand_b_fw_mux_sel_o(operand_b_fw_mux_sel), 
        .reg_d_ex_is_reg_a_i(reg_d_ex_is_reg_a_id), .reg_d_ex_is_reg_b_i(
        reg_d_ex_is_reg_b_id), .reg_d_ex_is_reg_c_i(reg_d_ex_is_reg_c_id), 
        .reg_d_wb_is_reg_a_i(reg_d_wb_is_reg_a_id), .reg_d_wb_is_reg_b_i(
        reg_d_wb_is_reg_b_id), .reg_d_wb_is_reg_c_i(reg_d_wb_is_reg_c_id), 
        .reg_d_alu_is_reg_a_i(reg_d_alu_is_reg_a_id), .reg_d_alu_is_reg_b_i(
        reg_d_alu_is_reg_b_id), .reg_d_alu_is_reg_c_i(reg_d_alu_is_reg_c_id), 
        .halt_if_o(halt_if_o), .jr_stall_o(jr_stall), .load_stall_o(load_stall), .ex_valid_i(ex_valid_i), .wb_ready_i(wb_ready_i), .perf_jump_o(perf_jump_o), 
        .perf_jr_stall_o(perf_jr_stall_o), .perf_ld_stall_o(perf_ld_stall_o), 
        .perf_pipeline_stall_o(perf_pipeline_stall_o), .irq_ack_o_BAR(
        irq_ack_o_BAR), .exc_ack_o_BAR(exc_ack), .csr_cause_o_5__BAR(
        csr_cause_o_5__BAR), .csr_cause_o_4_(csr_cause_o_4_), .csr_cause_o_3_(
        csr_cause_o_3_), .csr_cause_o_2_(csr_cause_o_2_), .csr_cause_o_0_(
        csr_cause_o_0_), .id_ready_i_BAR(n2577), .data_err_ack_o_BAR(
        data_err_ack_o_BAR), .csr_save_ex_o_BAR(csr_save_ex_o_BAR), 
        .data_err_i_BAR(data_err_i_BAR), .csr_cause_o_1__BAR(
        csr_cause_o_1__BAR), .halt_id_o_BAR(n55), .operand_c_fw_mux_sel_o_1_(
        operand_c_fw_mux_sel[1]), .operand_c_fw_mux_sel_o_0__BAR(
        operand_c_fw_mux_sel[0]), .is_decoding_o(is_decoding_o_BAR) );
  riscv_int_controller_PULP_SECURE1 int_controller_i ( .clk(clk), .rst_n(rst_n), .irq_req_ctrl_o(irq_req_ctrl), .irq_sec_ctrl_o(irq_sec_ctrl), 
        .irq_id_ctrl_o(irq_id_ctrl), .ctrl_kill_i(exc_kill), .irq_i(irq_i), 
        .irq_sec_i(irq_sec_i), .irq_id_i(irq_id_i), .m_IE_i(m_irq_enable_i), 
        .u_IE_i(u_irq_enable_i), .current_priv_lvl_i(current_priv_lvl_i), 
        .ctrl_ack_i_BAR(exc_ack) );
  riscv_hwloop_regs_N_REGS2 hwloop_regs_i ( .clk(clk), .rst_n(rst_n), 
        .hwlp_start_data_i(hwloop_start), .hwlp_end_data_i(hwloop_end), 
        .hwlp_cnt_data_i(hwloop_cnt), .hwlp_we_i(hwloop_we), .hwlp_regid_i(
        hwloop_regid_0_), .valid_i(hwloop_valid), .hwlp_dec_cnt_i(
        hwlp_dec_cnt_i), .hwlp_start_addr_o(hwlp_start_o), .hwlp_end_addr_o(
        hwlp_end_o), .hwlp_counter_o(hwlp_cnt_o) );
  SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_0 clk_gate_mult_dot_op_a_ex_o_reg_8_ ( 
        .CLK(clk), .EN(n2652), .ENCLK(n3540), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_1 clk_gate_mult_operand_b_ex_o_reg_15_ ( 
        .CLK(clk), .EN(n2650), .ENCLK(n3538), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_2 clk_gate_alu_operand_c_ex_o_reg_14_ ( 
        .CLK(clk), .EN(n778), .ENCLK(n3530), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_3 clk_gate_pc_ex_o_reg_0_ ( 
        .CLK(clk), .EN(n2571), .ENCLK(n3518), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_4 clk_gate_mult_operand_c_ex_o_reg_31_ ( 
        .CLK(clk), .EN(n3517), .ENCLK(n3515), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_5 clk_gate_alu_operand_b_ex_o_reg_26_ ( 
        .CLK(clk), .EN(n2533), .ENCLK(n3513), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_6 clk_gate_alu_operand_a_ex_o_reg_8_ ( 
        .CLK(clk), .EN(n2694), .ENCLK(n3507), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_7 clk_gate_data_load_event_ex_o_reg ( 
        .CLK(clk), .EN(n3506), .ENCLK(n3504), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_8 clk_gate_alu_operator_ex_o_reg_1_ ( 
        .CLK(clk), .EN(n3498), .ENCLK(n3496), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_9 clk_gate_regfile_waddr_ex_o_reg_4_ ( 
        .CLK(clk), .EN(n2693), .ENCLK(n3487), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_10 clk_gate_regfile_alu_waddr_ex_o_reg_4_ ( 
        .CLK(clk), .EN(n3486), .ENCLK(n3484), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_11 clk_gate_data_sign_ext_ex_o_reg_0_ ( 
        .CLK(clk), .EN(n3483), .ENCLK(n3481), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5_12 clk_gate_mult_operator_ex_o_reg_2_ ( 
        .CLK(clk), .EN(n2692), .ENCLK(n3479), .TE(1'b0) );
  SDFFR_X2 csr_access_ex_o_reg ( .D(n1626), .SI(1'b0), .SE(1'b0), .CK(n3504), 
        .RN(rst_n), .Q(csr_access_ex_o), .QN(csr_access_ex_o_BAR) );
  SDFFR_X2 alu_operand_a_ex_o_reg_24_ ( .D(n2560), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[24]) );
  SDFFR_X2 alu_operand_b_ex_o_reg_10_ ( .D(n2509), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[10]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_19_ ( .D(n2555), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[19]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_17_ ( .D(n2553), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[17]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_2_ ( .D(n2536), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[2]) );
  SDFFR_X2 alu_operand_b_ex_o_reg_28_ ( .D(n2528), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[28]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_28_ ( .D(n2528), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[28]) );
  SDFFR_X2 mult_operand_b_ex_o_reg_28_ ( .D(n2528), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[28]) );
  SDFFR_X2 alu_operand_b_ex_o_reg_25_ ( .D(n2526), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[25]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_25_ ( .D(n2526), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[25]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_31_ ( .D(n150), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[31]) );
  SDFFR_X2 mult_operand_b_ex_o_reg_31_ ( .D(n150), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[31]) );
  SDFFR_X2 alu_operand_b_ex_o_reg_15_ ( .D(n2514), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[15]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_15_ ( .D(n2514), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[15]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_9_ ( .D(n3537), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[9]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_12_ ( .D(n2511), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[12]) );
  SDFFR_X2 mult_operand_b_ex_o_reg_12_ ( .D(n2511), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[12]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_26_ ( .D(n162), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[26]) );
  SDFFR_X2 mult_operand_b_ex_o_reg_26_ ( .D(n162), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[26]) );
  SDFFR_X2 alu_operand_b_ex_o_reg_20_ ( .D(n2520), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[20]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_20_ ( .D(n2520), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[20]) );
  SDFFR_X2 mult_operand_b_ex_o_reg_20_ ( .D(n2520), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[20]) );
  SDFFR_X2 alu_operand_b_ex_o_reg_23_ ( .D(n2524), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[23]) );
  SDFFR_X2 mult_operand_b_ex_o_reg_23_ ( .D(n2524), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[23]) );
  SDFFR_X2 alu_operand_b_ex_o_reg_19_ ( .D(n2519), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[19]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_21_ ( .D(n2557), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[21]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_27_ ( .D(n2563), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[27]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_1_ ( .D(n2535), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[1]) );
  SDFFR_X2 alu_operand_b_ex_o_reg_1_ ( .D(n1874), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[1]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_11_ ( .D(n2546), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[11]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_15_ ( .D(n2550), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[15]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_22_ ( .D(n2558), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[22]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_30_ ( .D(n2566), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[30]) );
  SDFFR_X2 alu_vec_mode_ex_o_reg_1_ ( .D(alu_vec_mode[1]), .SI(1'b0), .SE(1'b0), .CK(n3530), .RN(rst_n), .Q(alu_vec_mode_ex_o[1]) );
  SDFFR_X2 mult_dot_op_c_ex_o_reg_5_ ( .D(n2474), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[5]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_8_ ( .D(n2507), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[8]) );
  SDFFR_X2 mult_operand_b_ex_o_reg_17_ ( .D(n2517), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[17]) );
  SDFFR_X2 mult_operand_b_ex_o_reg_19_ ( .D(n2519), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[19]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_28_ ( .D(n2564), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[28]) );
  SDFFR_X2 mult_operand_b_ex_o_reg_7_ ( .D(n2506), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[7]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_7_ ( .D(n2506), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[7]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_7_ ( .D(n2506), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[7]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_17_ ( .D(n2666), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[17]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_17_ ( .D(n2517), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[17]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_1_ ( .D(n1874), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[1]) );
  SDFFR_X1 alu_operand_b_ex_o_reg_12_ ( .D(n2511), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[12]) );
  SDFFR_X2 alu_operand_b_ex_o_reg_5_ ( .D(n2661), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[5]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_5_ ( .D(n2661), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[5]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_4_ ( .D(n1940), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[4]) );
  SDFFR_X2 mult_operand_b_ex_o_reg_4_ ( .D(n1940), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[4]) );
  SDFFR_X2 alu_operand_b_ex_o_reg_4_ ( .D(n1940), .SI(1'b0), .SE(1'b0), .CK(
        n3513), .RN(rst_n), .Q(alu_operand_b_ex_o[4]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_13_ ( .D(n2512), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[13]) );
  SDFFR_X2 mult_operand_b_ex_o_reg_13_ ( .D(n2512), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[13]) );
  SDFFR_X2 mult_dot_op_a_ex_o_reg_29_ ( .D(n2565), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_a_ex_o[29]) );
  SDFFR_X2 mult_operand_a_ex_o_reg_29_ ( .D(n2565), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_a_ex_o[29]) );
  SDFFR_X2 alu_operand_a_ex_o_reg_29_ ( .D(n2565), .SI(1'b0), .SE(1'b0), .CK(
        n3507), .RN(rst_n), .Q(alu_operand_a_ex_o[29]) );
  SDFFR_X2 mult_clpx_shift_ex_o_reg_1_ ( .D(instr_rdata_i[14]), .SI(1'b0), 
        .SE(1'b0), .CK(n3540), .RN(rst_n), .Q(mult_clpx_shift_ex_o[1]) );
  SDFFR_X2 alu_clpx_shift_ex_o_reg_1_ ( .D(instr_rdata_i[14]), .SI(1'b0), .SE(
        1'b0), .CK(n3530), .RN(rst_n), .Q(alu_clpx_shift_ex_o[1]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_3_ ( .D(n1925), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[3]) );
  SDFFR_X2 mult_dot_op_b_ex_o_reg_11_ ( .D(n2510), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_b_ex_o[11]) );
  SDFFR_X2 mult_dot_op_c_ex_o_reg_0_ ( .D(n2469), .SI(1'b0), .SE(1'b0), .CK(
        n3540), .RN(rst_n), .Q(mult_dot_op_c_ex_o[0]) );
  SDFFR_X2 mult_operand_c_ex_o_reg_0_ ( .D(n2469), .SI(1'b0), .SE(1'b0), .CK(
        n3515), .RN(rst_n), .Q(mult_operand_c_ex_o[0]) );
  SDFFR_X2 alu_operand_c_ex_o_reg_0_ ( .D(n2656), .SI(1'b0), .SE(1'b0), .CK(
        n3530), .RN(rst_n), .Q(alu_operand_c_ex_o[0]) );
  INV_X1 U383 ( .A(n292), .ZN(n277) );
  OAI21_X1 U25 ( .B1(n528), .B2(n597), .A(n529), .ZN(n521) );
  OAI211_X1 U64 ( .C1(n743), .C2(n2430), .A(n732), .B(n731), .ZN(n1635) );
  AND2_X1 U99 ( .A1(n602), .A2(operand_b_fw_mux_sel[1]), .ZN(n2207) );
  OR2_X1 U97 ( .A1(n2140), .A2(n2219), .ZN(n2299) );
  NAND2_X1 U14 ( .A1(n1125), .A2(n1073), .ZN(n1160) );
  INV_X2 U763 ( .A(hwloop_we_int[1]), .ZN(n854) );
  INV_X1 U63 ( .A(n854), .ZN(n860) );
  OR2_X1 U93 ( .A1(n719), .A2(n1884), .ZN(n814) );
  INV_X1 U378 ( .A(n211), .ZN(n1005) );
  AND2_X2 U72 ( .A1(n1005), .A2(hwloop_start_mux_sel), .ZN(n900) );
  BUF_X1 U77 ( .A(instr_rdata_i[16]), .Z(n80) );
  SDFFR_X2 alu_operator_ex_o_reg_1_ ( .D(n3495), .SI(1'b0), .SE(1'b0), .CK(
        n3496), .RN(rst_n), .QN(alu_operator_ex_o[1]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_1_ ( .D(n1874), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[1]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_16_ ( .D(n3510), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[16]) );
  SDFFR_X1 mult_operand_b_ex_o_reg_5_ ( .D(n2662), .SI(1'b0), .SE(1'b0), .CK(
        n3538), .RN(rst_n), .Q(mult_operand_b_ex_o[5]) );
  CLKBUF_X1 U3 ( .A(regfile_data_ra_id[2]), .Z(n2627) );
  BUF_X1 U4 ( .A(n272), .Z(n2673) );
  BUF_X1 U5 ( .A(instr_rdata_i[17]), .Z(n110) );
  BUF_X1 U6 ( .A(n1647), .Z(n2147) );
  BUF_X2 U7 ( .A(regfile_alu_wdata_fw_i[28]), .Z(n2667) );
  CLKBUF_X1 U8 ( .A(ex_ready_i), .Z(n2671) );
  CLKBUF_X2 U9 ( .A(n995), .Z(n1000) );
  CLKBUF_X2 U10 ( .A(n318), .Z(n48) );
  BUF_X2 U11 ( .A(jump_target_mux_sel[0]), .Z(n90) );
  CLKBUF_X1 U12 ( .A(instr_rdata_i[27]), .Z(n2678) );
  OAI21_X1 U13 ( .B1(n2188), .B2(n1881), .A(n1731), .ZN(n2506) );
  OR2_X1 U20 ( .A1(n605), .A2(n185), .ZN(n638) );
  OR2_X1 U21 ( .A1(n2360), .A2(n814), .ZN(n2682) );
  NOR2_X1 U22 ( .A1(n455), .A2(n451), .ZN(n327) );
  NOR2_X1 U23 ( .A1(n320), .A2(n319), .ZN(n576) );
  CLKBUF_X1 U24 ( .A(n811), .Z(n788) );
  CLKBUF_X1 U28 ( .A(regfile_data_ra_id[7]), .Z(n31) );
  INV_X1 U33 ( .A(n2299), .ZN(n107) );
  AND2_X1 U37 ( .A1(n1764), .A2(n1882), .ZN(n2209) );
  OR2_X1 U38 ( .A1(n2387), .A2(n814), .ZN(n2684) );
  NOR3_X1 U44 ( .A1(hwloop_we_int[2]), .A2(hwloop_we_int[0]), .A3(
        hwloop_we_int[1]), .ZN(n2574) );
  INV_X1 U45 ( .A(n638), .ZN(n778) );
  AND2_X1 U46 ( .A1(n2462), .A2(n2668), .ZN(n2647) );
  AND2_X1 U47 ( .A1(n2462), .A2(n2678), .ZN(n2648) );
  AND2_X1 U50 ( .A1(n2462), .A2(n2683), .ZN(n2649) );
  NOR2_X1 U51 ( .A1(n2427), .A2(n2426), .ZN(n2650) );
  AND2_X1 U52 ( .A1(n2462), .A2(instr_rdata_i[29]), .ZN(n2651) );
  NOR2_X1 U54 ( .A1(n2427), .A2(n1035), .ZN(n2652) );
  OR2_X1 U57 ( .A1(n2063), .A2(n2125), .ZN(n2655) );
  OAI21_X1 U58 ( .B1(n1046), .B2(n1101), .A(n1045), .ZN(n2656) );
  OAI21_X1 U59 ( .B1(n1046), .B2(n1101), .A(n1045), .ZN(n2469) );
  INV_X1 U61 ( .A(n2631), .ZN(n2657) );
  NAND2_X1 U65 ( .A1(n724), .A2(n723), .ZN(n2658) );
  XOR2_X1 U66 ( .A(n210), .B(pc_id_i[31]), .Z(n2659) );
  NAND2_X1 U67 ( .A1(n657), .A2(n656), .ZN(n2660) );
  NAND4_X1 U68 ( .A1(n1712), .A2(n1711), .A3(n1710), .A4(n1709), .ZN(n2661) );
  NAND4_X1 U69 ( .A1(n1712), .A2(n1711), .A3(n1710), .A4(n1709), .ZN(n2662) );
  NAND4_X1 U70 ( .A1(n1712), .A2(n1711), .A3(n1710), .A4(n1709), .ZN(n1971) );
  BUF_X1 U71 ( .A(regfile_alu_wdata_fw_i[15]), .Z(n2663) );
  AND3_X1 U75 ( .A1(n2076), .A2(n2075), .A3(n2655), .ZN(n2077) );
  NAND2_X1 U76 ( .A1(n2506), .A2(n1848), .ZN(n2664) );
  AND4_X1 U78 ( .A1(n1632), .A2(n1396), .A3(n1328), .A4(n1243), .ZN(n2665) );
  OAI21_X1 U81 ( .B1(n2665), .B2(n1983), .A(n1911), .ZN(n2666) );
  AND3_X1 U82 ( .A1(n2686), .A2(n2032), .A3(n2031), .ZN(n2034) );
  CLKBUF_X1 U84 ( .A(instr_rdata_i[28]), .Z(n2668) );
  NOR2_X1 U85 ( .A1(n2650), .A2(n2456), .ZN(n2435) );
  INV_X1 U87 ( .A(n2435), .ZN(n3517) );
  INV_X1 U88 ( .A(n311), .ZN(n2669) );
  OR2_X1 U89 ( .A1(n105), .A2(n104), .ZN(n2670) );
  INV_X1 U90 ( .A(n349), .ZN(n2672) );
  AND2_X1 U91 ( .A1(n272), .A2(n318), .ZN(n292) );
  NAND2_X1 U92 ( .A1(jump_target_mux_sel[1]), .A2(jump_target_mux_sel[0]), 
        .ZN(n272) );
  CLKBUF_X3 U98 ( .A(id_ready_o_BAR), .Z(n2577) );
  CLKBUF_X1 U114 ( .A(instr_rdata_i[19]), .Z(n116) );
  NOR2_X1 U115 ( .A1(n239), .A2(n238), .ZN(n490) );
  INV_X1 U116 ( .A(n2452), .ZN(n3486) );
  NAND3_X1 U142 ( .A1(n2681), .A2(n2682), .A3(n625), .ZN(hwloop_cnt[25]) );
  NAND2_X1 U144 ( .A1(regfile_alu_wdata_fw_i[25]), .A2(n788), .ZN(n2681) );
  NAND2_X1 U159 ( .A1(n473), .A2(n288), .ZN(n289) );
  OAI21_X1 U160 ( .B1(n108), .B2(n534), .A(n287), .ZN(n473) );
  BUF_X1 U161 ( .A(instr_rdata_i[26]), .Z(n2683) );
  INV_X1 U171 ( .A(n2569), .ZN(n3499) );
  NAND3_X1 U193 ( .A1(n2685), .A2(n646), .A3(n2684), .ZN(hwloop_cnt[28]) );
  NAND2_X1 U194 ( .A1(regfile_alu_wdata_fw_i[28]), .A2(n788), .ZN(n2685) );
  NAND2_X1 U195 ( .A1(n2014), .A2(n2033), .ZN(n2686) );
  NOR2_X1 U196 ( .A1(bmask_b_mux[1]), .A2(n1904), .ZN(n2688) );
  MUX2_X1 U197 ( .A(n2651), .B(n2688), .S(n3470), .Z(n3473) );
  NOR2_X1 U203 ( .A1(bmask_b_mux[1]), .A2(n1991), .ZN(n2689) );
  MUX2_X1 U204 ( .A(n2647), .B(n2689), .S(n3470), .Z(n3472) );
  NOR2_X1 U205 ( .A1(bmask_b_mux[1]), .A2(n1984), .ZN(n2690) );
  MUX2_X1 U221 ( .A(n2648), .B(n2690), .S(n3470), .Z(n3471) );
  NOR2_X1 U227 ( .A1(bmask_b_mux[1]), .A2(n1738), .ZN(n2691) );
  MUX2_X1 U228 ( .A(n2649), .B(n2691), .S(n3470), .Z(n3469) );
  OR2_X1 U240 ( .A1(n2652), .A2(n2650), .ZN(n2692) );
  AND2_X1 U261 ( .A1(n1032), .A2(regfile_we_id), .ZN(n2693) );
  INV_X1 U262 ( .A(n2570), .ZN(n3483) );
  AND2_X1 U263 ( .A1(n2533), .A2(n2532), .ZN(n2694) );
  INV_X1 U272 ( .A(n1822), .ZN(n3509) );
  INV_X1 U273 ( .A(n2521), .ZN(n3512) );
  INV_X1 U274 ( .A(n2508), .ZN(n3537) );
  INV_X1 U277 ( .A(n2515), .ZN(n3510) );
  AND2_X1 U2990 ( .A1(n778), .A2(alu_operator[2]), .ZN(n3489) );
  AND2_X1 U2991 ( .A1(n778), .A2(alu_operator[3]), .ZN(n3490) );
  AND2_X1 U2992 ( .A1(n778), .A2(alu_operator[4]), .ZN(n3491) );
  AND2_X1 U2993 ( .A1(n778), .A2(alu_operator[5]), .ZN(n3492) );
  AND2_X1 U2994 ( .A1(n778), .A2(alu_operator[6]), .ZN(n3493) );
  INV_X1 U2995 ( .A(n3460), .ZN(n3494) );
  AOI211_X1 U2996 ( .C1(n185), .C2(n1032), .A(alu_operator[0]), .B(n187), .ZN(
        n3460) );
  NOR2_X1 U2997 ( .A1(alu_operator[1]), .A2(n3461), .ZN(n3495) );
  INV_X1 U2998 ( .A(n2448), .ZN(n3461) );
  NAND2_X1 U2999 ( .A1(n605), .A2(n3462), .ZN(n3498) );
  INV_X1 U3000 ( .A(n187), .ZN(n3462) );
  AND2_X1 U3001 ( .A1(id_valid_o), .A2(csr_op[0]), .ZN(n3500) );
  AND2_X1 U3002 ( .A1(id_valid_o), .A2(csr_op[1]), .ZN(n3501) );
  NAND2_X1 U3003 ( .A1(id_valid_o), .A2(n605), .ZN(n3502) );
  NOR2_X1 U3004 ( .A1(n1034), .A2(n2570), .ZN(n3503) );
  NAND2_X1 U3005 ( .A1(n810), .A2(n605), .ZN(n3506) );
  NAND2_X1 U3006 ( .A1(n1923), .A2(n3463), .ZN(n3511) );
  AOI21_X1 U3007 ( .B1(scalar_replication), .B2(n1912), .A(n173), .ZN(n3463)
         );
  OAI21_X1 U3008 ( .B1(n3464), .B2(n3465), .A(n3466), .ZN(n3520) );
  NAND2_X1 U3009 ( .A1(n3465), .A2(n1205), .ZN(n3466) );
  INV_X1 U3010 ( .A(alu_bmask_b_mux_sel), .ZN(n3465) );
  AOI22_X1 U3011 ( .A1(n2462), .A2(n3467), .B1(bmask_b_mux[0]), .B2(n3468), 
        .ZN(n3464) );
  NAND2_X1 U3012 ( .A1(n2462), .A2(n2463), .ZN(n3468) );
  NOR2_X1 U3013 ( .A1(bmask_b_mux[0]), .A2(n2467), .ZN(n3467) );
  MUX2_X1 U3014 ( .A(n1229), .B(n3469), .S(alu_bmask_b_mux_sel), .Z(n3521) );
  INV_X1 U3015 ( .A(bmask_b_mux[0]), .ZN(n3470) );
  MUX2_X1 U3016 ( .A(n713), .B(n3471), .S(alu_bmask_b_mux_sel), .Z(n3522) );
  MUX2_X1 U3017 ( .A(n643), .B(n3472), .S(alu_bmask_b_mux_sel), .Z(n3523) );
  MUX2_X1 U3018 ( .A(n701), .B(n3473), .S(alu_bmask_b_mux_sel), .Z(n3524) );
  OAI21_X1 U3019 ( .B1(n659), .B2(alu_bmask_a_mux_sel), .A(n3474), .ZN(n3525)
         );
  NAND3_X1 U3020 ( .A1(alu_bmask_a_mux_sel), .A2(instr_rdata_i[25]), .A3(
        bmask_a_mux_0_), .ZN(n3474) );
  OAI21_X1 U3021 ( .B1(n2173), .B2(alu_bmask_a_mux_sel), .A(n3475), .ZN(n3526)
         );
  NAND3_X1 U3022 ( .A1(alu_bmask_a_mux_sel), .A2(n2683), .A3(bmask_a_mux_0_), 
        .ZN(n3475) );
  OAI21_X1 U3023 ( .B1(n2188), .B2(alu_bmask_a_mux_sel), .A(n3476), .ZN(n3527)
         );
  NAND3_X1 U3024 ( .A1(alu_bmask_a_mux_sel), .A2(n2678), .A3(bmask_a_mux_0_), 
        .ZN(n3476) );
  OAI21_X1 U3025 ( .B1(n2198), .B2(alu_bmask_a_mux_sel), .A(n3477), .ZN(n3528)
         );
  NAND3_X1 U3026 ( .A1(alu_bmask_a_mux_sel), .A2(n2668), .A3(bmask_a_mux_0_), 
        .ZN(n3477) );
  OAI21_X1 U3027 ( .B1(n2204), .B2(alu_bmask_a_mux_sel), .A(n3478), .ZN(n3529)
         );
  NAND3_X1 U3028 ( .A1(alu_bmask_a_mux_sel), .A2(instr_rdata_i[29]), .A3(
        bmask_a_mux_0_), .ZN(n3478) );
  NOR2_X1 U3029 ( .A1(n2463), .A2(mult_imm_mux_0_), .ZN(n3532) );
  NOR2_X1 U3030 ( .A1(n2428), .A2(mult_imm_mux_0_), .ZN(n3533) );
  NOR2_X1 U3031 ( .A1(n2429), .A2(mult_imm_mux_0_), .ZN(n3534) );
  NOR2_X1 U3032 ( .A1(n2430), .A2(mult_imm_mux_0_), .ZN(n3535) );
  NOR2_X1 U3033 ( .A1(n2431), .A2(mult_imm_mux_0_), .ZN(n3536) );
endmodule


module riscv_if_stage_2_128_0_1a110800 ( clk, rst_n, m_trap_base_addr_i, 
        u_trap_base_addr_i, trap_addr_mux_i, boot_addr_i, req_i, instr_req_o, 
        instr_addr_o, instr_gnt_i, instr_rvalid_i, instr_rdata_i, 
        instr_err_pmp_i, hwlp_dec_cnt_id_o, is_hwlp_id_o, instr_valid_id_o, 
        instr_rdata_id_o, is_compressed_id_o, illegal_c_insn_id_o, pc_if_o, 
        pc_id_o, is_fetch_failed_o, clear_instr_valid_i, pc_set_i, mepc_i, 
        uepc_i, depc_i, pc_mux_i, exc_pc_mux_i, exc_vec_pc_mux_i, 
        jump_target_id_i, jump_target_ex_i, hwlp_start_i, hwlp_end_i, 
        hwlp_cnt_i, halt_if_i, if_busy_o, perf_imiss_o, id_ready_i_BAR );
  input [23:0] m_trap_base_addr_i;
  input [23:0] u_trap_base_addr_i;
  input [30:0] boot_addr_i;
  output [31:0] instr_addr_o;
  input [127:0] instr_rdata_i;
  output [1:0] hwlp_dec_cnt_id_o;
  output [31:0] instr_rdata_id_o;
  output [31:0] pc_if_o;
  output [31:0] pc_id_o;
  input [31:0] mepc_i;
  input [31:0] uepc_i;
  input [31:0] depc_i;
  input [2:0] pc_mux_i;
  input [2:0] exc_pc_mux_i;
  input [4:0] exc_vec_pc_mux_i;
  input [31:0] jump_target_id_i;
  input [31:0] jump_target_ex_i;
  input [63:0] hwlp_start_i;
  input [63:0] hwlp_end_i;
  input [63:0] hwlp_cnt_i;
  input clk, rst_n, trap_addr_mux_i, req_i, instr_gnt_i, instr_rvalid_i,
         instr_err_pmp_i, clear_instr_valid_i, pc_set_i, halt_if_i,
         id_ready_i_BAR;
  output instr_req_o, is_hwlp_id_o, instr_valid_id_o, is_compressed_id_o,
         illegal_c_insn_id_o, is_fetch_failed_o, if_busy_o, perf_imiss_o;
  wire   branch_req, hwlp_jump, fetch_ready, fetch_valid, fetch_is_hwlp,
         offset_fsm_cs_0_, offset_fsm_ns_0_, n_2_net__1_, n_2_net__0_,
         instr_compressed_int, illegal_c_insn, is_hwlp_id_q, n243, n245, n246,
         n247, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n6,
         n7, n9, n10, n13, n14, n15, n16, n20, n21, n22, n23, n24, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n87, n88, n89, n90, n91, n93, n94, n95, n96, n97, n98, n99, n100,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n314, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n555, n561, n567, n572, n573, n574, n575,
         n584, n585, n586, n587, n589, n590, n591, n592, n593, n594, n595,
         n599, n600, n611, n620, n621, n625, n626, n627, n773, n774;
  wire   [31:0] hwlp_target;
  wire   [31:0] fetch_rdata;
  wire   [31:1] instr_decompressed;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4;

  AOI22_X1 U4 ( .A1(n479), .A2(m_trap_base_addr_i[7]), .B1(n507), .B2(
        boot_addr_i[14]), .ZN(n236) );
  NOR2_X1 U6 ( .A1(n69), .A2(pc_mux_i[1]), .ZN(n174) );
  AND2_X1 U8 ( .A1(pc_mux_i[1]), .A2(n40), .ZN(n223) );
  OR2_X1 U9 ( .A1(n38), .A2(n37), .ZN(n82) );
  CLKBUF_X1 U11 ( .A(id_ready_i_BAR), .Z(n38) );
  CLKBUF_X1 U12 ( .A(n501), .Z(n371) );
  AND2_X1 U13 ( .A1(pc_mux_i[1]), .A2(n14), .ZN(n132) );
  AND3_X1 U15 ( .A1(n372), .A2(n374), .A3(n373), .ZN(n13) );
  INV_X1 U16 ( .A(n60), .ZN(n14) );
  NAND2_X1 U17 ( .A1(pc_mux_i[0]), .A2(n423), .ZN(n60) );
  AOI22_X1 U19 ( .A1(n479), .A2(m_trap_base_addr_i[11]), .B1(boot_addr_i[18]), 
        .B2(n480), .ZN(n372) );
  BUF_X2 U20 ( .A(n132), .Z(n491) );
  AND2_X1 U21 ( .A1(req_i), .A2(offset_fsm_cs_0_), .ZN(n73) );
  AND4_X1 U22 ( .A1(n29), .A2(n58), .A3(n66), .A4(n28), .ZN(n27) );
  NOR2_X1 U23 ( .A1(pc_mux_i[0]), .A2(n67), .ZN(n96) );
  CLKBUF_X1 U24 ( .A(n510), .Z(n93) );
  AND2_X1 U25 ( .A1(n423), .A2(n376), .ZN(n15) );
  AND2_X1 U26 ( .A1(n379), .A2(n378), .ZN(n16) );
  NAND3_X1 U27 ( .A1(n426), .A2(n377), .A3(n15), .ZN(n379) );
  NOR3_X1 U28 ( .A1(n20), .A2(n21), .A3(n22), .ZN(n71) );
  AND2_X1 U29 ( .A1(n433), .A2(uepc_i[17]), .ZN(n20) );
  AND2_X1 U30 ( .A1(n471), .A2(jump_target_ex_i[17]), .ZN(n21) );
  AND2_X1 U31 ( .A1(n497), .A2(u_trap_base_addr_i[9]), .ZN(n22) );
  NOR2_X1 U32 ( .A1(n41), .A2(pc_mux_i[1]), .ZN(n204) );
  AND2_X1 U33 ( .A1(n237), .A2(n238), .ZN(n24) );
  NAND3_X1 U34 ( .A1(n57), .A2(n55), .A3(n56), .ZN(n335) );
  AOI21_X1 U35 ( .B1(m_trap_base_addr_i[12]), .B2(n479), .A(n23), .ZN(n384) );
  NAND2_X1 U36 ( .A1(n380), .A2(n16), .ZN(n23) );
  NAND3_X1 U37 ( .A1(n239), .A2(n236), .A3(n24), .ZN(n332) );
  NAND2_X1 U38 ( .A1(jump_target_id_i[30]), .A2(n410), .ZN(n487) );
  AOI21_X1 U39 ( .B1(jump_target_id_i[25]), .B2(n508), .A(n26), .ZN(n440) );
  AND2_X1 U40 ( .A1(n466), .A2(n437), .ZN(n26) );
  NAND3_X1 U41 ( .A1(n27), .A2(n71), .A3(n72), .ZN(n330) );
  NAND2_X1 U42 ( .A1(n463), .A2(mepc_i[17]), .ZN(n28) );
  NAND2_X1 U43 ( .A1(jump_target_id_i[17]), .A2(n476), .ZN(n29) );
  NAND2_X1 U44 ( .A1(n96), .A2(trap_addr_mux_i), .ZN(n70) );
  NAND2_X1 U45 ( .A1(n96), .A2(n68), .ZN(n69) );
  NOR2_X1 U46 ( .A1(n70), .A2(pc_mux_i[1]), .ZN(n167) );
  INV_X1 U47 ( .A(exc_pc_mux_i[0]), .ZN(n94) );
  AOI21_X1 U49 ( .B1(n368), .B2(u_trap_base_addr_i[11]), .A(n367), .ZN(n375)
         );
  AND2_X1 U50 ( .A1(n96), .A2(n95), .ZN(n154) );
  OR2_X2 U51 ( .A1(pc_set_i), .A2(n73), .ZN(branch_req) );
  INV_X1 U52 ( .A(n7), .ZN(n74) );
  INV_X1 U53 ( .A(halt_if_i), .ZN(n36) );
  NAND4_X1 U54 ( .A1(fetch_valid), .A2(n74), .A3(n36), .A4(n561), .ZN(n37) );
  NAND2_X1 U59 ( .A1(pc_mux_i[0]), .A2(pc_mux_i[2]), .ZN(n59) );
  INV_X1 U60 ( .A(n59), .ZN(n40) );
  BUF_X2 U61 ( .A(n223), .Z(n199) );
  NOR2_X1 U62 ( .A1(pc_mux_i[0]), .A2(pc_mux_i[2]), .ZN(n43) );
  INV_X1 U63 ( .A(n43), .ZN(n41) );
  BUF_X2 U64 ( .A(n204), .Z(n480) );
  AOI22_X1 U65 ( .A1(n432), .A2(depc_i[12]), .B1(n480), .B2(boot_addr_i[11]), 
        .ZN(n57) );
  INV_X1 U66 ( .A(pc_mux_i[2]), .ZN(n423) );
  NOR2_X1 U67 ( .A1(pc_mux_i[0]), .A2(n423), .ZN(n42) );
  AND2_X1 U68 ( .A1(pc_mux_i[1]), .A2(n42), .ZN(n139) );
  BUF_X2 U69 ( .A(n139), .Z(n433) );
  AOI22_X1 U70 ( .A1(n433), .A2(uepc_i[12]), .B1(n491), .B2(
        jump_target_ex_i[12]), .ZN(n56) );
  AND2_X1 U71 ( .A1(pc_mux_i[1]), .A2(n43), .ZN(n140) );
  BUF_X2 U72 ( .A(n140), .Z(n508) );
  INV_X1 U73 ( .A(pc_mux_i[1]), .ZN(n426) );
  INV_X1 U74 ( .A(exc_pc_mux_i[1]), .ZN(n44) );
  NAND2_X1 U75 ( .A1(pc_mux_i[2]), .A2(n44), .ZN(n67) );
  INV_X1 U76 ( .A(trap_addr_mux_i), .ZN(n68) );
  AOI22_X1 U77 ( .A1(n68), .A2(m_trap_base_addr_i[4]), .B1(
        u_trap_base_addr_i[4]), .B2(trap_addr_mux_i), .ZN(n45) );
  OR2_X1 U78 ( .A1(n67), .A2(n45), .ZN(n53) );
  NAND2_X1 U79 ( .A1(pc_id_o[6]), .A2(pc_id_o[7]), .ZN(n171) );
  NAND2_X1 U80 ( .A1(pc_id_o[8]), .A2(pc_id_o[9]), .ZN(n46) );
  NOR2_X1 U81 ( .A1(n171), .A2(n46), .ZN(n48) );
  NAND2_X1 U82 ( .A1(pc_id_o[4]), .A2(pc_id_o[5]), .ZN(n47) );
  NAND2_X1 U83 ( .A1(pc_id_o[3]), .A2(pc_id_o[2]), .ZN(n141) );
  NOR2_X1 U84 ( .A1(n47), .A2(n141), .ZN(n155) );
  NAND2_X1 U85 ( .A1(n48), .A2(n155), .ZN(n358) );
  INV_X1 U86 ( .A(n358), .ZN(n202) );
  NAND2_X1 U87 ( .A1(pc_id_o[10]), .A2(pc_id_o[11]), .ZN(n62) );
  INV_X1 U88 ( .A(n62), .ZN(n49) );
  NAND2_X1 U89 ( .A1(n202), .A2(n49), .ZN(n213) );
  XOR2_X1 U90 ( .A(n213), .B(n592), .Z(n50) );
  NAND3_X1 U91 ( .A1(n377), .A2(n50), .A3(n423), .ZN(n52) );
  NAND3_X1 U92 ( .A1(n377), .A2(pc_mux_i[2]), .A3(mepc_i[12]), .ZN(n51) );
  OAI211_X1 U93 ( .C1(n377), .C2(n53), .A(n52), .B(n51), .ZN(n54) );
  AOI22_X1 U94 ( .A1(n508), .A2(jump_target_id_i[12]), .B1(n426), .B2(n54), 
        .ZN(n55) );
  BUF_X2 U95 ( .A(n223), .Z(n432) );
  NAND2_X1 U96 ( .A1(n432), .A2(depc_i[17]), .ZN(n58) );
  BUF_X2 U97 ( .A(n140), .Z(n410) );
  NOR2_X1 U98 ( .A1(pc_mux_i[1]), .A2(n59), .ZN(n133) );
  NOR2_X1 U100 ( .A1(pc_mux_i[1]), .A2(n60), .ZN(n87) );
  NAND2_X1 U102 ( .A1(pc_id_o[12]), .A2(pc_id_o[13]), .ZN(n61) );
  NOR2_X1 U103 ( .A1(n62), .A2(n61), .ZN(n357) );
  NAND2_X1 U104 ( .A1(n202), .A2(n357), .ZN(n233) );
  INV_X1 U105 ( .A(n233), .ZN(n224) );
  NAND2_X1 U106 ( .A1(pc_id_o[14]), .A2(pc_id_o[15]), .ZN(n355) );
  INV_X1 U107 ( .A(n355), .ZN(n63) );
  NAND2_X1 U108 ( .A1(n224), .A2(n63), .ZN(n240) );
  NOR2_X1 U109 ( .A1(n240), .A2(n590), .ZN(n64) );
  XNOR2_X1 U110 ( .A(n64), .B(n586), .ZN(n65) );
  NAND2_X1 U111 ( .A1(n627), .A2(n65), .ZN(n66) );
  AOI22_X1 U114 ( .A1(n507), .A2(boot_addr_i[16]), .B1(n509), .B2(
        m_trap_base_addr_i[9]), .ZN(n72) );
  BUF_X2 U115 ( .A(n167), .Z(n497) );
  NAND3_X1 U116 ( .A1(n74), .A2(req_i), .A3(n561), .ZN(n75) );
  NOR2_X1 U117 ( .A1(halt_if_i), .A2(n75), .ZN(n76) );
  NAND2_X1 U118 ( .A1(fetch_valid), .A2(n76), .ZN(n77) );
  NOR2_X1 U119 ( .A1(id_ready_i_BAR), .A2(n77), .ZN(fetch_ready) );
  AND2_X1 U120 ( .A1(instr_valid_id_o), .A2(is_hwlp_id_q), .ZN(is_hwlp_id_o)
         );
  AND2_X1 U121 ( .A1(is_hwlp_id_o), .A2(hwlp_dec_cnt_id_o[0]), .ZN(n_2_net__0_) );
  AND2_X1 U122 ( .A1(is_hwlp_id_o), .A2(hwlp_dec_cnt_id_o[1]), .ZN(n_2_net__1_) );
  INV_X1 U123 ( .A(req_i), .ZN(n78) );
  NAND2_X1 U124 ( .A1(n78), .A2(offset_fsm_cs_0_), .ZN(n79) );
  NOR2_X1 U125 ( .A1(n7), .A2(n79), .ZN(offset_fsm_ns_0_) );
  NAND2_X1 U126 ( .A1(hwlp_jump), .A2(n10), .ZN(n80) );
  OAI21_X1 U127 ( .B1(hwlp_jump), .B2(n599), .A(n80), .ZN(n246) );
  NAND2_X1 U128 ( .A1(n555), .A2(fetch_is_hwlp), .ZN(n85) );
  NAND2_X1 U129 ( .A1(n85), .A2(hwlp_dec_cnt_id_o[0]), .ZN(n81) );
  OAI21_X1 U130 ( .B1(n85), .B2(n599), .A(n81), .ZN(n315) );
  OAI21_X1 U131 ( .B1(clear_instr_valid_i), .B2(n611), .A(n82), .ZN(n247) );
  INV_X1 U132 ( .A(n82), .ZN(n555) );
  NAND2_X1 U134 ( .A1(n9), .A2(hwlp_jump), .ZN(n83) );
  OAI21_X1 U135 ( .B1(hwlp_jump), .B2(n600), .A(n83), .ZN(n245) );
  NAND2_X1 U136 ( .A1(n85), .A2(hwlp_dec_cnt_id_o[1]), .ZN(n84) );
  OAI21_X1 U137 ( .B1(n85), .B2(n600), .A(n84), .ZN(n243) );
  AOI22_X1 U140 ( .A1(n508), .A2(jump_target_id_i[1]), .B1(n491), .B2(
        jump_target_ex_i[1]), .ZN(n91) );
  BUF_X2 U141 ( .A(n139), .Z(n496) );
  BUF_X2 U142 ( .A(n87), .Z(n501) );
  AOI22_X1 U143 ( .A1(n496), .A2(uepc_i[1]), .B1(n371), .B2(pc_id_o[1]), .ZN(
        n90) );
  AOI22_X1 U144 ( .A1(n506), .A2(depc_i[1]), .B1(n6), .B2(boot_addr_i[0]), 
        .ZN(n89) );
  NAND2_X1 U145 ( .A1(n93), .A2(mepc_i[1]), .ZN(n88) );
  NAND4_X1 U146 ( .A1(n91), .A2(n90), .A3(n89), .A4(n88), .ZN(n346) );
  BUF_X2 U150 ( .A(n132), .Z(n471) );
  AOI22_X1 U151 ( .A1(n496), .A2(uepc_i[2]), .B1(n505), .B2(
        jump_target_ex_i[2]), .ZN(n100) );
  AOI22_X1 U152 ( .A1(n199), .A2(depc_i[2]), .B1(n476), .B2(
        jump_target_id_i[2]), .ZN(n99) );
  AOI22_X1 U153 ( .A1(mepc_i[2]), .A2(n93), .B1(n371), .B2(n567), .ZN(n98) );
  NOR2_X1 U154 ( .A1(pc_mux_i[1]), .A2(n94), .ZN(n95) );
  AOI22_X1 U155 ( .A1(n6), .A2(boot_addr_i[1]), .B1(n154), .B2(
        exc_vec_pc_mux_i[0]), .ZN(n97) );
  NAND4_X1 U156 ( .A1(n100), .A2(n99), .A3(n98), .A4(n97), .ZN(n345) );
  BUF_X2 U220 ( .A(n132), .Z(n505) );
  AOI22_X1 U221 ( .A1(n496), .A2(uepc_i[3]), .B1(n505), .B2(
        jump_target_ex_i[3]), .ZN(n138) );
  AOI22_X1 U222 ( .A1(n506), .A2(depc_i[3]), .B1(n410), .B2(
        jump_target_id_i[3]), .ZN(n137) );
  XNOR2_X1 U224 ( .A(n30), .B(pc_id_o[2]), .ZN(n134) );
  AOI22_X1 U225 ( .A1(n93), .A2(mepc_i[3]), .B1(n371), .B2(n134), .ZN(n136) );
  AOI22_X1 U226 ( .A1(n6), .A2(boot_addr_i[2]), .B1(n154), .B2(
        exc_vec_pc_mux_i[1]), .ZN(n135) );
  NAND4_X1 U227 ( .A1(n138), .A2(n137), .A3(n136), .A4(n135), .ZN(n344) );
  BUF_X2 U228 ( .A(n139), .Z(n451) );
  AOI22_X1 U229 ( .A1(n451), .A2(uepc_i[4]), .B1(n505), .B2(
        jump_target_ex_i[4]), .ZN(n146) );
  BUF_X2 U230 ( .A(n140), .Z(n476) );
  AOI22_X1 U231 ( .A1(n199), .A2(depc_i[4]), .B1(n508), .B2(
        jump_target_id_i[4]), .ZN(n145) );
  INV_X1 U232 ( .A(n141), .ZN(n147) );
  XNOR2_X1 U233 ( .A(n572), .B(n147), .ZN(n142) );
  AOI22_X1 U234 ( .A1(n626), .A2(mepc_i[4]), .B1(n501), .B2(n142), .ZN(n144)
         );
  AOI22_X1 U235 ( .A1(n480), .A2(boot_addr_i[3]), .B1(n154), .B2(
        exc_vec_pc_mux_i[2]), .ZN(n143) );
  NAND4_X1 U236 ( .A1(n144), .A2(n145), .A3(n146), .A4(n143), .ZN(n343) );
  AOI22_X1 U237 ( .A1(n433), .A2(uepc_i[5]), .B1(n505), .B2(
        jump_target_ex_i[5]), .ZN(n153) );
  AOI22_X1 U238 ( .A1(n199), .A2(depc_i[5]), .B1(n476), .B2(
        jump_target_id_i[5]), .ZN(n152) );
  NAND2_X1 U239 ( .A1(n147), .A2(pc_id_o[4]), .ZN(n148) );
  XOR2_X1 U240 ( .A(n148), .B(n587), .Z(n149) );
  AOI22_X1 U241 ( .A1(n463), .A2(mepc_i[5]), .B1(n627), .B2(n149), .ZN(n151)
         );
  AOI22_X1 U242 ( .A1(n507), .A2(boot_addr_i[4]), .B1(n154), .B2(
        exc_vec_pc_mux_i[3]), .ZN(n150) );
  NAND4_X1 U243 ( .A1(n150), .A2(n152), .A3(n151), .A4(n153), .ZN(n342) );
  AOI22_X1 U244 ( .A1(n433), .A2(uepc_i[6]), .B1(n505), .B2(
        jump_target_ex_i[6]), .ZN(n160) );
  AOI22_X1 U245 ( .A1(n199), .A2(depc_i[6]), .B1(n508), .B2(
        jump_target_id_i[6]), .ZN(n159) );
  AOI22_X1 U246 ( .A1(n480), .A2(boot_addr_i[5]), .B1(n154), .B2(
        exc_vec_pc_mux_i[4]), .ZN(n158) );
  INV_X1 U247 ( .A(n155), .ZN(n172) );
  XOR2_X1 U248 ( .A(n172), .B(n593), .Z(n156) );
  AOI22_X1 U249 ( .A1(n626), .A2(mepc_i[6]), .B1(n466), .B2(n156), .ZN(n157)
         );
  NAND4_X1 U250 ( .A1(n160), .A2(n159), .A3(n158), .A4(n157), .ZN(n341) );
  AOI22_X1 U251 ( .A1(n508), .A2(jump_target_id_i[7]), .B1(n433), .B2(
        uepc_i[7]), .ZN(n166) );
  NOR2_X1 U252 ( .A1(n172), .A2(n593), .ZN(n161) );
  XNOR2_X1 U253 ( .A(n161), .B(n589), .ZN(n162) );
  AOI22_X1 U254 ( .A1(n491), .A2(jump_target_ex_i[7]), .B1(n466), .B2(n162), 
        .ZN(n165) );
  AOI22_X1 U255 ( .A1(n432), .A2(depc_i[7]), .B1(n485), .B2(boot_addr_i[6]), 
        .ZN(n164) );
  NAND2_X1 U256 ( .A1(n510), .A2(mepc_i[7]), .ZN(n163) );
  NAND4_X1 U257 ( .A1(n166), .A2(n165), .A3(n164), .A4(n163), .ZN(n340) );
  NAND2_X1 U258 ( .A1(n505), .A2(jump_target_ex_i[8]), .ZN(n170) );
  NAND2_X1 U259 ( .A1(n451), .A2(uepc_i[8]), .ZN(n169) );
  NAND2_X1 U261 ( .A1(n497), .A2(u_trap_base_addr_i[0]), .ZN(n168) );
  AND3_X1 U262 ( .A1(n170), .A2(n169), .A3(n168), .ZN(n178) );
  AOI22_X1 U263 ( .A1(n506), .A2(depc_i[8]), .B1(n508), .B2(
        jump_target_id_i[8]), .ZN(n177) );
  NOR2_X1 U264 ( .A1(n172), .A2(n171), .ZN(n182) );
  XNOR2_X1 U265 ( .A(n182), .B(n575), .ZN(n173) );
  AOI22_X1 U266 ( .A1(n626), .A2(mepc_i[8]), .B1(n501), .B2(n173), .ZN(n176)
         );
  BUF_X2 U267 ( .A(n174), .Z(n479) );
  AOI22_X1 U268 ( .A1(n480), .A2(boot_addr_i[7]), .B1(n479), .B2(
        m_trap_base_addr_i[0]), .ZN(n175) );
  NAND4_X1 U269 ( .A1(n178), .A2(n177), .A3(n176), .A4(n175), .ZN(n339) );
  NAND2_X1 U270 ( .A1(n433), .A2(uepc_i[9]), .ZN(n181) );
  NAND2_X1 U271 ( .A1(n471), .A2(jump_target_ex_i[9]), .ZN(n180) );
  NAND2_X1 U272 ( .A1(n497), .A2(u_trap_base_addr_i[1]), .ZN(n179) );
  AND3_X1 U273 ( .A1(n180), .A2(n181), .A3(n179), .ZN(n188) );
  AOI22_X1 U274 ( .A1(n506), .A2(depc_i[9]), .B1(n410), .B2(
        jump_target_id_i[9]), .ZN(n187) );
  NAND2_X1 U275 ( .A1(n182), .A2(pc_id_o[8]), .ZN(n183) );
  XOR2_X1 U276 ( .A(n183), .B(n31), .Z(n184) );
  AOI22_X1 U277 ( .A1(n510), .A2(mepc_i[9]), .B1(n627), .B2(n184), .ZN(n186)
         );
  AOI22_X1 U278 ( .A1(n480), .A2(boot_addr_i[8]), .B1(n479), .B2(
        m_trap_base_addr_i[1]), .ZN(n185) );
  NAND4_X1 U279 ( .A1(n188), .A2(n187), .A3(n186), .A4(n185), .ZN(n338) );
  NAND2_X1 U280 ( .A1(n496), .A2(uepc_i[10]), .ZN(n191) );
  NAND2_X1 U281 ( .A1(n491), .A2(jump_target_ex_i[10]), .ZN(n190) );
  NAND2_X1 U282 ( .A1(n497), .A2(u_trap_base_addr_i[2]), .ZN(n189) );
  AND3_X1 U283 ( .A1(n191), .A2(n190), .A3(n189), .ZN(n196) );
  AOI22_X1 U284 ( .A1(n506), .A2(depc_i[10]), .B1(n476), .B2(
        jump_target_id_i[10]), .ZN(n195) );
  XNOR2_X1 U285 ( .A(n202), .B(n574), .ZN(n192) );
  AOI22_X1 U286 ( .A1(n463), .A2(mepc_i[10]), .B1(n501), .B2(n192), .ZN(n194)
         );
  AOI22_X1 U287 ( .A1(n507), .A2(boot_addr_i[9]), .B1(n509), .B2(
        m_trap_base_addr_i[2]), .ZN(n193) );
  NAND4_X1 U288 ( .A1(n196), .A2(n195), .A3(n194), .A4(n193), .ZN(n337) );
  INV_X1 U289 ( .A(n377), .ZN(n425) );
  NAND3_X1 U290 ( .A1(n94), .A2(exc_pc_mux_i[1]), .A3(pc_mux_i[2]), .ZN(n197)
         );
  NOR2_X1 U291 ( .A1(pc_mux_i[1]), .A2(n197), .ZN(n198) );
  AND2_X2 U292 ( .A1(n425), .A2(n198), .ZN(n460) );
  AOI21_X1 U293 ( .B1(n451), .B2(uepc_i[11]), .A(n460), .ZN(n201) );
  AOI22_X1 U294 ( .A1(n432), .A2(depc_i[11]), .B1(n471), .B2(
        jump_target_ex_i[11]), .ZN(n200) );
  AND2_X1 U295 ( .A1(n200), .A2(n201), .ZN(n209) );
  AOI22_X1 U296 ( .A1(n410), .A2(jump_target_id_i[11]), .B1(n510), .B2(
        mepc_i[11]), .ZN(n208) );
  NAND2_X1 U297 ( .A1(n202), .A2(pc_id_o[10]), .ZN(n203) );
  XOR2_X1 U298 ( .A(n203), .B(n32), .Z(n205) );
  BUF_X1 U299 ( .A(n204), .Z(n485) );
  AOI22_X1 U300 ( .A1(n627), .A2(n205), .B1(n480), .B2(boot_addr_i[10]), .ZN(
        n207) );
  AOI22_X1 U301 ( .A1(n509), .A2(m_trap_base_addr_i[3]), .B1(n472), .B2(
        u_trap_base_addr_i[3]), .ZN(n206) );
  NAND4_X1 U302 ( .A1(n209), .A2(n208), .A3(n207), .A4(n206), .ZN(n336) );
  NAND2_X1 U303 ( .A1(n496), .A2(uepc_i[13]), .ZN(n212) );
  NAND2_X1 U304 ( .A1(n491), .A2(jump_target_ex_i[13]), .ZN(n211) );
  NAND2_X1 U305 ( .A1(n497), .A2(u_trap_base_addr_i[5]), .ZN(n210) );
  AND3_X1 U306 ( .A1(n212), .A2(n211), .A3(n210), .ZN(n219) );
  AOI22_X1 U307 ( .A1(n199), .A2(depc_i[13]), .B1(n476), .B2(
        jump_target_id_i[13]), .ZN(n218) );
  NOR2_X1 U308 ( .A1(n213), .A2(n592), .ZN(n214) );
  XNOR2_X1 U309 ( .A(n214), .B(n33), .ZN(n215) );
  AOI22_X1 U310 ( .A1(n626), .A2(mepc_i[13]), .B1(n501), .B2(n215), .ZN(n217)
         );
  AOI22_X1 U311 ( .A1(n507), .A2(boot_addr_i[12]), .B1(n479), .B2(
        m_trap_base_addr_i[5]), .ZN(n216) );
  NAND4_X1 U312 ( .A1(n219), .A2(n218), .A3(n217), .A4(n216), .ZN(n334) );
  NAND2_X1 U313 ( .A1(n471), .A2(jump_target_ex_i[14]), .ZN(n222) );
  NAND2_X1 U314 ( .A1(n451), .A2(uepc_i[14]), .ZN(n221) );
  NAND2_X1 U315 ( .A1(n497), .A2(u_trap_base_addr_i[6]), .ZN(n220) );
  AND3_X1 U316 ( .A1(n220), .A2(n221), .A3(n222), .ZN(n229) );
  BUF_X1 U317 ( .A(n223), .Z(n506) );
  AOI22_X1 U318 ( .A1(n199), .A2(depc_i[14]), .B1(n410), .B2(
        jump_target_id_i[14]), .ZN(n228) );
  XNOR2_X1 U319 ( .A(n224), .B(n34), .ZN(n225) );
  AOI22_X1 U320 ( .A1(n510), .A2(mepc_i[14]), .B1(n627), .B2(n225), .ZN(n227)
         );
  AOI22_X1 U321 ( .A1(n507), .A2(boot_addr_i[13]), .B1(n479), .B2(
        m_trap_base_addr_i[6]), .ZN(n226) );
  NAND4_X1 U322 ( .A1(n229), .A2(n228), .A3(n227), .A4(n226), .ZN(n333) );
  NAND2_X1 U323 ( .A1(n471), .A2(jump_target_ex_i[15]), .ZN(n231) );
  NAND2_X1 U324 ( .A1(n433), .A2(uepc_i[15]), .ZN(n230) );
  NAND2_X1 U325 ( .A1(n231), .A2(n230), .ZN(n232) );
  AOI21_X1 U326 ( .B1(n368), .B2(u_trap_base_addr_i[7]), .A(n232), .ZN(n239)
         );
  AOI22_X1 U327 ( .A1(n199), .A2(depc_i[15]), .B1(n410), .B2(
        jump_target_id_i[15]), .ZN(n238) );
  NOR2_X1 U328 ( .A1(n233), .A2(n34), .ZN(n234) );
  XNOR2_X1 U329 ( .A(n234), .B(n35), .ZN(n235) );
  AOI22_X1 U330 ( .A1(n510), .A2(mepc_i[15]), .B1(n501), .B2(n235), .ZN(n237)
         );
  AOI22_X1 U331 ( .A1(n463), .A2(mepc_i[16]), .B1(n485), .B2(boot_addr_i[15]), 
        .ZN(n314) );
  XOR2_X1 U332 ( .A(n240), .B(n590), .Z(n241) );
  AOI22_X1 U333 ( .A1(n432), .A2(depc_i[16]), .B1(n466), .B2(n241), .ZN(n242)
         );
  AND2_X1 U334 ( .A1(n242), .A2(n314), .ZN(n350) );
  AOI22_X1 U335 ( .A1(n509), .A2(m_trap_base_addr_i[8]), .B1(n472), .B2(
        u_trap_base_addr_i[8]), .ZN(n349) );
  AOI21_X1 U336 ( .B1(n451), .B2(uepc_i[16]), .A(n460), .ZN(n348) );
  AOI22_X1 U337 ( .A1(n508), .A2(jump_target_id_i[16]), .B1(n491), .B2(
        jump_target_ex_i[16]), .ZN(n347) );
  NAND4_X1 U338 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(n331) );
  NAND2_X1 U339 ( .A1(n433), .A2(uepc_i[18]), .ZN(n353) );
  NAND2_X1 U340 ( .A1(n505), .A2(jump_target_ex_i[18]), .ZN(n352) );
  NAND2_X1 U341 ( .A1(n497), .A2(u_trap_base_addr_i[10]), .ZN(n351) );
  AND3_X1 U342 ( .A1(n351), .A2(n353), .A3(n352), .ZN(n364) );
  AOI22_X1 U343 ( .A1(n199), .A2(depc_i[18]), .B1(n410), .B2(
        jump_target_id_i[18]), .ZN(n363) );
  NAND2_X1 U344 ( .A1(pc_id_o[16]), .A2(pc_id_o[17]), .ZN(n354) );
  NOR2_X1 U345 ( .A1(n355), .A2(n354), .ZN(n356) );
  NAND2_X1 U346 ( .A1(n357), .A2(n356), .ZN(n359) );
  NOR2_X1 U347 ( .A1(n359), .A2(n358), .ZN(n420) );
  INV_X1 U348 ( .A(n420), .ZN(n412) );
  XOR2_X1 U349 ( .A(n412), .B(n591), .Z(n360) );
  AOI22_X1 U350 ( .A1(n626), .A2(mepc_i[18]), .B1(n627), .B2(n360), .ZN(n362)
         );
  AOI22_X1 U351 ( .A1(n480), .A2(boot_addr_i[17]), .B1(n479), .B2(
        m_trap_base_addr_i[10]), .ZN(n361) );
  NAND4_X1 U352 ( .A1(n364), .A2(n363), .A3(n362), .A4(n361), .ZN(n329) );
  NAND2_X1 U353 ( .A1(n471), .A2(jump_target_ex_i[19]), .ZN(n366) );
  AOI22_X1 U356 ( .A1(n199), .A2(depc_i[19]), .B1(jump_target_id_i[19]), .B2(
        n508), .ZN(n374) );
  NOR2_X1 U357 ( .A1(n412), .A2(n591), .ZN(n369) );
  XNOR2_X1 U358 ( .A(n369), .B(n585), .ZN(n370) );
  AOI22_X1 U359 ( .A1(n463), .A2(mepc_i[19]), .B1(n627), .B2(n370), .ZN(n373)
         );
  INV_X1 U360 ( .A(n460), .ZN(n380) );
  NAND2_X1 U361 ( .A1(pc_id_o[18]), .A2(pc_id_o[19]), .ZN(n399) );
  NOR2_X1 U362 ( .A1(n412), .A2(n399), .ZN(n388) );
  XNOR2_X1 U363 ( .A(n388), .B(n573), .ZN(n376) );
  NAND4_X1 U364 ( .A1(pc_mux_i[1]), .A2(pc_mux_i[2]), .A3(n377), .A4(
        depc_i[20]), .ZN(n378) );
  AOI22_X1 U365 ( .A1(n496), .A2(uepc_i[20]), .B1(n507), .B2(boot_addr_i[19]), 
        .ZN(n383) );
  AOI22_X1 U366 ( .A1(n476), .A2(jump_target_id_i[20]), .B1(n510), .B2(
        mepc_i[20]), .ZN(n382) );
  AOI22_X1 U367 ( .A1(n491), .A2(jump_target_ex_i[20]), .B1(n472), .B2(
        u_trap_base_addr_i[12]), .ZN(n381) );
  NAND4_X1 U368 ( .A1(n384), .A2(n383), .A3(n382), .A4(n381), .ZN(n327) );
  NAND2_X1 U369 ( .A1(n433), .A2(uepc_i[21]), .ZN(n387) );
  NAND2_X1 U370 ( .A1(n505), .A2(jump_target_ex_i[21]), .ZN(n386) );
  NAND2_X1 U371 ( .A1(n472), .A2(u_trap_base_addr_i[13]), .ZN(n385) );
  AND3_X1 U372 ( .A1(n387), .A2(n386), .A3(n385), .ZN(n394) );
  AOI22_X1 U373 ( .A1(n506), .A2(depc_i[21]), .B1(n410), .B2(
        jump_target_id_i[21]), .ZN(n393) );
  NAND2_X1 U374 ( .A1(n388), .A2(pc_id_o[20]), .ZN(n389) );
  XOR2_X1 U375 ( .A(n389), .B(n584), .Z(n390) );
  AOI22_X1 U376 ( .A1(n626), .A2(mepc_i[21]), .B1(n627), .B2(n390), .ZN(n392)
         );
  AOI22_X1 U377 ( .A1(n507), .A2(boot_addr_i[20]), .B1(n479), .B2(
        m_trap_base_addr_i[13]), .ZN(n391) );
  NAND4_X1 U378 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(n326) );
  NAND2_X1 U379 ( .A1(n451), .A2(uepc_i[22]), .ZN(n397) );
  NAND2_X1 U380 ( .A1(n491), .A2(jump_target_ex_i[22]), .ZN(n396) );
  NAND2_X1 U381 ( .A1(n472), .A2(u_trap_base_addr_i[14]), .ZN(n395) );
  AND3_X1 U382 ( .A1(n397), .A2(n396), .A3(n395), .ZN(n406) );
  AOI22_X1 U383 ( .A1(n506), .A2(depc_i[22]), .B1(n410), .B2(
        jump_target_id_i[22]), .ZN(n405) );
  NAND2_X1 U384 ( .A1(pc_id_o[20]), .A2(pc_id_o[21]), .ZN(n398) );
  NOR2_X1 U385 ( .A1(n399), .A2(n398), .ZN(n411) );
  INV_X1 U386 ( .A(n411), .ZN(n400) );
  NOR2_X1 U387 ( .A1(n412), .A2(n400), .ZN(n401) );
  XNOR2_X1 U388 ( .A(n401), .B(n594), .ZN(n402) );
  AOI22_X1 U389 ( .A1(n626), .A2(mepc_i[22]), .B1(n501), .B2(n402), .ZN(n404)
         );
  AOI22_X1 U390 ( .A1(n507), .A2(boot_addr_i[21]), .B1(n509), .B2(
        m_trap_base_addr_i[14]), .ZN(n403) );
  NAND4_X1 U391 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(n325) );
  NAND2_X1 U392 ( .A1(n491), .A2(jump_target_ex_i[23]), .ZN(n409) );
  NAND2_X1 U393 ( .A1(n451), .A2(uepc_i[23]), .ZN(n408) );
  NAND2_X1 U394 ( .A1(n472), .A2(u_trap_base_addr_i[15]), .ZN(n407) );
  AND3_X1 U395 ( .A1(n409), .A2(n408), .A3(n407), .ZN(n418) );
  AOI22_X1 U396 ( .A1(n199), .A2(depc_i[23]), .B1(n410), .B2(
        jump_target_id_i[23]), .ZN(n417) );
  NAND2_X1 U397 ( .A1(n411), .A2(pc_id_o[22]), .ZN(n419) );
  NOR2_X1 U398 ( .A1(n412), .A2(n419), .ZN(n413) );
  XNOR2_X1 U399 ( .A(n413), .B(n595), .ZN(n414) );
  AOI22_X1 U400 ( .A1(n626), .A2(mepc_i[23]), .B1(n627), .B2(n414), .ZN(n416)
         );
  AOI22_X1 U401 ( .A1(n507), .A2(boot_addr_i[22]), .B1(n509), .B2(
        m_trap_base_addr_i[15]), .ZN(n415) );
  NAND4_X1 U402 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(n324) );
  AOI22_X1 U403 ( .A1(n506), .A2(depc_i[24]), .B1(n491), .B2(
        jump_target_ex_i[24]), .ZN(n431) );
  AOI22_X1 U404 ( .A1(n476), .A2(jump_target_id_i[24]), .B1(n480), .B2(
        boot_addr_i[23]), .ZN(n430) );
  AOI22_X1 U405 ( .A1(n509), .A2(m_trap_base_addr_i[16]), .B1(n472), .B2(
        u_trap_base_addr_i[16]), .ZN(n429) );
  NOR2_X1 U406 ( .A1(n419), .A2(n595), .ZN(n421) );
  AND2_X1 U407 ( .A1(n421), .A2(n420), .ZN(n436) );
  AOI22_X1 U408 ( .A1(n423), .A2(n422), .B1(mepc_i[24]), .B2(pc_mux_i[2]), 
        .ZN(n424) );
  NOR2_X1 U409 ( .A1(n425), .A2(n424), .ZN(n427) );
  AOI22_X1 U410 ( .A1(n451), .A2(uepc_i[24]), .B1(n427), .B2(n426), .ZN(n428)
         );
  NAND4_X1 U411 ( .A1(n431), .A2(n430), .A3(n429), .A4(n428), .ZN(n323) );
  AOI22_X1 U412 ( .A1(n199), .A2(depc_i[25]), .B1(n471), .B2(
        jump_target_ex_i[25]), .ZN(n435) );
  AOI21_X1 U413 ( .B1(n433), .B2(uepc_i[25]), .A(n460), .ZN(n434) );
  AND2_X1 U414 ( .A1(n435), .A2(n434), .ZN(n441) );
  HA_X1 U415 ( .A(n436), .B(pc_id_o[24]), .CO(n445), .S(n422) );
  AOI22_X1 U416 ( .A1(n463), .A2(mepc_i[25]), .B1(n480), .B2(boot_addr_i[24]), 
        .ZN(n439) );
  AOI22_X1 U417 ( .A1(n509), .A2(m_trap_base_addr_i[17]), .B1(n472), .B2(
        u_trap_base_addr_i[17]), .ZN(n438) );
  NAND4_X1 U418 ( .A1(n441), .A2(n440), .A3(n439), .A4(n438), .ZN(n322) );
  NAND2_X1 U419 ( .A1(n505), .A2(jump_target_ex_i[26]), .ZN(n444) );
  NAND2_X1 U420 ( .A1(n451), .A2(uepc_i[26]), .ZN(n443) );
  NAND2_X1 U421 ( .A1(n472), .A2(u_trap_base_addr_i[18]), .ZN(n442) );
  AND3_X1 U422 ( .A1(n444), .A2(n443), .A3(n442), .ZN(n450) );
  AOI22_X1 U423 ( .A1(n506), .A2(depc_i[26]), .B1(n476), .B2(
        jump_target_id_i[26]), .ZN(n449) );
  HA_X1 U424 ( .A(n445), .B(pc_id_o[25]), .CO(n454), .S(n437) );
  AOI22_X1 U425 ( .A1(n510), .A2(mepc_i[26]), .B1(n501), .B2(n446), .ZN(n448)
         );
  AOI22_X1 U426 ( .A1(n507), .A2(boot_addr_i[25]), .B1(n479), .B2(
        m_trap_base_addr_i[18]), .ZN(n447) );
  NAND4_X1 U427 ( .A1(n450), .A2(n449), .A3(n448), .A4(n447), .ZN(n321) );
  AOI21_X1 U428 ( .B1(n451), .B2(uepc_i[27]), .A(n460), .ZN(n453) );
  AOI22_X1 U429 ( .A1(n432), .A2(depc_i[27]), .B1(n505), .B2(
        jump_target_ex_i[27]), .ZN(n452) );
  AND2_X1 U430 ( .A1(n452), .A2(n453), .ZN(n459) );
  HA_X1 U431 ( .A(n454), .B(pc_id_o[26]), .CO(n464), .S(n446) );
  AOI22_X1 U432 ( .A1(n476), .A2(jump_target_id_i[27]), .B1(n501), .B2(n455), 
        .ZN(n458) );
  AOI22_X1 U433 ( .A1(n510), .A2(mepc_i[27]), .B1(n507), .B2(boot_addr_i[26]), 
        .ZN(n457) );
  AOI22_X1 U434 ( .A1(n509), .A2(m_trap_base_addr_i[19]), .B1(n472), .B2(
        u_trap_base_addr_i[19]), .ZN(n456) );
  NAND4_X1 U435 ( .A1(n459), .A2(n458), .A3(n457), .A4(n456), .ZN(n320) );
  AOI21_X1 U437 ( .B1(n496), .B2(uepc_i[28]), .A(n460), .ZN(n461) );
  AOI22_X1 U439 ( .A1(n410), .A2(jump_target_id_i[28]), .B1(n626), .B2(
        mepc_i[28]), .ZN(n469) );
  HA_X1 U440 ( .A(n464), .B(pc_id_o[27]), .CO(n477), .S(n455) );
  AOI22_X1 U441 ( .A1(n627), .A2(n465), .B1(n507), .B2(boot_addr_i[27]), .ZN(
        n468) );
  AOI22_X1 U442 ( .A1(n509), .A2(m_trap_base_addr_i[20]), .B1(n472), .B2(
        u_trap_base_addr_i[20]), .ZN(n467) );
  NAND4_X1 U443 ( .A1(n470), .A2(n469), .A3(n468), .A4(n467), .ZN(n319) );
  NAND2_X1 U444 ( .A1(n491), .A2(jump_target_ex_i[29]), .ZN(n475) );
  NAND2_X1 U445 ( .A1(n496), .A2(uepc_i[29]), .ZN(n474) );
  NAND2_X1 U446 ( .A1(n497), .A2(u_trap_base_addr_i[21]), .ZN(n473) );
  AND3_X1 U447 ( .A1(n475), .A2(n474), .A3(n473), .ZN(n484) );
  AOI22_X1 U448 ( .A1(n506), .A2(depc_i[29]), .B1(n476), .B2(
        jump_target_id_i[29]), .ZN(n483) );
  HA_X1 U449 ( .A(n477), .B(pc_id_o[28]), .CO(n489), .S(n465) );
  AOI22_X1 U450 ( .A1(n510), .A2(mepc_i[29]), .B1(n627), .B2(n478), .ZN(n482)
         );
  AOI22_X1 U451 ( .A1(n507), .A2(boot_addr_i[28]), .B1(n479), .B2(
        m_trap_base_addr_i[21]), .ZN(n481) );
  NAND4_X1 U452 ( .A1(n484), .A2(n483), .A3(n482), .A4(n481), .ZN(n318) );
  NAND2_X1 U453 ( .A1(n485), .A2(boot_addr_i[29]), .ZN(n488) );
  NAND2_X1 U454 ( .A1(n626), .A2(mepc_i[30]), .ZN(n486) );
  AND3_X1 U455 ( .A1(n487), .A2(n488), .A3(n486), .ZN(n495) );
  AOI22_X1 U456 ( .A1(n509), .A2(m_trap_base_addr_i[22]), .B1(n472), .B2(
        u_trap_base_addr_i[22]), .ZN(n494) );
  HA_X1 U457 ( .A(n489), .B(pc_id_o[29]), .CO(n498), .S(n478) );
  AOI22_X1 U458 ( .A1(n471), .A2(jump_target_ex_i[30]), .B1(n501), .B2(n490), 
        .ZN(n493) );
  AOI22_X1 U459 ( .A1(n432), .A2(depc_i[30]), .B1(n451), .B2(uepc_i[30]), .ZN(
        n492) );
  NAND4_X1 U460 ( .A1(n495), .A2(n494), .A3(n493), .A4(n492), .ZN(n317) );
  NAND2_X1 U461 ( .A1(n496), .A2(uepc_i[31]), .ZN(n504) );
  NAND2_X1 U462 ( .A1(n497), .A2(u_trap_base_addr_i[23]), .ZN(n503) );
  HA_X1 U463 ( .A(n498), .B(pc_id_o[30]), .CO(n499), .S(n490) );
  XOR2_X1 U464 ( .A(n499), .B(pc_id_o[31]), .Z(n500) );
  NAND2_X1 U465 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND3_X1 U466 ( .A1(n502), .A2(n503), .A3(n504), .ZN(n514) );
  AOI22_X1 U467 ( .A1(n506), .A2(depc_i[31]), .B1(n505), .B2(
        jump_target_ex_i[31]), .ZN(n513) );
  AOI22_X1 U468 ( .A1(n508), .A2(jump_target_id_i[31]), .B1(n480), .B2(
        boot_addr_i[30]), .ZN(n512) );
  AOI22_X1 U469 ( .A1(n510), .A2(mepc_i[31]), .B1(n509), .B2(
        m_trap_base_addr_i[23]), .ZN(n511) );
  NAND4_X1 U470 ( .A1(n514), .A2(n513), .A3(n512), .A4(n511), .ZN(n316) );
  INV_X1 U471 ( .A(branch_req), .ZN(n515) );
  NAND2_X1 U472 ( .A1(fetch_valid), .A2(n515), .ZN(perf_imiss_o) );
  SDFFS_X1 offset_fsm_cs_reg_0_ ( .D(offset_fsm_ns_0_), .SI(1'b0), .SE(1'b0), 
        .CK(clk), .SN(rst_n), .Q(offset_fsm_cs_0_), .QN(n561) );
  SDFFR_X1 hwlp_dec_cnt_id_o_reg_0_ ( .D(n315), .SI(1'b0), .SE(1'b0), .CK(n774), .RN(rst_n), .Q(hwlp_dec_cnt_id_o[0]) );
  SDFFR_X1 instr_rdata_id_o_reg_2_ ( .D(instr_decompressed[2]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[2]) );
  SDFFR_X1 instr_rdata_id_o_reg_4_ ( .D(instr_decompressed[4]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[4]) );
  SDFFR_X1 instr_rdata_id_o_reg_5_ ( .D(instr_decompressed[5]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[5]) );
  SDFFR_X1 instr_rdata_id_o_reg_6_ ( .D(instr_decompressed[6]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[6]) );
  SDFFR_X1 instr_rdata_id_o_reg_7_ ( .D(instr_decompressed[7]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[7]) );
  SDFFR_X1 instr_rdata_id_o_reg_8_ ( .D(instr_decompressed[8]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[8]) );
  SDFFR_X1 instr_rdata_id_o_reg_9_ ( .D(instr_decompressed[9]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[9]) );
  SDFFR_X1 instr_rdata_id_o_reg_10_ ( .D(instr_decompressed[10]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[10]) );
  SDFFR_X1 instr_rdata_id_o_reg_11_ ( .D(instr_decompressed[11]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[11]) );
  SDFFR_X1 instr_rdata_id_o_reg_14_ ( .D(instr_decompressed[14]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[14]) );
  SDFFR_X1 instr_rdata_id_o_reg_22_ ( .D(instr_decompressed[22]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[22]) );
  SDFFR_X1 instr_rdata_id_o_reg_23_ ( .D(instr_decompressed[23]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[23]) );
  SDFFR_X1 instr_rdata_id_o_reg_24_ ( .D(instr_decompressed[24]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[24]) );
  SDFFR_X1 illegal_c_insn_id_o_reg ( .D(illegal_c_insn), .SI(1'b0), .SE(1'b0), 
        .CK(n774), .RN(rst_n), .Q(illegal_c_insn_id_o) );
  SDFFR_X1 is_compressed_id_o_reg ( .D(instr_compressed_int), .SI(1'b0), .SE(
        1'b0), .CK(n774), .RN(rst_n), .Q(is_compressed_id_o) );
  SDFFR_X1 pc_id_o_reg_0_ ( .D(pc_if_o[0]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[0]) );
  SDFFR_X1 pc_id_o_reg_1_ ( .D(pc_if_o[1]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[1]) );
  SDFFR_X1 pc_id_o_reg_3_ ( .D(pc_if_o[3]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[3]), .QN(n30) );
  SDFFR_X1 pc_id_o_reg_5_ ( .D(pc_if_o[5]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[5]), .QN(n587) );
  SDFFR_X1 pc_id_o_reg_6_ ( .D(pc_if_o[6]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[6]), .QN(n593) );
  SDFFR_X1 pc_id_o_reg_7_ ( .D(pc_if_o[7]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[7]), .QN(n589) );
  SDFFR_X1 pc_id_o_reg_9_ ( .D(pc_if_o[9]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[9]), .QN(n31) );
  SDFFR_X1 pc_id_o_reg_11_ ( .D(pc_if_o[11]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[11]), .QN(n32) );
  SDFFR_X1 pc_id_o_reg_12_ ( .D(pc_if_o[12]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[12]), .QN(n592) );
  SDFFR_X1 pc_id_o_reg_13_ ( .D(pc_if_o[13]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[13]), .QN(n33) );
  SDFFR_X1 pc_id_o_reg_14_ ( .D(pc_if_o[14]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[14]), .QN(n34) );
  SDFFR_X1 pc_id_o_reg_15_ ( .D(pc_if_o[15]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[15]), .QN(n35) );
  SDFFR_X1 pc_id_o_reg_16_ ( .D(pc_if_o[16]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[16]), .QN(n590) );
  SDFFR_X1 pc_id_o_reg_17_ ( .D(pc_if_o[17]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[17]), .QN(n586) );
  SDFFR_X1 pc_id_o_reg_18_ ( .D(pc_if_o[18]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[18]), .QN(n591) );
  SDFFR_X1 pc_id_o_reg_19_ ( .D(pc_if_o[19]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[19]), .QN(n585) );
  SDFFR_X1 pc_id_o_reg_21_ ( .D(pc_if_o[21]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[21]), .QN(n584) );
  SDFFR_X1 pc_id_o_reg_22_ ( .D(pc_if_o[22]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[22]), .QN(n594) );
  SDFFR_X1 pc_id_o_reg_23_ ( .D(pc_if_o[23]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[23]), .QN(n595) );
  SDFFR_X1 pc_id_o_reg_24_ ( .D(pc_if_o[24]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[24]) );
  SDFFR_X1 pc_id_o_reg_25_ ( .D(pc_if_o[25]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[25]) );
  SDFFR_X1 pc_id_o_reg_26_ ( .D(pc_if_o[26]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[26]) );
  SDFFR_X1 pc_id_o_reg_28_ ( .D(pc_if_o[28]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[28]) );
  SDFFR_X1 pc_id_o_reg_29_ ( .D(pc_if_o[29]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[29]) );
  SDFFR_X1 pc_id_o_reg_30_ ( .D(pc_if_o[30]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[30]) );
  SDFFR_X1 pc_id_o_reg_31_ ( .D(pc_if_o[31]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[31]) );
  SDFFR_X1 instr_rdata_id_o_reg_0_ ( .D(instr_decompressed[1]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[0]) );
  SDFFR_X1 instr_valid_id_o_reg ( .D(n247), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(rst_n), .Q(instr_valid_id_o), .QN(n611) );
  SDFFR_X1 is_hwlp_id_q_reg ( .D(fetch_is_hwlp), .SI(1'b0), .SE(1'b0), .CK(
        n774), .RN(rst_n), .Q(is_hwlp_id_q) );
  SDFFR_X1 hwlp_dec_cnt_if_reg_0_ ( .D(n246), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(rst_n), .QN(n599) );
  SDFFR_X1 hwlp_dec_cnt_if_reg_1_ ( .D(n245), .SI(1'b0), .SE(1'b0), .CK(clk), 
        .RN(rst_n), .QN(n600) );
  SDFFR_X1 hwlp_dec_cnt_id_o_reg_1_ ( .D(n243), .SI(1'b0), .SE(1'b0), .CK(n774), .RN(rst_n), .Q(hwlp_dec_cnt_id_o[1]) );
  SDFFR_X1 instr_rdata_id_o_reg_30_ ( .D(instr_decompressed[30]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[30]) );
  SDFFR_X1 pc_id_o_reg_27_ ( .D(pc_if_o[27]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[27]) );
  SDFFR_X1 pc_id_o_reg_8_ ( .D(pc_if_o[8]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[8]), .QN(n575) );
  SDFFR_X1 pc_id_o_reg_10_ ( .D(pc_if_o[10]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[10]), .QN(n574) );
  SDFFR_X1 pc_id_o_reg_4_ ( .D(pc_if_o[4]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[4]), .QN(n572) );
  SDFFR_X1 instr_rdata_id_o_reg_20_ ( .D(instr_decompressed[20]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[20]) );
  SDFFR_X1 instr_rdata_id_o_reg_27_ ( .D(instr_decompressed[27]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[27]) );
  SDFFR_X1 instr_rdata_id_o_reg_28_ ( .D(instr_decompressed[28]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[28]) );
  SDFFR_X1 instr_rdata_id_o_reg_21_ ( .D(instr_decompressed[21]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[21]) );
  SDFFR_X1 instr_rdata_id_o_reg_3_ ( .D(instr_decompressed[3]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[3]) );
  SDFFR_X1 pc_id_o_reg_2_ ( .D(pc_if_o[2]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[2]), .QN(n567) );
  SDFFR_X1 pc_id_o_reg_20_ ( .D(pc_if_o[20]), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .RN(rst_n), .Q(pc_id_o[20]), .QN(n573) );
  SDFFS_X1 instr_rdata_id_o_reg_1_ ( .D(n773), .SI(1'b0), .SE(1'b0), .CK(n774), 
        .SN(rst_n), .QN(instr_rdata_id_o[1]) );
  SDFFR_X1 instr_rdata_id_o_reg_15_ ( .D(instr_decompressed[15]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[15]) );
  SDFFR_X1 instr_rdata_id_o_reg_18_ ( .D(instr_decompressed[18]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[18]) );
  SDFFR_X1 instr_rdata_id_o_reg_19_ ( .D(instr_decompressed[19]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[19]) );
  SDFFR_X1 instr_rdata_id_o_reg_17_ ( .D(instr_decompressed[17]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[17]) );
  SDFFR_X2 instr_rdata_id_o_reg_31_ ( .D(instr_decompressed[31]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[31]) );
  SDFFR_X2 instr_rdata_id_o_reg_29_ ( .D(instr_decompressed[29]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[29]) );
  CLKBUF_X3 U260 ( .A(n167), .Z(n472) );
  riscv_prefetch_L0_buffer prefetch_128_prefetch_buffer_i ( .clk(clk), .rst_n(
        rst_n), .req_i(1'b1), .branch_i(branch_req), .addr_i({n316, n317, n318, 
        n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
        n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
        n343, n344, n345, n346, 1'b0}), .hwloop_i(hwlp_jump), 
        .hwloop_target_i(hwlp_target), .ready_i(fetch_ready), .valid_o(
        fetch_valid), .rdata_o(fetch_rdata), .addr_o(pc_if_o), .is_hwlp_o(
        fetch_is_hwlp), .instr_req_o(instr_req_o), .instr_addr_o({
        instr_addr_o[31:4], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3}), .instr_gnt_i(
        instr_gnt_i), .instr_rvalid_i(instr_rvalid_i), .instr_rdata_i(
        instr_rdata_i), .busy_o(if_busy_o) );
  riscv_hwloop_controller_N_REGS2 hwloop_controller_i ( .current_pc_i(pc_if_o), 
        .hwlp_start_addr_i(hwlp_start_i), .hwlp_end_addr_i(hwlp_end_i), 
        .hwlp_counter_i(hwlp_cnt_i), .hwlp_dec_cnt_id_i({n_2_net__1_, 
        n_2_net__0_}), .hwlp_jump_o(hwlp_jump), .hwlp_targ_addr_o(hwlp_target), 
        .hwlp_dec_cnt_o_1_(n9), .hwlp_dec_cnt_o_0_(n10) );
  riscv_compressed_decoder_FPU0 compressed_decoder_i ( .instr_i(fetch_rdata), 
        .instr_o({instr_decompressed, SYNOPSYS_UNCONNECTED__4}), 
        .is_compressed_o(instr_compressed_int), .illegal_instr_o(
        illegal_c_insn) );
  SNPS_CLOCK_GATE_HIGH_riscv_if_stage_2_128_0_1a110800_0 clk_gate_instr_rdata_id_o_reg_17_ ( 
        .CLK(clk), .EN(n555), .ENCLK(n774), .TE(1'b0) );
  SDFFR_X1 instr_rdata_id_o_reg_16_ ( .D(instr_decompressed[16]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[16]) );
  SDFFR_X2 instr_rdata_id_o_reg_25_ ( .D(instr_decompressed[25]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[25]) );
  SDFFR_X1 instr_rdata_id_o_reg_26_ ( .D(instr_decompressed[26]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[26]) );
  SDFFR_X2 instr_rdata_id_o_reg_12_ ( .D(instr_decompressed[12]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[12]) );
  SDFFR_X2 instr_rdata_id_o_reg_13_ ( .D(instr_decompressed[13]), .SI(1'b0), 
        .SE(1'b0), .CK(n774), .RN(rst_n), .Q(instr_rdata_id_o[13]) );
  CLKBUF_X1 U5 ( .A(pc_set_i), .Z(n7) );
  AND3_X1 U3 ( .A1(n461), .A2(n621), .A3(n620), .ZN(n470) );
  NAND2_X1 U7 ( .A1(n471), .A2(jump_target_ex_i[28]), .ZN(n620) );
  NAND2_X1 U10 ( .A1(n432), .A2(depc_i[28]), .ZN(n621) );
  BUF_X2 U14 ( .A(n133), .Z(n510) );
  BUF_X2 U18 ( .A(n133), .Z(n463) );
  CLKBUF_X1 U48 ( .A(n472), .Z(n368) );
  NAND2_X1 U55 ( .A1(n625), .A2(n366), .ZN(n367) );
  NAND2_X1 U56 ( .A1(n496), .A2(uepc_i[19]), .ZN(n625) );
  BUF_X1 U57 ( .A(n87), .Z(n466) );
  CLKBUF_X1 U58 ( .A(n480), .Z(n6) );
  BUF_X2 U99 ( .A(n174), .Z(n509) );
  BUF_X2 U101 ( .A(n133), .Z(n626) );
  CLKBUF_X1 U112 ( .A(pc_mux_i[0]), .Z(n377) );
  BUF_X2 U113 ( .A(n87), .Z(n627) );
  BUF_X2 U133 ( .A(n204), .Z(n507) );
  INV_X1 U138 ( .A(instr_decompressed[1]), .ZN(n773) );
  NAND2_X1 U147 ( .A1(n13), .A2(n375), .ZN(n328) );
endmodule


module cluster_clock_gating ( clk_i, en_i, test_en_i, clk_o );
  input clk_i, en_i, test_en_i;
  output clk_o;


  CLKGATETST_X1 cgc ( .CK(clk_i), .E(en_i), .SE(test_en_i), .GCK(clk_o) );
endmodule


module riscv_core_0_128_1_16_1_1_0_0_0_0_0_0_0_0_0_3_6_15_5_1a110800 ( clk_i, 
        rst_ni, clock_en_i, test_en_i, fregfile_disable_i, boot_addr_i, 
        core_id_i, cluster_id_i, instr_req_o, instr_gnt_i, instr_rvalid_i, 
        instr_addr_o, instr_rdata_i, data_req_o, data_gnt_i, data_rvalid_i, 
        data_we_o, data_be_o, data_addr_o, data_wdata_o, data_rdata_i, 
        apu_master_req_o, apu_master_ready_o, apu_master_gnt_i, 
        apu_master_operands_o, apu_master_op_o, apu_master_type_o, 
        apu_master_flags_o, apu_master_valid_i, apu_master_result_i, 
        apu_master_flags_i, irq_i, irq_id_i, irq_ack_o, irq_id_o, irq_sec_i, 
        sec_lvl_o, debug_req_i, fetch_enable_i, core_busy_o, 
        ext_perf_counters_i, test_mode_tp );
  input [31:0] boot_addr_i;
  input [3:0] core_id_i;
  input [5:0] cluster_id_i;
  output [31:0] instr_addr_o;
  input [127:0] instr_rdata_i;
  output [3:0] data_be_o;
  output [31:0] data_addr_o;
  output [31:0] data_wdata_o;
  input [31:0] data_rdata_i;
  output [95:0] apu_master_operands_o;
  output [5:0] apu_master_op_o;
  output [1:2] apu_master_type_o;
  output [14:0] apu_master_flags_o;
  input [31:0] apu_master_result_i;
  input [4:0] apu_master_flags_i;
  input [4:0] irq_id_i;
  output [4:0] irq_id_o;
  input [1:2] ext_perf_counters_i;
  input clk_i, rst_ni, clock_en_i, test_en_i, fregfile_disable_i, instr_gnt_i,
         instr_rvalid_i, data_gnt_i, data_rvalid_i, apu_master_gnt_i,
         apu_master_valid_i, irq_i, irq_sec_i, debug_req_i, fetch_enable_i,
         test_mode_tp;
  output instr_req_o, data_req_o, data_we_o, apu_master_req_o,
         apu_master_ready_o, irq_ack_o, sec_lvl_o, core_busy_o;
  wire   n316, n317, n318, n319, n332, core_ctrl_firstfetch, core_busy_q,
         data_load_event_ex, if_busy, core_busy_int, ctrl_busy, lsu_busy,
         clock_en, clk, trap_addr_mux, instr_req_int, instr_req_pmp,
         instr_gnt_pmp, is_hwlp_id, instr_valid_id, is_compressed_id,
         illegal_c_insn_id, clear_instr_valid, pc_set, halt_if, id_ready,
         perf_imiss, is_decoding, branch_in_ex, branch_decision, ex_ready,
         lsu_ready_wb, id_valid, ex_valid, alu_en_ex, alu_is_clpx_ex,
         alu_is_subrot_ex, regfile_we_ex, regfile_alu_we_ex, mult_en_ex,
         mult_sel_subword_ex, mult_is_clpx_ex, mult_clpx_img_ex, csr_access_ex,
         csr_irq_sec, csr_save_if, csr_save_id, csr_save_ex,
         csr_restore_mret_id, csr_restore_uret_id, csr_restore_dret_id,
         csr_save_cause, csr_hwlp_regid_0_, data_req_ex, data_we_ex,
         data_sign_ext_ex_0_, data_misaligned_ex, useincr_addr_ex,
         data_misaligned, data_err_pmp, data_err_ack, m_irq_enable,
         u_irq_enable, debug_csr_save, debug_single_step, debug_ebreakm,
         debug_ebreaku, regfile_we_wb, regfile_alu_we_fw, mult_multicycle,
         perf_jump, perf_jr_stall, perf_ld_stall, perf_pipeline_stall,
         lsu_ready_ex, data_req_pmp, data_gnt_pmp, n_0_net_, n_1_net_, n255,
         n256, n257, n258, n259, n260, n261, n262, n270, n271, n273, n276,
         n278, n280, n282, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n308, n309, n310,
         n311, n312, n313, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351;
  wire   [23:0] mtvec;
  wire   [23:0] utvec;
  wire   [31:4] instr_addr_pmp;
  wire   [1:0] hwlp_dec_cnt_id;
  wire   [31:0] instr_rdata_id;
  wire   [31:0] pc_if;
  wire   [31:0] pc_id;
  wire   [31:1] mepc;
  wire   [31:1] uepc;
  wire   [31:1] depc;
  wire   [2:0] pc_mux_id;
  wire   [1:0] exc_pc_mux_id;
  wire   [4:0] exc_cause;
  wire   [63:0] hwlp_start;
  wire   [63:0] hwlp_end;
  wire   [63:0] hwlp_cnt;
  wire   [31:1] jump_target_id;
  wire   [31:1] jump_target_ex;
  wire   [31:0] pc_ex;
  wire   [6:0] alu_operator_ex;
  wire   [31:0] alu_operand_a_ex;
  wire   [31:0] alu_operand_b_ex;
  wire   [31:0] alu_operand_c_ex;
  wire   [4:0] bmask_a_ex;
  wire   [4:0] bmask_b_ex;
  wire   [1:0] imm_vec_ext_ex;
  wire   [1:0] alu_vec_mode_ex;
  wire   [1:0] alu_clpx_shift_ex;
  wire   [4:0] regfile_waddr_ex;
  wire   [4:0] regfile_alu_waddr_ex;
  wire   [2:0] mult_operator_ex;
  wire   [1:0] mult_signed_mode_ex;
  wire   [31:0] mult_operand_a_ex;
  wire   [31:0] mult_operand_b_ex;
  wire   [31:0] mult_operand_c_ex;
  wire   [4:0] mult_imm_ex;
  wire   [31:0] mult_dot_op_a_ex;
  wire   [31:0] mult_dot_op_b_ex;
  wire   [31:0] mult_dot_op_c_ex;
  wire   [1:0] mult_dot_signed_ex;
  wire   [1:0] mult_clpx_shift_ex;
  wire   [1:0] csr_op_ex;
  wire   [1:0] current_priv_lvl;
  wire   [5:0] csr_cause;
  wire   [2:0] csr_hwlp_we;
  wire   [31:0] csr_hwlp_data;
  wire   [1:0] data_type_ex;
  wire   [2:1] debug_cause;
  wire   [4:0] regfile_waddr_fw_wb_o;
  wire   [31:0] regfile_wdata;
  wire   [4:0] regfile_alu_waddr_fw;
  wire   [31:0] regfile_alu_wdata_fw;
  wire   [31:0] lsu_rdata;
  wire   [31:0] csr_rdata;
  wire   [31:0] data_addr_pmp;
  wire   [11:0] csr_addr;
  wire   [511:0] pmp_addr;
  wire   [79:0] pmp_cfg;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64;
  assign apu_master_ready_o = 1'b1;
  assign apu_master_flags_o[0] = 1'b0;
  assign apu_master_flags_o[1] = 1'b0;
  assign apu_master_flags_o[2] = 1'b0;
  assign apu_master_flags_o[3] = 1'b0;
  assign apu_master_flags_o[4] = 1'b0;
  assign apu_master_flags_o[5] = 1'b0;
  assign apu_master_flags_o[6] = 1'b0;
  assign apu_master_flags_o[7] = 1'b0;
  assign apu_master_flags_o[8] = 1'b0;
  assign apu_master_flags_o[9] = 1'b0;
  assign apu_master_flags_o[10] = 1'b0;
  assign apu_master_flags_o[11] = 1'b0;
  assign apu_master_flags_o[12] = 1'b0;
  assign apu_master_flags_o[13] = 1'b0;
  assign apu_master_flags_o[14] = 1'b0;
  assign apu_master_type_o[2] = 1'b0;
  assign apu_master_type_o[1] = 1'b0;
  assign apu_master_op_o[0] = 1'b0;
  assign apu_master_op_o[1] = 1'b0;
  assign apu_master_op_o[2] = 1'b0;
  assign apu_master_op_o[3] = 1'b0;
  assign apu_master_op_o[4] = 1'b0;
  assign apu_master_op_o[5] = 1'b0;
  assign apu_master_operands_o[0] = 1'b0;
  assign apu_master_operands_o[1] = 1'b0;
  assign apu_master_operands_o[2] = 1'b0;
  assign apu_master_operands_o[3] = 1'b0;
  assign apu_master_operands_o[4] = 1'b0;
  assign apu_master_operands_o[5] = 1'b0;
  assign apu_master_operands_o[6] = 1'b0;
  assign apu_master_operands_o[7] = 1'b0;
  assign apu_master_operands_o[8] = 1'b0;
  assign apu_master_operands_o[9] = 1'b0;
  assign apu_master_operands_o[10] = 1'b0;
  assign apu_master_operands_o[11] = 1'b0;
  assign apu_master_operands_o[12] = 1'b0;
  assign apu_master_operands_o[13] = 1'b0;
  assign apu_master_operands_o[14] = 1'b0;
  assign apu_master_operands_o[15] = 1'b0;
  assign apu_master_operands_o[16] = 1'b0;
  assign apu_master_operands_o[17] = 1'b0;
  assign apu_master_operands_o[18] = 1'b0;
  assign apu_master_operands_o[19] = 1'b0;
  assign apu_master_operands_o[20] = 1'b0;
  assign apu_master_operands_o[21] = 1'b0;
  assign apu_master_operands_o[22] = 1'b0;
  assign apu_master_operands_o[23] = 1'b0;
  assign apu_master_operands_o[24] = 1'b0;
  assign apu_master_operands_o[25] = 1'b0;
  assign apu_master_operands_o[26] = 1'b0;
  assign apu_master_operands_o[27] = 1'b0;
  assign apu_master_operands_o[28] = 1'b0;
  assign apu_master_operands_o[29] = 1'b0;
  assign apu_master_operands_o[30] = 1'b0;
  assign apu_master_operands_o[31] = 1'b0;
  assign apu_master_operands_o[32] = 1'b0;
  assign apu_master_operands_o[33] = 1'b0;
  assign apu_master_operands_o[34] = 1'b0;
  assign apu_master_operands_o[35] = 1'b0;
  assign apu_master_operands_o[36] = 1'b0;
  assign apu_master_operands_o[37] = 1'b0;
  assign apu_master_operands_o[38] = 1'b0;
  assign apu_master_operands_o[39] = 1'b0;
  assign apu_master_operands_o[40] = 1'b0;
  assign apu_master_operands_o[41] = 1'b0;
  assign apu_master_operands_o[42] = 1'b0;
  assign apu_master_operands_o[43] = 1'b0;
  assign apu_master_operands_o[44] = 1'b0;
  assign apu_master_operands_o[45] = 1'b0;
  assign apu_master_operands_o[46] = 1'b0;
  assign apu_master_operands_o[47] = 1'b0;
  assign apu_master_operands_o[48] = 1'b0;
  assign apu_master_operands_o[49] = 1'b0;
  assign apu_master_operands_o[50] = 1'b0;
  assign apu_master_operands_o[51] = 1'b0;
  assign apu_master_operands_o[52] = 1'b0;
  assign apu_master_operands_o[53] = 1'b0;
  assign apu_master_operands_o[54] = 1'b0;
  assign apu_master_operands_o[55] = 1'b0;
  assign apu_master_operands_o[56] = 1'b0;
  assign apu_master_operands_o[57] = 1'b0;
  assign apu_master_operands_o[58] = 1'b0;
  assign apu_master_operands_o[59] = 1'b0;
  assign apu_master_operands_o[60] = 1'b0;
  assign apu_master_operands_o[61] = 1'b0;
  assign apu_master_operands_o[62] = 1'b0;
  assign apu_master_operands_o[63] = 1'b0;
  assign apu_master_operands_o[64] = 1'b0;
  assign apu_master_operands_o[65] = 1'b0;
  assign apu_master_operands_o[66] = 1'b0;
  assign apu_master_operands_o[67] = 1'b0;
  assign apu_master_operands_o[68] = 1'b0;
  assign apu_master_operands_o[69] = 1'b0;
  assign apu_master_operands_o[70] = 1'b0;
  assign apu_master_operands_o[71] = 1'b0;
  assign apu_master_operands_o[72] = 1'b0;
  assign apu_master_operands_o[73] = 1'b0;
  assign apu_master_operands_o[74] = 1'b0;
  assign apu_master_operands_o[75] = 1'b0;
  assign apu_master_operands_o[76] = 1'b0;
  assign apu_master_operands_o[77] = 1'b0;
  assign apu_master_operands_o[78] = 1'b0;
  assign apu_master_operands_o[79] = 1'b0;
  assign apu_master_operands_o[80] = 1'b0;
  assign apu_master_operands_o[81] = 1'b0;
  assign apu_master_operands_o[82] = 1'b0;
  assign apu_master_operands_o[83] = 1'b0;
  assign apu_master_operands_o[84] = 1'b0;
  assign apu_master_operands_o[85] = 1'b0;
  assign apu_master_operands_o[86] = 1'b0;
  assign apu_master_operands_o[87] = 1'b0;
  assign apu_master_operands_o[88] = 1'b0;
  assign apu_master_operands_o[89] = 1'b0;
  assign apu_master_operands_o[90] = 1'b0;
  assign apu_master_operands_o[91] = 1'b0;
  assign apu_master_operands_o[92] = 1'b0;
  assign apu_master_operands_o[93] = 1'b0;
  assign apu_master_operands_o[94] = 1'b0;
  assign apu_master_operands_o[95] = 1'b0;
  assign apu_master_req_o = 1'b0;
  assign instr_addr_o[0] = 1'b0;
  assign instr_addr_o[1] = 1'b0;
  assign instr_addr_o[2] = 1'b0;
  assign instr_addr_o[3] = 1'b0;
  assign instr_addr_o[18] = n316;
  assign instr_addr_o[14] = n317;
  assign instr_addr_o[4] = n318;
  assign data_addr_o[31] = n319;

  CLKBUF_X1 U27 ( .A(alu_operand_a_ex[16]), .Z(n313) );
  AND2_X1 U33 ( .A1(n351), .A2(alu_operand_b_ex[10]), .ZN(csr_addr[10]) );
  AND2_X1 U34 ( .A1(n351), .A2(alu_operand_b_ex[0]), .ZN(csr_addr[0]) );
  AND2_X1 U35 ( .A1(n351), .A2(alu_operand_b_ex[3]), .ZN(csr_addr[3]) );
  AND2_X1 U36 ( .A1(n351), .A2(alu_operand_b_ex[2]), .ZN(csr_addr[2]) );
  AND2_X1 U37 ( .A1(n351), .A2(alu_operand_b_ex[11]), .ZN(csr_addr[11]) );
  CLKBUF_X1 U39 ( .A(branch_decision), .Z(n308) );
  OR2_X1 U40 ( .A1(core_ctrl_firstfetch), .A2(core_busy_q), .ZN(core_busy_o)
         );
  OR2_X1 U41 ( .A1(clock_en_i), .A2(core_busy_o), .ZN(clock_en) );
  INV_X1 U42 ( .A(n332), .ZN(irq_ack_o) );
  AND2_X1 U44 ( .A1(n351), .A2(alu_operand_b_ex[6]), .ZN(csr_addr[6]) );
  AND2_X1 U45 ( .A1(n351), .A2(alu_operand_b_ex[5]), .ZN(csr_addr[5]) );
  AND2_X1 U46 ( .A1(n351), .A2(alu_operand_b_ex[7]), .ZN(csr_addr[7]) );
  AND2_X1 U47 ( .A1(n351), .A2(alu_operand_b_ex[4]), .ZN(csr_addr[4]) );
  AND2_X1 U48 ( .A1(n351), .A2(alu_operand_b_ex[8]), .ZN(csr_addr[8]) );
  AND2_X1 U49 ( .A1(n351), .A2(n350), .ZN(csr_addr[9]) );
  NOR2_X1 U50 ( .A1(ctrl_busy), .A2(lsu_busy), .ZN(n309) );
  AOI21_X1 U51 ( .B1(data_req_o), .B2(data_load_event_ex), .A(n309), .ZN(n310)
         );
  OR2_X1 U52 ( .A1(if_busy), .A2(n310), .ZN(core_busy_int) );
  INV_X1 U53 ( .A(data_we_o), .ZN(n311) );
  AND3_X1 U54 ( .A1(data_req_o), .A2(data_gnt_i), .A3(n311), .ZN(n_0_net_) );
  AND3_X1 U55 ( .A1(data_req_o), .A2(data_we_o), .A3(data_gnt_i), .ZN(n_1_net_) );
  SDFFR_X1 core_busy_q_reg ( .D(core_busy_int), .SI(1'b0), .SE(1'b0), .CK(
        clk_i), .RN(rst_ni), .Q(core_busy_q) );
  cluster_clock_gating core_clock_gate_i ( .clk_i(clk_i), .en_i(clock_en), 
        .test_en_i(test_en_i), .clk_o(clk) );
  riscv_if_stage_2_128_0_1a110800 if_stage_i ( .clk(clk), .rst_n(rst_ni), 
        .m_trap_base_addr_i(mtvec), .u_trap_base_addr_i(utvec), 
        .trap_addr_mux_i(trap_addr_mux), .boot_addr_i(boot_addr_i[31:1]), 
        .req_i(instr_req_int), .instr_req_o(instr_req_pmp), .instr_addr_o({
        instr_addr_pmp[31:21], n335, instr_addr_pmp[19:7], n336, 
        instr_addr_pmp[5:4], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3}), .instr_gnt_i(
        instr_gnt_pmp), .instr_rvalid_i(instr_rvalid_i), .instr_rdata_i(
        instr_rdata_i), .instr_err_pmp_i(1'b0), .hwlp_dec_cnt_id_o(
        hwlp_dec_cnt_id), .is_hwlp_id_o(is_hwlp_id), .instr_valid_id_o(
        instr_valid_id), .instr_rdata_id_o(instr_rdata_id), 
        .is_compressed_id_o(is_compressed_id), .illegal_c_insn_id_o(
        illegal_c_insn_id), .pc_if_o(pc_if), .pc_id_o(pc_id), 
        .clear_instr_valid_i(clear_instr_valid), .pc_set_i(pc_set), .mepc_i({
        mepc, 1'b0}), .uepc_i({uepc, 1'b0}), .depc_i({depc, 1'b0}), .pc_mux_i(
        pc_mux_id), .exc_pc_mux_i({1'b0, exc_pc_mux_id}), .exc_vec_pc_mux_i({
        n337, exc_cause[3:0]}), .jump_target_id_i({jump_target_id, 1'b0}), 
        .jump_target_ex_i({jump_target_ex, 1'b0}), .hwlp_start_i(hwlp_start), 
        .hwlp_end_i(hwlp_end), .hwlp_cnt_i(hwlp_cnt), .halt_if_i(halt_if), 
        .if_busy_o(if_busy), .perf_imiss_o(perf_imiss), .id_ready_i_BAR(
        id_ready) );
  riscv_id_stage_N_HWLP2_PULP_SECURE1_APU0_FPU0_Zfinx0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_MULT0_SHARED_INT_DIV0_SHARED_FP_DIVSQRT0_WAPUTYPE0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5 id_stage_i ( 
        .clk(clk), .rst_n(rst_ni), .test_en_i(1'b0), .fregfile_disable_i(1'b0), 
        .fetch_enable_i(fetch_enable_i), .ctrl_busy_o(ctrl_busy), 
        .core_ctrl_firstfetch_o(core_ctrl_firstfetch), .hwlp_dec_cnt_i(
        hwlp_dec_cnt_id), .is_hwlp_i(is_hwlp_id), .instr_valid_i(
        instr_valid_id), .instr_rdata_i(instr_rdata_id), .instr_req_o(
        instr_req_int), .branch_in_ex_o(branch_in_ex), .branch_decision_i(
        branch_decision), .jump_target_o({jump_target_id, 
        SYNOPSYS_UNCONNECTED__4}), .clear_instr_valid_o(clear_instr_valid), 
        .pc_set_o(pc_set), .pc_mux_o(pc_mux_id), .exc_pc_mux_o({
        SYNOPSYS_UNCONNECTED__5, exc_pc_mux_id}), .trap_addr_mux_o(
        trap_addr_mux), .illegal_c_insn_i(illegal_c_insn_id), 
        .is_compressed_i(is_compressed_id), .is_fetch_failed_i(1'b0), 
        .pc_if_i(pc_if), .pc_id_i(pc_id), .halt_if_o(halt_if), .ex_ready_i(
        ex_ready), .wb_ready_i(lsu_ready_wb), .id_valid_o(id_valid), 
        .ex_valid_i(ex_valid), .pc_ex_o(pc_ex), .alu_operand_a_ex_o(
        alu_operand_a_ex), .alu_operand_b_ex_o(alu_operand_b_ex), 
        .alu_operand_c_ex_o(alu_operand_c_ex), .bmask_a_ex_o(bmask_a_ex), 
        .bmask_b_ex_o(bmask_b_ex), .imm_vec_ext_ex_o(imm_vec_ext_ex), 
        .alu_vec_mode_ex_o(alu_vec_mode_ex), .regfile_waddr_ex_o({
        SYNOPSYS_UNCONNECTED__6, regfile_waddr_ex}), .regfile_we_ex_o(
        regfile_we_ex), .regfile_alu_waddr_ex_o({SYNOPSYS_UNCONNECTED__7, 
        regfile_alu_waddr_ex}), .alu_operator_ex_o(alu_operator_ex), 
        .alu_is_clpx_ex_o(alu_is_clpx_ex), .alu_is_subrot_ex_o(
        alu_is_subrot_ex), .alu_clpx_shift_ex_o(alu_clpx_shift_ex), 
        .mult_operator_ex_o(mult_operator_ex), .mult_operand_a_ex_o(
        mult_operand_a_ex), .mult_operand_b_ex_o(mult_operand_b_ex), 
        .mult_operand_c_ex_o(mult_operand_c_ex), .mult_en_ex_o(mult_en_ex), 
        .mult_signed_mode_ex_o(mult_signed_mode_ex), .mult_imm_ex_o(
        mult_imm_ex), .mult_dot_op_a_ex_o(mult_dot_op_a_ex), 
        .mult_dot_op_b_ex_o(mult_dot_op_b_ex), .mult_dot_op_c_ex_o(
        mult_dot_op_c_ex), .mult_dot_signed_ex_o(mult_dot_signed_ex), 
        .mult_is_clpx_ex_o(mult_is_clpx_ex), .mult_clpx_shift_ex_o(
        mult_clpx_shift_ex), .mult_clpx_img_ex_o(mult_clpx_img_ex), 
        .apu_read_dep_i(1'b0), .apu_write_dep_i(1'b0), .apu_busy_i(1'b0), 
        .frm_i({1'b0, 1'b0, 1'b0}), .csr_op_ex_o(csr_op_ex), 
        .current_priv_lvl_i(current_priv_lvl), .csr_irq_sec_o(csr_irq_sec), 
        .csr_save_if_o(csr_save_if), .csr_save_id_o(csr_save_id), 
        .csr_restore_mret_id_o(csr_restore_mret_id), .csr_restore_uret_id_o(
        csr_restore_uret_id), .csr_restore_dret_id_o(csr_restore_dret_id), 
        .csr_save_cause_o(csr_save_cause), .hwlp_start_o(hwlp_start), 
        .hwlp_end_o(hwlp_end), .hwlp_cnt_o(hwlp_cnt), .csr_hwlp_regid_i(
        csr_hwlp_regid_0_), .csr_hwlp_we_i(csr_hwlp_we), .csr_hwlp_data_i({
        csr_hwlp_data[31:13], n347, n346, csr_hwlp_data[10:5], n348, 
        csr_hwlp_data[3:0]}), .data_req_ex_o(data_req_ex), .data_we_ex_o(
        data_we_ex), .data_type_ex_o(data_type_ex), .data_sign_ext_ex_o({
        SYNOPSYS_UNCONNECTED__8, data_sign_ext_ex_0_}), .data_load_event_ex_o(
        data_load_event_ex), .data_misaligned_i(data_misaligned), .irq_i(irq_i), .irq_sec_i(irq_sec_i), .irq_id_i(irq_id_i), .m_irq_enable_i(m_irq_enable), 
        .u_irq_enable_i(u_irq_enable), .irq_id_o(irq_id_o), .exc_cause_o({
        SYNOPSYS_UNCONNECTED__9, n337, exc_cause[3:0]}), .debug_cause_o({
        debug_cause, SYNOPSYS_UNCONNECTED__10}), .debug_csr_save_o(
        debug_csr_save), .debug_req_i(debug_req_i), .debug_single_step_i(
        debug_single_step), .debug_ebreakm_i(debug_ebreakm), .debug_ebreaku_i(
        debug_ebreaku), .regfile_waddr_wb_i({1'b0, regfile_waddr_fw_wb_o}), 
        .regfile_we_wb_i(regfile_we_wb), .regfile_wdata_wb_i({
        regfile_wdata[31:24], n258, n256, regfile_wdata[21], n270, 
        regfile_wdata[19:15], n288, n295, n291, n293, n299, n297, n301, 
        regfile_wdata[7:0]}), .regfile_alu_waddr_fw_i({1'b0, 
        regfile_alu_waddr_fw}), .regfile_alu_we_fw_i(regfile_alu_we_fw), 
        .regfile_alu_wdata_fw_i({regfile_alu_wdata_fw[31], n342, n333, n343, 
        regfile_alu_wdata_fw[27:21], n341, regfile_alu_wdata_fw[19], n339, 
        regfile_alu_wdata_fw[17:13], n340, n262, regfile_alu_wdata_fw[10:8], 
        n334, n261, regfile_alu_wdata_fw[5], n260, regfile_alu_wdata_fw[3:2], 
        n345, n344}), .mult_multicycle_i(mult_multicycle), .perf_jump_o(
        perf_jump), .perf_jr_stall_o(perf_jr_stall), .perf_ld_stall_o(
        perf_ld_stall), .perf_pipeline_stall_o(perf_pipeline_stall), 
        .irq_ack_o_BAR(n332), .csr_cause_o_5__BAR(csr_cause[5]), 
        .csr_cause_o_4_(n338), .csr_cause_o_3_(csr_cause[3]), .csr_cause_o_2_(
        csr_cause[2]), .csr_cause_o_0_(csr_cause[0]), .id_ready_o_BAR(id_ready), .data_err_ack_o_BAR(data_err_ack), .csr_save_ex_o_BAR(csr_save_ex), 
        .data_err_i_BAR(data_err_pmp), .regfile_alu_we_ex_o(regfile_alu_we_ex), 
        .alu_en_ex_o_BAR(alu_en_ex), .mult_sel_subword_ex_o_BAR(
        mult_sel_subword_ex), .csr_cause_o_1__BAR(csr_cause[1]), 
        .is_decoding_o(is_decoding), .csr_access_ex_o_BAR(csr_access_ex), 
        .data_misaligned_ex_o_BAR(data_misaligned_ex), .prepost_useincr_ex_o(
        useincr_addr_ex) );
  riscv_ex_stage_FPU0_FP_DIVSQRT0_SHARED_FP0_SHARED_DSP_MULT0_SHARED_INT_DIV0_APU_NARGS_CPU3_APU_WOP_CPU6_APU_NDSFLAGS_CPU15_APU_NUSFLAGS_CPU5 ex_stage_i ( 
        .clk(clk), .rst_n(rst_ni), .alu_operator_i(alu_operator_ex), 
        .alu_operand_a_i(alu_operand_a_ex), .alu_operand_b_i(alu_operand_b_ex), 
        .alu_operand_c_i(alu_operand_c_ex), .bmask_a_i(bmask_a_ex), 
        .bmask_b_i(bmask_b_ex), .imm_vec_ext_i(imm_vec_ext_ex), 
        .alu_vec_mode_i(alu_vec_mode_ex), .alu_is_clpx_i(alu_is_clpx_ex), 
        .alu_is_subrot_i(alu_is_subrot_ex), .alu_clpx_shift_i(
        alu_clpx_shift_ex), .mult_operator_i(mult_operator_ex), 
        .mult_operand_a_i(mult_operand_a_ex), .mult_operand_b_i(
        mult_operand_b_ex), .mult_operand_c_i(mult_operand_c_ex), .mult_en_i(
        mult_en_ex), .mult_signed_mode_i(mult_signed_mode_ex), .mult_imm_i(
        mult_imm_ex), .mult_dot_op_a_i(mult_dot_op_a_ex), .mult_dot_op_b_i(
        mult_dot_op_b_ex), .mult_dot_op_c_i(mult_dot_op_c_ex), 
        .mult_dot_signed_i(mult_dot_signed_ex), .mult_is_clpx_i(
        mult_is_clpx_ex), .mult_clpx_shift_i(mult_clpx_shift_ex), 
        .mult_clpx_img_i(mult_clpx_img_ex), .mult_multicycle_o(mult_multicycle), .fpu_prec_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .apu_en_i(1'b0), .apu_op_i({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .apu_lat_i({1'b0, 1'b0}), 
        .apu_operands_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .apu_waddr_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .apu_flags_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .apu_read_regs_i({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .apu_read_regs_valid_i({1'b0, 1'b0, 1'b0}), 
        .apu_write_regs_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .apu_write_regs_valid_i({1'b0, 1'b0}), 
        .apu_master_gnt_i(1'b0), .apu_master_valid_i(1'b0), 
        .apu_master_result_i({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .lsu_en_i(data_req_ex), .lsu_rdata_i({lsu_rdata[31:24], n259, n257, 
        lsu_rdata[21], n271, lsu_rdata[19:15], n289, n296, n292, n294, n300, 
        n298, n302, lsu_rdata[7:0]}), .branch_in_ex_i(branch_in_ex), 
        .regfile_alu_waddr_i({1'b0, regfile_alu_waddr_ex}), .regfile_we_i(
        regfile_we_ex), .regfile_waddr_i({1'b0, regfile_waddr_ex}), 
        .csr_rdata_i(csr_rdata), .regfile_waddr_wb_o({SYNOPSYS_UNCONNECTED__11, 
        regfile_waddr_fw_wb_o}), .regfile_we_wb_o(regfile_we_wb), 
        .regfile_wdata_wb_o({regfile_wdata[31:24], n258, n256, 
        regfile_wdata[21], n270, regfile_wdata[19:15], n288, n295, n291, n293, 
        n299, n297, n301, regfile_wdata[7:0]}), .regfile_alu_waddr_fw_o({
        SYNOPSYS_UNCONNECTED__12, regfile_alu_waddr_fw}), 
        .regfile_alu_we_fw_o(regfile_alu_we_fw), .regfile_alu_wdata_fw_o({
        regfile_alu_wdata_fw[31], n342, n333, n343, 
        regfile_alu_wdata_fw[27:21], n341, regfile_alu_wdata_fw[19], n339, 
        regfile_alu_wdata_fw[17:13], n340, n262, regfile_alu_wdata_fw[10:8], 
        n334, n261, regfile_alu_wdata_fw[5], n260, regfile_alu_wdata_fw[3:2], 
        n345, n344}), .jump_target_o({jump_target_ex, SYNOPSYS_UNCONNECTED__13}), .branch_decision_o(branch_decision), .lsu_ready_ex_i(lsu_ready_ex), 
        .ex_ready_o(ex_ready), .ex_valid_o(ex_valid), .wb_ready_i(lsu_ready_wb), .lsu_err_i_BAR(data_err_pmp), .regfile_alu_we_i(regfile_alu_we_ex), 
        .alu_en_i_BAR(alu_en_ex), .mult_sel_subword_i_BAR(mult_sel_subword_ex), 
        .csr_access_i_BAR(csr_access_ex) );
  riscv_load_store_unit load_store_unit_i ( .clk(clk), .rst_n(rst_ni), 
        .data_req_o(data_req_pmp), .data_gnt_i(data_gnt_pmp), .data_rvalid_i(
        data_rvalid_i), .data_addr_o({data_addr_pmp[31:29], n280, n287, 
        data_addr_pmp[26:25], n276, data_addr_pmp[23], n273, n282, 
        data_addr_pmp[20], n278, data_addr_pmp[18:14], n290, 
        data_addr_pmp[12:0]}), .data_we_o(data_we_o), .data_be_o(data_be_o), 
        .data_wdata_o(data_wdata_o), .data_rdata_i(data_rdata_i), 
        .data_we_ex_i(data_we_ex), .data_type_ex_i(data_type_ex), 
        .data_wdata_ex_i(alu_operand_c_ex), .data_reg_offset_ex_i({1'b0, 1'b0}), .data_sign_ext_ex_i({1'b0, data_sign_ext_ex_0_}), .data_rdata_ex_o({
        lsu_rdata[31:24], n259, n257, lsu_rdata[21], n271, lsu_rdata[19:15], 
        n289, n296, n292, n294, n300, n298, n302, lsu_rdata[7:0]}), 
        .data_req_ex_i(data_req_ex), .operand_a_ex_i({n349, 
        alu_operand_a_ex[30:17], n313, n255, alu_operand_a_ex[14:10], n312, 
        alu_operand_a_ex[8:0]}), .operand_b_ex_i({alu_operand_b_ex[31:10], 
        n350, alu_operand_b_ex[8:0]}), .data_misaligned_o(data_misaligned), 
        .lsu_ready_ex_o(lsu_ready_ex), .lsu_ready_wb_o(lsu_ready_wb), 
        .ex_valid_i(ex_valid), .busy_o(lsu_busy), .data_err_i_BAR(data_err_pmp), .data_misaligned_ex_i_BAR(data_misaligned_ex), .addr_useincr_ex_i(
        useincr_addr_ex) );
  riscv_cs_registers_N_EXT_CNT0_APU0_FPU0_PULP_SECURE1_USE_PMP1_N_PMP_ENTRIES16 cs_registers_i ( 
        .clk(clk), .rst_n(rst_ni), .core_id_i(core_id_i), .cluster_id_i(
        cluster_id_i), .mtvec_o(mtvec), .utvec_o(utvec), .boot_addr_i({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .csr_addr_i(csr_addr), 
        .csr_wdata_i({n349, alu_operand_a_ex[30:17], n313, n255, 
        alu_operand_a_ex[14:10], n312, alu_operand_a_ex[8:0]}), .csr_op_i(
        csr_op_ex), .csr_rdata_o(csr_rdata), .fflags_i({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .fflags_we_i(1'b0), .m_irq_enable_o(m_irq_enable), 
        .u_irq_enable_o(u_irq_enable), .csr_irq_sec_i(csr_irq_sec), 
        .sec_lvl_o(sec_lvl_o), .mepc_o({mepc, SYNOPSYS_UNCONNECTED__14}), 
        .uepc_o({uepc, SYNOPSYS_UNCONNECTED__15}), .debug_mode_i(1'b0), 
        .debug_cause_i({debug_cause, 1'b0}), .debug_csr_save_i(debug_csr_save), 
        .depc_o({depc, SYNOPSYS_UNCONNECTED__16}), .debug_single_step_o(
        debug_single_step), .debug_ebreakm_o(debug_ebreakm), .debug_ebreaku_o(
        debug_ebreaku), .pmp_addr_o(pmp_addr), .pmp_cfg_o({
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, pmp_cfg[79:75], SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, pmp_cfg[74:70], 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, pmp_cfg[69:65], SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, pmp_cfg[64:60], 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, pmp_cfg[59:55], SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, pmp_cfg[54:50], 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, pmp_cfg[49:45], SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, pmp_cfg[44:40], 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, pmp_cfg[39:35], SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, pmp_cfg[34:30], 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, pmp_cfg[29:25], SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, pmp_cfg[24:20], 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, pmp_cfg[19:15], SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, pmp_cfg[14:10], 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, pmp_cfg[9:5], SYNOPSYS_UNCONNECTED__62, 
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, pmp_cfg[4:0]}), 
        .priv_lvl_o(current_priv_lvl), .pc_if_i(pc_if), .pc_id_i(pc_id), 
        .pc_ex_i(pc_ex), .csr_save_if_i(csr_save_if), .csr_save_id_i(
        csr_save_id), .csr_restore_mret_i(csr_restore_mret_id), 
        .csr_restore_uret_i(csr_restore_uret_id), .csr_restore_dret_i(
        csr_restore_dret_id), .csr_save_cause_i(csr_save_cause), 
        .hwlp_start_i(hwlp_start), .hwlp_end_i(hwlp_end), .hwlp_cnt_i(hwlp_cnt), .hwlp_data_o({csr_hwlp_data[31:13], n347, n346, csr_hwlp_data[10:5], n348, 
        csr_hwlp_data[3:0]}), .hwlp_regid_o(csr_hwlp_regid_0_), .hwlp_we_o(
        csr_hwlp_we), .id_valid_i(id_valid), .is_compressed_i(is_compressed_id), .imiss_i(perf_imiss), .pc_set_i(pc_set), .jump_i(perf_jump), .branch_i(
        branch_in_ex), .branch_taken_i(n308), .ld_stall_i(perf_ld_stall), 
        .jr_stall_i(perf_jr_stall), .pipeline_stall_i(perf_pipeline_stall), 
        .apu_typeconflict_i(1'b0), .apu_contention_i(1'b0), .apu_dep_i(1'b0), 
        .apu_wb_i(1'b0), .mem_load_i(n_0_net_), .mem_store_i(n_1_net_), 
        .ext_counters_i({1'b0, 1'b0}), .csr_cause_i_5__BAR(csr_cause[5]), 
        .csr_cause_i_4_(n338), .csr_cause_i_3_(csr_cause[3]), .csr_cause_i_2_(
        csr_cause[2]), .csr_cause_i_0_(csr_cause[0]), .csr_save_ex_i_BAR(
        csr_save_ex), .csr_cause_i_1__BAR(csr_cause[1]), .is_decoding_i(
        is_decoding), .csr_access_i_BAR(csr_access_ex) );
  riscv_pmp_N_PMP_ENTRIES16 RISCY_PMP_pmp_unit_i ( .clk(clk), .rst_n(rst_ni), 
        .pmp_privil_mode_i(current_priv_lvl), .pmp_addr_i(pmp_addr), 
        .pmp_cfg_i({1'b0, 1'b0, 1'b0, pmp_cfg[79:75], 1'b0, 1'b0, 1'b0, 
        pmp_cfg[74:70], 1'b0, 1'b0, 1'b0, pmp_cfg[69:65], 1'b0, 1'b0, 1'b0, 
        pmp_cfg[64:60], 1'b0, 1'b0, 1'b0, pmp_cfg[59:55], 1'b0, 1'b0, 1'b0, 
        pmp_cfg[54:50], 1'b0, 1'b0, 1'b0, pmp_cfg[49:45], 1'b0, 1'b0, 1'b0, 
        pmp_cfg[44:40], 1'b0, 1'b0, 1'b0, pmp_cfg[39:35], 1'b0, 1'b0, 1'b0, 
        pmp_cfg[34:30], 1'b0, 1'b0, 1'b0, pmp_cfg[29:25], 1'b0, 1'b0, 1'b0, 
        pmp_cfg[24:20], 1'b0, 1'b0, 1'b0, pmp_cfg[19:15], 1'b0, 1'b0, 1'b0, 
        pmp_cfg[14:10], 1'b0, 1'b0, 1'b0, pmp_cfg[9:5], 1'b0, 1'b0, 1'b0, 
        pmp_cfg[4:0]}), .data_req_i(data_req_pmp), .data_addr_i({
        data_addr_pmp[31:29], n280, n287, data_addr_pmp[26:25], n276, 
        data_addr_pmp[23], n273, n282, data_addr_pmp[20], n278, 
        data_addr_pmp[18:14], n290, data_addr_pmp[12:0]}), .data_we_i(
        data_we_o), .data_gnt_o(data_gnt_pmp), .data_req_o(data_req_o), 
        .data_gnt_i(data_gnt_i), .instr_req_i(instr_req_pmp), .instr_addr_i({
        instr_addr_pmp[31:21], n335, instr_addr_pmp[19:7], n336, 
        instr_addr_pmp[5:4], 1'b0, 1'b0, 1'b0, 1'b0}), .instr_gnt_o(
        instr_gnt_pmp), .instr_req_o(instr_req_o), .instr_gnt_i(instr_gnt_i), 
        .data_err_ack_i_BAR(data_err_ack), .data_err_o_BAR(data_err_pmp), 
        .instr_addr_o_31_(instr_addr_o[31]), .instr_addr_o_30_(
        instr_addr_o[30]), .instr_addr_o_29_(instr_addr_o[29]), 
        .instr_addr_o_28_(instr_addr_o[28]), .instr_addr_o_27_(
        instr_addr_o[27]), .instr_addr_o_26_(instr_addr_o[26]), 
        .instr_addr_o_25_(instr_addr_o[25]), .instr_addr_o_24_(
        instr_addr_o[24]), .instr_addr_o_23_(instr_addr_o[23]), 
        .instr_addr_o_22_(instr_addr_o[22]), .instr_addr_o_21_(
        instr_addr_o[21]), .instr_addr_o_20_(instr_addr_o[20]), 
        .instr_addr_o_19_(instr_addr_o[19]), .instr_addr_o_17_(
        instr_addr_o[17]), .instr_addr_o_16_(instr_addr_o[16]), 
        .instr_addr_o_15_(instr_addr_o[15]), .instr_addr_o_13_(
        instr_addr_o[13]), .instr_addr_o_12_(instr_addr_o[12]), 
        .instr_addr_o_11_(instr_addr_o[11]), .instr_addr_o_10_(
        instr_addr_o[10]), .instr_addr_o_9_(instr_addr_o[9]), 
        .instr_addr_o_8_(instr_addr_o[8]), .instr_addr_o_7_(instr_addr_o[7]), 
        .instr_addr_o_6_(instr_addr_o[6]), .instr_addr_o_5_(instr_addr_o[5]), 
        .data_addr_o_30_(data_addr_o[30]), .data_addr_o_29_(data_addr_o[29]), 
        .data_addr_o_28_(data_addr_o[28]), .data_addr_o_27_(data_addr_o[27]), 
        .data_addr_o_26_(data_addr_o[26]), .data_addr_o_25_(data_addr_o[25]), 
        .data_addr_o_24_(data_addr_o[24]), .data_addr_o_23_(data_addr_o[23]), 
        .data_addr_o_22_(data_addr_o[22]), .data_addr_o_21_(data_addr_o[21]), 
        .data_addr_o_20_(data_addr_o[20]), .data_addr_o_19_(data_addr_o[19]), 
        .data_addr_o_18_(data_addr_o[18]), .data_addr_o_17_(data_addr_o[17]), 
        .data_addr_o_16_(data_addr_o[16]), .data_addr_o_15_(data_addr_o[15]), 
        .data_addr_o_14_(data_addr_o[14]), .data_addr_o_13_(data_addr_o[13]), 
        .data_addr_o_12_(data_addr_o[12]), .data_addr_o_11_(data_addr_o[11]), 
        .data_addr_o_10_(data_addr_o[10]), .data_addr_o_9_(data_addr_o[9]), 
        .data_addr_o_8_(data_addr_o[8]), .data_addr_o_7_(data_addr_o[7]), 
        .data_addr_o_6_(data_addr_o[6]), .data_addr_o_5_(data_addr_o[5]), 
        .data_addr_o_4_(data_addr_o[4]), .data_addr_o_3_(data_addr_o[3]), 
        .data_addr_o_2_(data_addr_o[2]), .data_addr_o_1_(data_addr_o[1]), 
        .data_addr_o_0_(data_addr_o[0]), .instr_addr_o_18_(n316), 
        .instr_addr_o_14_(n317), .instr_addr_o_4_(n318), .data_addr_o_31_(n319) );
  BUF_X1 U26 ( .A(alu_operand_a_ex[9]), .Z(n312) );
  AND2_X1 U28 ( .A1(n351), .A2(alu_operand_b_ex[1]), .ZN(csr_addr[1]) );
  CLKBUF_X1 U29 ( .A(alu_operand_a_ex[31]), .Z(n349) );
  CLKBUF_X1 U30 ( .A(alu_operand_a_ex[15]), .Z(n255) );
  CLKBUF_X1 U31 ( .A(alu_operand_b_ex[9]), .Z(n350) );
  INV_X1 U32 ( .A(csr_access_ex), .ZN(n351) );
endmodule

