library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
 
entity misr is
-- NON HO ANCORA CAPITO COME FARLO
end misr;